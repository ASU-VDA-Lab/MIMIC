module fake_netlist_5_667_n_1793 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1793);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1793;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_20),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_41),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_79),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_22),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_5),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_4),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_95),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_50),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_32),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_45),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_6),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_135),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_47),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_54),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_57),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_54),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_9),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_82),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_149),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_55),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_62),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_84),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_33),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_120),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_96),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_74),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_20),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_134),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_55),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_71),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_153),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_170),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_88),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_46),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_19),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_122),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_124),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_176),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_26),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_119),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_172),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_89),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_118),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_139),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_98),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_2),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_101),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_165),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_86),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_97),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_146),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_152),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_175),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_133),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_5),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_72),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_67),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_111),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_61),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_25),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_87),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_78),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_22),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_75),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_48),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_94),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_174),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_127),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_167),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_129),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_14),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_51),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_2),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_1),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_44),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_51),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_19),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_35),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_38),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_39),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_114),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_65),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_141),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_109),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_52),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_26),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_158),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_93),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_30),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_21),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_154),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_47),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_21),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_42),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_35),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_11),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_0),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_150),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_132),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_128),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_31),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_155),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_10),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_23),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_0),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_50),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_49),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_42),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_13),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_56),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_207),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_213),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_212),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_221),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_1),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_243),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_225),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_312),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_198),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_182),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_228),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_198),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_229),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_198),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_232),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_256),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_196),
.B(n_6),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_260),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_279),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_231),
.B(n_7),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_328),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_255),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_294),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_263),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_265),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_216),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_198),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_275),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_289),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_214),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_214),
.Y(n_389)
);

BUFx6f_ASAP7_75t_SL g390 ( 
.A(n_344),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_214),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_295),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_214),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_187),
.Y(n_394)
);

BUFx6f_ASAP7_75t_SL g395 ( 
.A(n_344),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_219),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_187),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_231),
.B(n_8),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_258),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_258),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_220),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_258),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_258),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_258),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_348),
.B(n_10),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_298),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_269),
.B(n_12),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_190),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_300),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_178),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_310),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_313),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_186),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_222),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_227),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_209),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_215),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_190),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_247),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_253),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_191),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_272),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_280),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_230),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_282),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_191),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_193),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_250),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_182),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_235),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_182),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_304),
.B(n_13),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_184),
.B(n_15),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_241),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_237),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_223),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_384),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_383),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_396),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_354),
.B(n_344),
.Y(n_447)
);

BUFx8_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_378),
.B(n_242),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_434),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_365),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_401),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_419),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_420),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_370),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_434),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_R g467 ( 
.A(n_380),
.B(n_251),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_323),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_376),
.A2(n_233),
.B(n_184),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

BUFx8_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_177),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_403),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_406),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_430),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_436),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_364),
.B(n_433),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_440),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_361),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_353),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_359),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_R g490 ( 
.A(n_356),
.B(n_252),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_363),
.B(n_354),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_356),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_418),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_421),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_357),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_422),
.Y(n_498)
);

CKINVDCx11_ASAP7_75t_R g499 ( 
.A(n_360),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_357),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_398),
.A2(n_283),
.B(n_233),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_411),
.B(n_238),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_438),
.B(n_323),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_355),
.B(n_362),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_362),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_367),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_428),
.B(n_181),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_367),
.B(n_285),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_358),
.B(n_286),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_375),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_369),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_369),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_394),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_454),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_513),
.B(n_283),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_468),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_512),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_451),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_371),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_513),
.B(n_307),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_492),
.B(n_372),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_451),
.B(n_372),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_307),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_483),
.B(n_374),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_329),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_519),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_503),
.B(n_374),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_447),
.B(n_381),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_382),
.C(n_381),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

BUFx4f_ASAP7_75t_L g545 ( 
.A(n_503),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_468),
.B(n_323),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_448),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_489),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_385),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_503),
.A2(n_236),
.B1(n_223),
.B2(n_352),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_518),
.B(n_329),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_504),
.B(n_373),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_487),
.B(n_394),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_462),
.B(n_427),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_503),
.B(n_385),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_495),
.Y(n_562)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_449),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_462),
.B(n_427),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_452),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_516),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_493),
.B(n_386),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_488),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_476),
.B(n_323),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_487),
.B(n_323),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_459),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_496),
.B(n_392),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_497),
.B(n_392),
.Y(n_578)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_516),
.B(n_435),
.C(n_366),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_505),
.B(n_408),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_468),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_463),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_507),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_507),
.B(n_407),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_503),
.B(n_408),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_509),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_498),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_450),
.B(n_286),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_463),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_498),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_450),
.B(n_185),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_500),
.B(n_414),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_414),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_467),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_476),
.B(n_416),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_445),
.B(n_377),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_506),
.B(n_416),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_468),
.B(n_417),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_517),
.B(n_417),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_517),
.B(n_424),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_446),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_490),
.B(n_192),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_468),
.B(n_250),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_514),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_498),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_501),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_463),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_498),
.B(n_197),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_482),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_508),
.B(n_424),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_458),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_517),
.B(n_432),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_458),
.B(n_199),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_515),
.B(n_202),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_460),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_342),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_464),
.Y(n_629)
);

AND3x2_ASAP7_75t_L g630 ( 
.A(n_465),
.B(n_314),
.C(n_236),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_499),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_482),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_466),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_469),
.B(n_211),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_453),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_444),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_448),
.B(n_226),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_469),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_448),
.B(n_183),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_471),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_471),
.B(n_254),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_453),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_444),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_444),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_474),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_234),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_472),
.B(n_224),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_475),
.Y(n_650)
);

AND3x2_ASAP7_75t_L g651 ( 
.A(n_475),
.B(n_345),
.C(n_314),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_501),
.B(n_345),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_485),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_455),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_477),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_478),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_470),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_472),
.B(n_239),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_478),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_484),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_470),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_600),
.B(n_549),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_432),
.C(n_472),
.Y(n_664)
);

NOR2x1p5_ASAP7_75t_L g665 ( 
.A(n_600),
.B(n_456),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_553),
.A2(n_352),
.B(n_330),
.C(n_327),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_549),
.B(n_457),
.Y(n_667)
);

AO22x1_ASAP7_75t_L g668 ( 
.A1(n_537),
.A2(n_472),
.B1(n_315),
.B2(n_316),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_529),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_537),
.A2(n_284),
.B1(n_308),
.B2(n_306),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_531),
.B(n_501),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_541),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_638),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_638),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_537),
.A2(n_262),
.B1(n_305),
.B2(n_302),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_526),
.B(n_250),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_537),
.B(n_501),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_537),
.B(n_484),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_526),
.B(n_250),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_520),
.B(n_179),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_537),
.A2(n_270),
.B1(n_261),
.B2(n_266),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_540),
.A2(n_288),
.B1(n_281),
.B2(n_278),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_526),
.B(n_250),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_534),
.B(n_250),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_607),
.B(n_473),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_SL g686 ( 
.A1(n_571),
.A2(n_246),
.B1(n_349),
.B2(n_309),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_557),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_602),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_562),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_526),
.B(n_250),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_607),
.B(n_473),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_526),
.B(n_560),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_638),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_629),
.B(n_240),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_520),
.B(n_194),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_629),
.B(n_245),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_520),
.B(n_244),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_558),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_567),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_543),
.B(n_276),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_539),
.B(n_437),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_558),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_522),
.B(n_248),
.Y(n_703)
);

BUFx5_ASAP7_75t_L g704 ( 
.A(n_534),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_608),
.B(n_441),
.C(n_510),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_560),
.B(n_250),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_523),
.B(n_249),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_533),
.B(n_257),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_527),
.B(n_259),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_652),
.B(n_292),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_577),
.B(n_180),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_652),
.B(n_296),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_568),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_611),
.A2(n_331),
.B1(n_326),
.B2(n_311),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_577),
.B(n_180),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_528),
.B(n_301),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_608),
.B(n_480),
.C(n_486),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_542),
.A2(n_287),
.B1(n_267),
.B2(n_268),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_528),
.B(n_585),
.Y(n_719)
);

INVx8_ASAP7_75t_L g720 ( 
.A(n_586),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_589),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_622),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_R g723 ( 
.A(n_563),
.B(n_481),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_558),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_626),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_566),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_555),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_560),
.B(n_303),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_623),
.A2(n_290),
.B1(n_271),
.B2(n_273),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_623),
.B(n_188),
.C(n_195),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_583),
.B(n_320),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_583),
.B(n_322),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_570),
.B(n_274),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_559),
.A2(n_332),
.B1(n_189),
.B2(n_195),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_633),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_555),
.Y(n_737)
);

INVxp33_ASAP7_75t_L g738 ( 
.A(n_564),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_583),
.B(n_485),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_580),
.A2(n_299),
.B1(n_297),
.B2(n_293),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_566),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_578),
.B(n_277),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_560),
.B(n_291),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_592),
.B(n_485),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_625),
.B(n_188),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_592),
.B(n_491),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_592),
.B(n_491),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_634),
.Y(n_748)
);

INVx6_ASAP7_75t_L g749 ( 
.A(n_561),
.Y(n_749)
);

NOR2x2_ASAP7_75t_L g750 ( 
.A(n_554),
.B(n_395),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_566),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_573),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_604),
.B(n_491),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_640),
.B(n_343),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_573),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_604),
.B(n_200),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_573),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_611),
.A2(n_350),
.B1(n_351),
.B2(n_319),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_200),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_552),
.A2(n_319),
.B1(n_351),
.B2(n_347),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_560),
.B(n_581),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_625),
.B(n_203),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_650),
.Y(n_763)
);

AND2x6_ASAP7_75t_SL g764 ( 
.A(n_595),
.B(n_237),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_654),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_661),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_584),
.B(n_203),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_584),
.B(n_205),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_660),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_660),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_615),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_615),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_615),
.B(n_205),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_587),
.A2(n_597),
.B1(n_606),
.B2(n_554),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_647),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_647),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_561),
.B(n_237),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_532),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_653),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_614),
.A2(n_347),
.B(n_204),
.C(n_206),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_616),
.B(n_210),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_581),
.B(n_210),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_616),
.B(n_264),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_616),
.B(n_264),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_324),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_550),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_653),
.Y(n_789)
);

AND2x6_ASAP7_75t_SL g790 ( 
.A(n_605),
.B(n_201),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_618),
.B(n_324),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_656),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_554),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_656),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_581),
.B(n_340),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_618),
.B(n_340),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_581),
.B(n_341),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_545),
.A2(n_341),
.B1(n_321),
.B2(n_339),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_632),
.B(n_201),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_655),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_632),
.B(n_204),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_206),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_572),
.B(n_395),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_636),
.B(n_208),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_645),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_545),
.A2(n_325),
.B1(n_339),
.B2(n_338),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_657),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_645),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_636),
.B(n_208),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_581),
.B(n_325),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_621),
.B(n_92),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_636),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_554),
.A2(n_395),
.B1(n_338),
.B2(n_337),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_614),
.B(n_337),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_545),
.B(n_335),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_658),
.B(n_335),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_658),
.B(n_334),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_524),
.B(n_334),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_637),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_586),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_658),
.B(n_333),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_669),
.B(n_641),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_669),
.B(n_601),
.C(n_579),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_685),
.B(n_691),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_739),
.A2(n_548),
.B(n_658),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_698),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_744),
.A2(n_548),
.B(n_603),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_749),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_794),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_628),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_710),
.A2(n_563),
.B1(n_586),
.B2(n_524),
.Y(n_833)
);

NOR2x1p5_ASAP7_75t_SL g834 ( 
.A(n_704),
.B(n_590),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_782),
.A2(n_818),
.B(n_823),
.C(n_819),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_671),
.A2(n_530),
.B(n_534),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_746),
.A2(n_603),
.B(n_525),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_794),
.B(n_530),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_747),
.A2(n_538),
.B(n_525),
.Y(n_839)
);

AOI21x1_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_593),
.B(n_598),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_677),
.A2(n_613),
.B(n_643),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_753),
.A2(n_535),
.B(n_525),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_692),
.A2(n_538),
.B(n_546),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_692),
.A2(n_538),
.B(n_546),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_727),
.B(n_649),
.Y(n_845)
);

OAI321xp33_ASAP7_75t_L g846 ( 
.A1(n_700),
.A2(n_659),
.A3(n_639),
.B1(n_553),
.B2(n_572),
.C(n_610),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_737),
.B(n_586),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_780),
.B(n_609),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_761),
.A2(n_535),
.B(n_546),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_715),
.B(n_534),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_782),
.A2(n_617),
.B(n_659),
.C(n_639),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_780),
.B(n_609),
.Y(n_852)
);

CKINVDCx10_ASAP7_75t_R g853 ( 
.A(n_800),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_761),
.A2(n_535),
.B(n_569),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_775),
.A2(n_601),
.B1(n_648),
.B2(n_617),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_672),
.B(n_648),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_818),
.A2(n_648),
.B(n_637),
.C(n_644),
.Y(n_858)
);

OAI321xp33_ASAP7_75t_L g859 ( 
.A1(n_700),
.A2(n_644),
.A3(n_521),
.B1(n_574),
.B2(n_544),
.C(n_620),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_788),
.B(n_793),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_713),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_678),
.A2(n_719),
.B(n_684),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_809),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_662),
.A2(n_556),
.B(n_569),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_662),
.A2(n_556),
.B(n_569),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_732),
.A2(n_556),
.B(n_582),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_733),
.A2(n_582),
.B(n_565),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_723),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_687),
.B(n_612),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_L g871 ( 
.A1(n_745),
.A2(n_315),
.B(n_316),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_771),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_734),
.B(n_631),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_816),
.A2(n_588),
.B(n_547),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_701),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_756),
.A2(n_599),
.B(n_574),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_742),
.B(n_619),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_689),
.B(n_591),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_699),
.B(n_591),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_702),
.A2(n_599),
.B(n_576),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_813),
.B(n_619),
.Y(n_881)
);

OAI321xp33_ASAP7_75t_L g882 ( 
.A1(n_745),
.A2(n_565),
.A3(n_521),
.B1(n_544),
.B2(n_620),
.C(n_596),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_749),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_724),
.A2(n_596),
.B(n_576),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_749),
.Y(n_886)
);

INVx11_ASAP7_75t_L g887 ( 
.A(n_667),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_762),
.A2(n_646),
.B(n_317),
.C(n_318),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_720),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_663),
.B(n_317),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_721),
.B(n_594),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_722),
.B(n_594),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_726),
.A2(n_594),
.B(n_635),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_741),
.A2(n_594),
.B(n_635),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_680),
.B(n_333),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_680),
.B(n_651),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_803),
.A2(n_321),
.B(n_318),
.C(n_624),
.Y(n_897)
);

CKINVDCx10_ASAP7_75t_R g898 ( 
.A(n_778),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_751),
.A2(n_755),
.B(n_752),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_757),
.A2(n_635),
.B(n_624),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_SL g901 ( 
.A1(n_817),
.A2(n_811),
.B(n_690),
.C(n_676),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_635),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_630),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_776),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_769),
.A2(n_624),
.B(n_575),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_772),
.A2(n_624),
.B(n_575),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_817),
.A2(n_575),
.B(n_60),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_575),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_773),
.A2(n_59),
.B(n_162),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_783),
.A2(n_163),
.B(n_160),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_812),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_714),
.A2(n_159),
.B1(n_156),
.B2(n_151),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_714),
.A2(n_147),
.B1(n_140),
.B2(n_130),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_785),
.A2(n_126),
.B(n_116),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_682),
.A2(n_112),
.B(n_110),
.C(n_108),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_736),
.B(n_16),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_786),
.A2(n_104),
.B(n_100),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_822),
.B(n_90),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_777),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_720),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_787),
.A2(n_85),
.B(n_77),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_791),
.A2(n_63),
.B(n_18),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_708),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_796),
.A2(n_17),
.B(n_23),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_767),
.A2(n_17),
.B(n_24),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_768),
.A2(n_24),
.B(n_25),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_748),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_774),
.A2(n_743),
.B(n_814),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_717),
.B(n_27),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_SL g930 ( 
.A(n_686),
.B(n_28),
.C(n_31),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_743),
.A2(n_34),
.B(n_36),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_695),
.B(n_34),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_792),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_779),
.A2(n_37),
.B(n_43),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_805),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_781),
.A2(n_43),
.B(n_44),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_695),
.B(n_45),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_763),
.B(n_46),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_697),
.B(n_48),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_697),
.B(n_52),
.Y(n_940)
);

NOR2x1_ASAP7_75t_SL g941 ( 
.A(n_728),
.B(n_53),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_688),
.B(n_53),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_765),
.B(n_57),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_789),
.A2(n_693),
.B(n_674),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_673),
.A2(n_690),
.B(n_676),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_758),
.A2(n_766),
.B1(n_730),
.B2(n_681),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_735),
.A2(n_804),
.B(n_801),
.C(n_802),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_708),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_808),
.B(n_810),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_758),
.A2(n_670),
.B1(n_675),
.B2(n_799),
.Y(n_950)
);

OA21x2_ASAP7_75t_L g951 ( 
.A1(n_703),
.A2(n_709),
.B(n_707),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_738),
.B(n_705),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_728),
.A2(n_679),
.B(n_706),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_754),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_754),
.B(n_778),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_679),
.A2(n_706),
.B(n_683),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_694),
.B(n_696),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_740),
.B(n_807),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_760),
.A2(n_729),
.B(n_718),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_683),
.A2(n_784),
.B(n_795),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_784),
.A2(n_795),
.B(n_797),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_820),
.A2(n_811),
.B(n_666),
.C(n_716),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_778),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_821),
.A2(n_797),
.B(n_759),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_815),
.B(n_798),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_664),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_803),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_790),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_760),
.A2(n_665),
.B1(n_704),
.B2(n_750),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_SL g970 ( 
.A(n_704),
.B(n_723),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_704),
.A2(n_668),
.B(n_764),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_704),
.A2(n_671),
.B(n_710),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_704),
.A2(n_545),
.B(n_739),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_669),
.B(n_727),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_669),
.B(n_685),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_727),
.B(n_737),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_739),
.A2(n_545),
.B(n_744),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_727),
.B(n_737),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_794),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_775),
.B(n_662),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_669),
.B(n_727),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_669),
.A2(n_762),
.B(n_745),
.C(n_711),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_669),
.A2(n_762),
.B(n_745),
.C(n_711),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_739),
.A2(n_746),
.B(n_744),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_739),
.A2(n_545),
.B(n_744),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_794),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_739),
.A2(n_545),
.B(n_744),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_794),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_794),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_669),
.B(n_685),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_669),
.A2(n_762),
.B(n_745),
.C(n_711),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_794),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_669),
.B(n_727),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_749),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_669),
.B(n_727),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_669),
.B(n_685),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_739),
.A2(n_545),
.B(n_744),
.Y(n_997)
);

O2A1O1Ixp5_ASAP7_75t_L g998 ( 
.A1(n_669),
.A2(n_671),
.B(n_817),
.C(n_691),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_794),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_669),
.A2(n_502),
.B(n_745),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_671),
.A2(n_712),
.B(n_710),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_895),
.A2(n_1000),
.B(n_871),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_862),
.A2(n_1001),
.B(n_985),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_841),
.A2(n_894),
.B(n_984),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_840),
.A2(n_928),
.B(n_964),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_982),
.B(n_991),
.C(n_983),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_861),
.B(n_889),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_1001),
.A2(n_987),
.B(n_977),
.Y(n_1009)
);

AOI221xp5_ASAP7_75t_SL g1010 ( 
.A1(n_959),
.A2(n_940),
.B1(n_888),
.B2(n_965),
.C(n_932),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_975),
.B(n_990),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_875),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_889),
.B(n_920),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_998),
.A2(n_996),
.B(n_836),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_832),
.B(n_826),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_970),
.B(n_846),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_867),
.A2(n_866),
.B(n_973),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_875),
.B(n_976),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_830),
.Y(n_1020)
);

AO31x2_ASAP7_75t_L g1021 ( 
.A1(n_855),
.A2(n_950),
.A3(n_897),
.B(n_946),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_974),
.B(n_981),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_853),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_864),
.A2(n_865),
.B(n_997),
.Y(n_1024)
);

NOR2xp67_ASAP7_75t_L g1025 ( 
.A(n_868),
.B(n_846),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_837),
.A2(n_827),
.B(n_839),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_957),
.A2(n_850),
.B(n_836),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_993),
.B(n_995),
.Y(n_1028)
);

OA21x2_ASAP7_75t_L g1029 ( 
.A1(n_972),
.A2(n_882),
.B(n_859),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_920),
.B(n_830),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_972),
.A2(n_901),
.B(n_842),
.Y(n_1031)
);

AOI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_835),
.A2(n_952),
.B(n_824),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_978),
.B(n_896),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_970),
.B(n_967),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_979),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_830),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_882),
.A2(n_859),
.B(n_874),
.Y(n_1037)
);

AOI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_947),
.A2(n_869),
.B(n_833),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_949),
.B(n_857),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_961),
.A2(n_960),
.B(n_893),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_900),
.A2(n_953),
.B(n_945),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_920),
.B(n_918),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_825),
.B(n_870),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_860),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_986),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_872),
.B(n_904),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_SL g1047 ( 
.A(n_883),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_848),
.B(n_852),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_851),
.A2(n_927),
.B(n_939),
.C(n_937),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_907),
.A2(n_929),
.B(n_931),
.C(n_926),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_988),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_907),
.A2(n_924),
.B(n_925),
.C(n_930),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_899),
.A2(n_844),
.B(n_849),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_881),
.A2(n_877),
.B(n_829),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_919),
.B(n_933),
.Y(n_1055)
);

NAND2x1_ASAP7_75t_L g1056 ( 
.A(n_828),
.B(n_999),
.Y(n_1056)
);

AOI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_962),
.A2(n_969),
.B(n_845),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_955),
.B(n_847),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_935),
.B(n_916),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_843),
.A2(n_854),
.B(n_880),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_885),
.A2(n_944),
.B(n_956),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_938),
.B(n_943),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_878),
.A2(n_879),
.B(n_992),
.Y(n_1063)
);

AO21x1_ASAP7_75t_L g1064 ( 
.A1(n_922),
.A2(n_921),
.B(n_917),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_884),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_954),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_884),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_902),
.A2(n_892),
.B(n_891),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_884),
.B(n_994),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_989),
.B(n_918),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_858),
.A2(n_838),
.B(n_908),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_905),
.A2(n_906),
.B(n_910),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_980),
.B(n_847),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_856),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_923),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_980),
.B(n_923),
.Y(n_1076)
);

AND2x2_ASAP7_75t_SL g1077 ( 
.A(n_942),
.B(n_966),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_954),
.B(n_923),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_948),
.A2(n_887),
.B1(n_828),
.B2(n_863),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_914),
.A2(n_909),
.B(n_915),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_971),
.A2(n_942),
.B(n_913),
.C(n_912),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_911),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_934),
.A2(n_936),
.B(n_834),
.C(n_890),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_951),
.A2(n_873),
.B(n_980),
.Y(n_1084)
);

BUFx4_ASAP7_75t_SL g1085 ( 
.A(n_963),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_980),
.A2(n_941),
.B(n_966),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_948),
.A2(n_954),
.B(n_886),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_948),
.B(n_966),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_968),
.A2(n_983),
.B(n_991),
.C(n_982),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_903),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_898),
.A2(n_894),
.B(n_876),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_968),
.A2(n_998),
.B(n_983),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_968),
.A2(n_894),
.B(n_876),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_982),
.B(n_983),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_875),
.B(n_727),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_982),
.A2(n_991),
.B(n_983),
.C(n_669),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_861),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_998),
.A2(n_983),
.B(n_982),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_975),
.B(n_669),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_841),
.A2(n_894),
.B(n_984),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_982),
.A2(n_991),
.B(n_983),
.C(n_669),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_SL g1102 ( 
.A1(n_895),
.A2(n_669),
.B(n_542),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_875),
.B(n_727),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_841),
.A2(n_894),
.B(n_984),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_841),
.A2(n_894),
.B(n_984),
.Y(n_1105)
);

CKINVDCx6p67_ASAP7_75t_R g1106 ( 
.A(n_853),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_982),
.A2(n_983),
.B1(n_991),
.B2(n_669),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_853),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_972),
.A2(n_1001),
.B(n_983),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_998),
.A2(n_983),
.B(n_982),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_875),
.B(n_727),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_862),
.A2(n_545),
.B(n_1001),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_862),
.A2(n_545),
.B(n_1001),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_830),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_975),
.B(n_669),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1000),
.A2(n_669),
.B1(n_959),
.B2(n_958),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_982),
.A2(n_991),
.B(n_983),
.C(n_669),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_975),
.B(n_669),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_831),
.Y(n_1119)
);

CKINVDCx8_ASAP7_75t_R g1120 ( 
.A(n_853),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_828),
.B(n_979),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_868),
.B(n_788),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1000),
.A2(n_669),
.B1(n_958),
.B2(n_982),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_875),
.B(n_727),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_875),
.B(n_727),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_875),
.B(n_727),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_979),
.Y(n_1127)
);

OAI22x1_ASAP7_75t_L g1128 ( 
.A1(n_940),
.A2(n_669),
.B1(n_965),
.B2(n_895),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_831),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_1000),
.A2(n_669),
.B(n_982),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_830),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_982),
.B(n_983),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_889),
.B(n_920),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_861),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_998),
.A2(n_983),
.B(n_982),
.Y(n_1135)
);

XOR2xp5_ASAP7_75t_L g1136 ( 
.A(n_868),
.B(n_514),
.Y(n_1136)
);

BUFx4f_ASAP7_75t_SL g1137 ( 
.A(n_861),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_861),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_841),
.A2(n_894),
.B(n_984),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_853),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_975),
.B(n_669),
.Y(n_1141)
);

AOI21x1_ASAP7_75t_L g1142 ( 
.A1(n_841),
.A2(n_840),
.B(n_826),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_875),
.B(n_727),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1077),
.B(n_1016),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1096),
.A2(n_1117),
.B(n_1101),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1137),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1035),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1102),
.A2(n_1128),
.B1(n_1002),
.B2(n_1116),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_1141),
.B2(n_1118),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1019),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1042),
.B(n_1133),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1137),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1098),
.A2(n_1135),
.B(n_1110),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1106),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1011),
.B(n_1033),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1097),
.Y(n_1157)
);

AOI22x1_ASAP7_75t_L g1158 ( 
.A1(n_1092),
.A2(n_1031),
.B1(n_1027),
.B2(n_1009),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1039),
.B(n_1130),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1096),
.B(n_1101),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_1023),
.B(n_1108),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1133),
.B(n_1008),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1095),
.B(n_1103),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1117),
.B(n_1107),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1045),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1046),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1111),
.B(n_1124),
.Y(n_1167)
);

OAI22x1_ASAP7_75t_L g1168 ( 
.A1(n_1048),
.A2(n_1006),
.B1(n_1028),
.B2(n_1022),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1007),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1138),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1012),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1077),
.A2(n_1089),
.B1(n_1094),
.B2(n_1132),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1134),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1043),
.B(n_1022),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1042),
.B(n_1133),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1042),
.B(n_1078),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1076),
.B(n_1007),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1028),
.B(n_1062),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1023),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1089),
.A2(n_1094),
.B1(n_1132),
.B2(n_1081),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1108),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_1007),
.B(n_1073),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1065),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1012),
.B(n_1125),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_SL g1185 ( 
.A(n_1034),
.B(n_1059),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1126),
.B(n_1143),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_SL g1187 ( 
.A(n_1034),
.B(n_1017),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1055),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1058),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1008),
.B(n_1090),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1048),
.B(n_1066),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1010),
.B(n_1032),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1088),
.B(n_1049),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1112),
.A2(n_1113),
.B(n_1003),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_1017),
.B(n_1057),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1013),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1120),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1140),
.Y(n_1198)
);

INVx3_ASAP7_75t_R g1199 ( 
.A(n_1085),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_1140),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1081),
.A2(n_1049),
.B1(n_1029),
.B2(n_1037),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1085),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1067),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1029),
.A2(n_1037),
.B1(n_1050),
.B2(n_1070),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1038),
.B(n_1075),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1067),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1029),
.A2(n_1037),
.B1(n_1050),
.B2(n_1052),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1025),
.A2(n_1044),
.B1(n_1090),
.B2(n_1109),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1067),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1066),
.B(n_1075),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1122),
.B(n_1082),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1036),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1047),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1014),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_1114),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1047),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1114),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1136),
.B(n_1079),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1051),
.B(n_1119),
.Y(n_1219)
);

HAxp5_ASAP7_75t_L g1220 ( 
.A(n_1069),
.B(n_1020),
.CON(n_1220),
.SN(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1074),
.B(n_1069),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1131),
.B(n_1030),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1014),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1052),
.B(n_1030),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1129),
.B(n_1087),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1083),
.A2(n_1086),
.B(n_1084),
.C(n_1071),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1127),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1127),
.A2(n_1083),
.B1(n_1121),
.B2(n_1056),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1093),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1021),
.B(n_1068),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1054),
.B(n_1142),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_1091),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1040),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1021),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1021),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1021),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1064),
.B(n_1063),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1072),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1041),
.B(n_1024),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1041),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_1026),
.B1(n_1018),
.B2(n_1061),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1005),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1053),
.A2(n_1080),
.B(n_1060),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1004),
.B(n_1100),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1004),
.Y(n_1245)
);

AOI222xp33_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_1102),
.B1(n_1000),
.B2(n_1128),
.C1(n_686),
.C2(n_1077),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1104),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1105),
.A2(n_1102),
.B(n_983),
.C(n_991),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1139),
.A2(n_1123),
.B1(n_1116),
.B2(n_983),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_983),
.B2(n_991),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1106),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1137),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1102),
.A2(n_669),
.B1(n_1128),
.B2(n_1002),
.Y(n_1256)
);

AOI221x1_ASAP7_75t_L g1257 ( 
.A1(n_1128),
.A2(n_1107),
.B1(n_983),
.B2(n_991),
.C(n_982),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_983),
.B2(n_991),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1012),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1076),
.B(n_1007),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1137),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1106),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_983),
.B2(n_991),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1035),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1137),
.Y(n_1266)
);

AOI222xp33_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_1000),
.B1(n_1128),
.B2(n_686),
.C1(n_1077),
.C2(n_669),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1065),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1035),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1019),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1033),
.B(n_1019),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1016),
.B(n_875),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1042),
.B(n_1133),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1023),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1046),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_983),
.B2(n_991),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_SL g1281 ( 
.A(n_1106),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_983),
.B2(n_991),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1033),
.B(n_1019),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1102),
.B(n_669),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1008),
.Y(n_1285)
);

BUFx8_ASAP7_75t_SL g1286 ( 
.A(n_1278),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1145),
.B(n_1172),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1219),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1197),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1196),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1284),
.A2(n_1174),
.B1(n_1254),
.B2(n_1255),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1173),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1227),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1256),
.A2(n_1267),
.B(n_1148),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1267),
.A2(n_1251),
.B1(n_1258),
.B2(n_1264),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1259),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1200),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1169),
.B(n_1209),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1147),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1274),
.B(n_1283),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1153),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1165),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1200),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1251),
.A2(n_1264),
.B1(n_1282),
.B2(n_1280),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1209),
.Y(n_1306)
);

BUFx8_ASAP7_75t_L g1307 ( 
.A(n_1202),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1161),
.Y(n_1308)
);

AOI222xp33_ASAP7_75t_L g1309 ( 
.A1(n_1258),
.A2(n_1280),
.B1(n_1282),
.B2(n_1172),
.C1(n_1156),
.C2(n_1168),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1253),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1149),
.A2(n_1272),
.B1(n_1273),
.B2(n_1275),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1179),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1265),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1269),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1246),
.A2(n_1180),
.B1(n_1150),
.B2(n_1164),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1166),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1252),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1157),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1235),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1163),
.B(n_1167),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1152),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1215),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1281),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1279),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1246),
.A2(n_1164),
.B1(n_1154),
.B2(n_1144),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1216),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1175),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1277),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1195),
.A2(n_1249),
.B(n_1192),
.C(n_1178),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1276),
.B(n_1184),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1262),
.B(n_1270),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1154),
.A2(n_1160),
.B1(n_1195),
.B2(n_1159),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1221),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1186),
.B(n_1151),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1241),
.A2(n_1243),
.B(n_1239),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1262),
.A2(n_1270),
.B1(n_1208),
.B2(n_1171),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1225),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1277),
.B(n_1176),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1176),
.B(n_1190),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1237),
.A2(n_1250),
.B(n_1204),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1191),
.Y(n_1342)
);

OR2x6_ASAP7_75t_L g1343 ( 
.A(n_1177),
.B(n_1260),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1170),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1210),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1193),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1257),
.A2(n_1226),
.B(n_1158),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1214),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1271),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1218),
.A2(n_1160),
.B(n_1211),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1159),
.A2(n_1201),
.B1(n_1236),
.B2(n_1205),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1233),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1224),
.A2(n_1201),
.B1(n_1187),
.B2(n_1207),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1189),
.B(n_1260),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1224),
.A2(n_1207),
.B1(n_1234),
.B2(n_1182),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1190),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1155),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1182),
.A2(n_1260),
.B1(n_1177),
.B2(n_1204),
.Y(n_1359)
);

CKINVDCx8_ASAP7_75t_R g1360 ( 
.A(n_1181),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1229),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1185),
.A2(n_1213),
.B1(n_1177),
.B2(n_1182),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_1212),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1199),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1229),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1213),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1222),
.B(n_1285),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1263),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1198),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1228),
.A2(n_1247),
.B(n_1244),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1238),
.B(n_1223),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1206),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1217),
.B(n_1214),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1162),
.B(n_1220),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1203),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1285),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1231),
.A2(n_1247),
.B(n_1244),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1203),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_R g1379 ( 
.A1(n_1146),
.A2(n_1266),
.B1(n_1261),
.B2(n_1240),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1268),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1206),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1268),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1214),
.A2(n_1232),
.B1(n_1183),
.B2(n_1242),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1232),
.A2(n_1242),
.B1(n_1248),
.B2(n_1245),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1248),
.A2(n_1102),
.B(n_669),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1219),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1219),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1174),
.B(n_1099),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1219),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1284),
.A2(n_1128),
.B1(n_1116),
.B2(n_1002),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1152),
.B(n_1175),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1219),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1172),
.A2(n_1077),
.B1(n_942),
.B2(n_669),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1194),
.A2(n_1110),
.B(n_1098),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1219),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1219),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1219),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1152),
.B(n_1175),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1342),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1291),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1292),
.B(n_1332),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1306),
.Y(n_1402)
);

BUFx2_ASAP7_75t_SL g1403 ( 
.A(n_1306),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1296),
.B(n_1287),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1306),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1306),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1296),
.B(n_1287),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1320),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1287),
.B(n_1305),
.Y(n_1409)
);

BUFx8_ASAP7_75t_L g1410 ( 
.A(n_1290),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1305),
.B(n_1353),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1353),
.B(n_1333),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1311),
.B(n_1388),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1333),
.B(n_1351),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1331),
.B(n_1288),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1371),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1343),
.B(n_1371),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1393),
.A2(n_1337),
.B1(n_1295),
.B2(n_1374),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1361),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1341),
.A2(n_1370),
.B(n_1330),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1318),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1394),
.B(n_1347),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1351),
.B(n_1309),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1394),
.A2(n_1352),
.B(n_1365),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1334),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1371),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1289),
.B(n_1386),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1338),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1377),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1294),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1359),
.A2(n_1356),
.B(n_1346),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1330),
.B(n_1350),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1356),
.A2(n_1326),
.B(n_1315),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1343),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1354),
.B(n_1345),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1359),
.B(n_1346),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1336),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1355),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1335),
.B(n_1390),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1393),
.A2(n_1390),
.B1(n_1379),
.B2(n_1354),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1336),
.A2(n_1395),
.B(n_1397),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1389),
.A2(n_1392),
.B(n_1396),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1316),
.B(n_1319),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1301),
.B(n_1321),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1325),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1297),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1300),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1360),
.B(n_1290),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1358),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1349),
.B(n_1297),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1303),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1313),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1314),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1384),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1312),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1384),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1383),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1376),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1380),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1383),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1293),
.Y(n_1463)
);

AOI21xp33_ASAP7_75t_L g1464 ( 
.A1(n_1362),
.A2(n_1375),
.B(n_1382),
.Y(n_1464)
);

INVx3_ASAP7_75t_SL g1465 ( 
.A(n_1381),
.Y(n_1465)
);

INVxp67_ASAP7_75t_R g1466 ( 
.A(n_1298),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1344),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1299),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1362),
.B(n_1357),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1378),
.A2(n_1367),
.B(n_1340),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1367),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1348),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1443),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1401),
.B(n_1372),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1443),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1412),
.B(n_1329),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1412),
.B(n_1322),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1413),
.B(n_1328),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1470),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1470),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_SL g1481 ( 
.A1(n_1444),
.A2(n_1416),
.B(n_1453),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1461),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1470),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1432),
.A2(n_1339),
.B(n_1391),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1470),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1422),
.B(n_1339),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1425),
.B(n_1398),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1425),
.B(n_1391),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_SL g1489 ( 
.A(n_1423),
.B(n_1364),
.Y(n_1489)
);

NOR4xp25_ASAP7_75t_SL g1490 ( 
.A(n_1430),
.B(n_1308),
.C(n_1312),
.D(n_1369),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1451),
.Y(n_1491)
);

CKINVDCx8_ASAP7_75t_R g1492 ( 
.A(n_1403),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1423),
.A2(n_1298),
.B1(n_1366),
.B2(n_1304),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1442),
.B(n_1366),
.Y(n_1494)
);

AOI222xp33_ASAP7_75t_L g1495 ( 
.A1(n_1424),
.A2(n_1441),
.B1(n_1404),
.B2(n_1407),
.C1(n_1414),
.C2(n_1409),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1429),
.B(n_1323),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1408),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1447),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1424),
.A2(n_1327),
.B1(n_1302),
.B2(n_1310),
.C(n_1363),
.Y(n_1499)
);

NOR2x2_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_1304),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1420),
.B(n_1373),
.Y(n_1501)
);

AND2x4_ASAP7_75t_SL g1502 ( 
.A(n_1417),
.B(n_1364),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1420),
.B(n_1310),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1408),
.B(n_1302),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1420),
.B(n_1414),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1419),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1489),
.A2(n_1433),
.B1(n_1418),
.B2(n_1495),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1505),
.B(n_1456),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1495),
.B(n_1433),
.C(n_1442),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1482),
.B(n_1474),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1426),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1489),
.B(n_1417),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1415),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1456),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1493),
.A2(n_1407),
.B(n_1404),
.Y(n_1515)
);

NAND4xp25_ASAP7_75t_SL g1516 ( 
.A(n_1493),
.B(n_1440),
.C(n_1459),
.D(n_1462),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1505),
.B(n_1419),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1476),
.B(n_1458),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1458),
.Y(n_1520)
);

OAI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1499),
.A2(n_1440),
.B1(n_1435),
.B2(n_1416),
.C(n_1450),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1499),
.B(n_1434),
.C(n_1429),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1523)
);

NOR3xp33_ASAP7_75t_L g1524 ( 
.A(n_1494),
.B(n_1427),
.C(n_1464),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1494),
.A2(n_1469),
.B1(n_1462),
.B2(n_1409),
.C(n_1436),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1478),
.B(n_1434),
.C(n_1448),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1504),
.B(n_1436),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1504),
.B(n_1437),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1504),
.B(n_1437),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1478),
.A2(n_1434),
.B1(n_1469),
.B2(n_1463),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1452),
.C(n_1399),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1439),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1487),
.B(n_1488),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1498),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1490),
.B(n_1463),
.C(n_1428),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1446),
.C(n_1467),
.D(n_1421),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1492),
.A2(n_1445),
.B1(n_1466),
.B2(n_1411),
.Y(n_1537)
);

OA211x2_ASAP7_75t_L g1538 ( 
.A1(n_1496),
.A2(n_1492),
.B(n_1466),
.C(n_1500),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_L g1539 ( 
.A(n_1503),
.B(n_1400),
.C(n_1454),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1486),
.B(n_1438),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1491),
.B(n_1421),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1480),
.B(n_1483),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1497),
.B(n_1431),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1503),
.B(n_1449),
.C(n_1455),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1480),
.B(n_1438),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1503),
.B(n_1449),
.C(n_1455),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1502),
.A2(n_1471),
.B1(n_1427),
.B2(n_1411),
.Y(n_1548)
);

NOR3xp33_ASAP7_75t_L g1549 ( 
.A(n_1501),
.B(n_1427),
.C(n_1468),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1545),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1544),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1534),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1533),
.B(n_1483),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1539),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1534),
.B(n_1479),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1543),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1542),
.A2(n_1485),
.B(n_1479),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1543),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1542),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1544),
.Y(n_1561)
);

AND2x4_ASAP7_75t_SL g1562 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1547),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1460),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1507),
.A2(n_1502),
.B1(n_1410),
.B2(n_1491),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1509),
.A2(n_1502),
.B1(n_1481),
.B2(n_1484),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1517),
.B(n_1473),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1484),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1484),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.B(n_1484),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1539),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1546),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1528),
.B(n_1473),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1475),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1551),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1569),
.B(n_1508),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1569),
.B(n_1514),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1562),
.B(n_1540),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1552),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1568),
.B(n_1575),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1568),
.B(n_1510),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1568),
.B(n_1527),
.Y(n_1585)
);

O2A1O1Ixp5_ASAP7_75t_L g1586 ( 
.A1(n_1551),
.A2(n_1525),
.B(n_1526),
.C(n_1512),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1552),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1514),
.Y(n_1590)
);

NAND2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1572),
.B(n_1501),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1518),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1523),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1552),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1566),
.A2(n_1509),
.B(n_1522),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1570),
.B(n_1518),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1556),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1556),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1556),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1560),
.B(n_1553),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1520),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1558),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1520),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1557),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1558),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1557),
.B(n_1513),
.Y(n_1608)
);

AOI32xp33_ASAP7_75t_L g1609 ( 
.A1(n_1572),
.A2(n_1530),
.A3(n_1524),
.B1(n_1537),
.B2(n_1521),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1557),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1559),
.B(n_1526),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1559),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1558),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1606),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1606),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1592),
.B(n_1608),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1577),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1610),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1610),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1612),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1597),
.A2(n_1565),
.B1(n_1522),
.B2(n_1566),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1574),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1587),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1590),
.B(n_1574),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1612),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1602),
.B(n_1553),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1587),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1595),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1580),
.A2(n_1516),
.B1(n_1565),
.B2(n_1537),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1561),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1595),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1611),
.B(n_1561),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1577),
.B(n_1573),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1595),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1602),
.B(n_1553),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1581),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1561),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1581),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1588),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1609),
.B(n_1563),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1589),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1580),
.B(n_1553),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1593),
.B(n_1584),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1580),
.B(n_1554),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1589),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1585),
.B(n_1567),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1621),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.B(n_1593),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1646),
.B(n_1594),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1661)
);

INVx3_ASAP7_75t_SL g1662 ( 
.A(n_1649),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1585),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1615),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.Y(n_1665)
);

INVx5_ASAP7_75t_L g1666 ( 
.A(n_1618),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1627),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1650),
.B(n_1594),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1639),
.B(n_1567),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1515),
.B1(n_1591),
.B2(n_1538),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1639),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1641),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1619),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1649),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1638),
.A2(n_1567),
.B1(n_1530),
.B2(n_1591),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1584),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1615),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1599),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1616),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1618),
.B(n_1586),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1616),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1578),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1578),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1648),
.B(n_1599),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1629),
.B(n_1596),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1653),
.B(n_1596),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1622),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1631),
.B(n_1575),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1657),
.Y(n_1690)
);

CKINVDCx16_ASAP7_75t_R g1691 ( 
.A(n_1652),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1657),
.B(n_1575),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_1652),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1662),
.B(n_1644),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1667),
.A2(n_1586),
.B(n_1655),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1675),
.A2(n_1591),
.B1(n_1515),
.B2(n_1531),
.Y(n_1696)
);

AOI222xp33_ASAP7_75t_L g1697 ( 
.A1(n_1675),
.A2(n_1562),
.B1(n_1620),
.B2(n_1644),
.C1(n_1564),
.C2(n_1531),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1662),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1681),
.A2(n_1655),
.B(n_1591),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1670),
.A2(n_1538),
.B1(n_1564),
.B2(n_1562),
.Y(n_1700)
);

INVxp33_ASAP7_75t_SL g1701 ( 
.A(n_1674),
.Y(n_1701)
);

NOR4xp25_ASAP7_75t_SL g1702 ( 
.A(n_1681),
.B(n_1623),
.C(n_1622),
.D(n_1624),
.Y(n_1702)
);

AOI221x1_ASAP7_75t_L g1703 ( 
.A1(n_1658),
.A2(n_1632),
.B1(n_1624),
.B2(n_1623),
.C(n_1643),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1672),
.A2(n_1358),
.B(n_1324),
.C(n_1541),
.Y(n_1704)
);

AO21x1_ASAP7_75t_L g1705 ( 
.A1(n_1669),
.A2(n_1632),
.B(n_1607),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1680),
.Y(n_1706)
);

OAI322xp33_ASAP7_75t_L g1707 ( 
.A1(n_1660),
.A2(n_1668),
.A3(n_1671),
.B1(n_1690),
.B2(n_1669),
.C1(n_1676),
.C2(n_1692),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1664),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1666),
.Y(n_1710)
);

OAI31xp33_ASAP7_75t_L g1711 ( 
.A1(n_1661),
.A2(n_1562),
.A3(n_1654),
.B(n_1536),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1666),
.A2(n_1535),
.B(n_1614),
.C(n_1604),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1691),
.B(n_1654),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1666),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1659),
.A2(n_1601),
.B(n_1600),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1693),
.B(n_1600),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1666),
.A2(n_1535),
.B1(n_1601),
.B2(n_1502),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1679),
.A2(n_1614),
.B1(n_1607),
.B2(n_1604),
.C(n_1645),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1661),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1698),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1701),
.B(n_1286),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1706),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1698),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1714),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1694),
.B(n_1663),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1708),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1710),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1709),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1702),
.A2(n_1687),
.B1(n_1686),
.B2(n_1684),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1683),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1703),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1695),
.B(n_1683),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1704),
.B(n_1286),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1707),
.B(n_1317),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1682),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1716),
.B(n_1688),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1705),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1700),
.B(n_1689),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1730),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1731),
.A2(n_1696),
.B1(n_1699),
.B2(n_1712),
.C(n_1715),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1738),
.A2(n_1696),
.B1(n_1718),
.B2(n_1711),
.C(n_1717),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1732),
.A2(n_1457),
.B(n_1678),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1735),
.A2(n_1685),
.B(n_1678),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1735),
.A2(n_1685),
.B(n_1665),
.C(n_1673),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1722),
.B(n_1596),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1720),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1727),
.B(n_1598),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1736),
.A2(n_1673),
.B(n_1665),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1723),
.A2(n_1614),
.B1(n_1607),
.B2(n_1604),
.C(n_1548),
.Y(n_1750)
);

OAI321xp33_ASAP7_75t_L g1751 ( 
.A1(n_1729),
.A2(n_1643),
.A3(n_1640),
.B1(n_1636),
.B2(n_1619),
.C(n_1630),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1747),
.B(n_1721),
.C(n_1724),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1741),
.A2(n_1737),
.B1(n_1739),
.B2(n_1726),
.C(n_1728),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1742),
.B(n_1724),
.C(n_1721),
.Y(n_1754)
);

XNOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1740),
.B(n_1725),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1744),
.A2(n_1733),
.B1(n_1734),
.B2(n_1739),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1749),
.B(n_1745),
.C(n_1743),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1746),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1748),
.A2(n_1733),
.B1(n_1750),
.B2(n_1457),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_L g1760 ( 
.A(n_1751),
.B(n_1324),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1742),
.A2(n_1656),
.B1(n_1651),
.B2(n_1645),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1740),
.Y(n_1762)
);

OAI211xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1761),
.A2(n_1410),
.B(n_1636),
.C(n_1640),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1753),
.A2(n_1635),
.B1(n_1628),
.B2(n_1630),
.C(n_1625),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1757),
.A2(n_1754),
.B(n_1752),
.C(n_1756),
.Y(n_1765)
);

NOR3x1_ASAP7_75t_L g1766 ( 
.A(n_1759),
.B(n_1762),
.C(n_1758),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1760),
.B(n_1410),
.C(n_1368),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1765),
.A2(n_1755),
.B1(n_1317),
.B2(n_1368),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1656),
.B1(n_1651),
.B2(n_1637),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1766),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1763),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1764),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1766),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1770),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1768),
.B(n_1560),
.Y(n_1775)
);

OAI222xp33_ASAP7_75t_L g1776 ( 
.A1(n_1773),
.A2(n_1625),
.B1(n_1628),
.B2(n_1637),
.C1(n_1635),
.C2(n_1647),
.Y(n_1776)
);

XNOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1771),
.B(n_1307),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1772),
.B(n_1560),
.Y(n_1778)
);

AND2x2_ASAP7_75t_SL g1779 ( 
.A(n_1774),
.B(n_1769),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1774),
.B(n_1307),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1780),
.A2(n_1775),
.B1(n_1778),
.B2(n_1776),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1782),
.B(n_1781),
.C(n_1779),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1465),
.B1(n_1647),
.B2(n_1613),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1783),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1465),
.B1(n_1613),
.B2(n_1550),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1784),
.B(n_1613),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1786),
.A2(n_1465),
.B1(n_1578),
.B2(n_1579),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1787),
.A2(n_1579),
.B(n_1605),
.Y(n_1789)
);

AOI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1788),
.A2(n_1576),
.B(n_1575),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1790),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1789),
.B1(n_1579),
.B2(n_1603),
.Y(n_1792)
);

AOI211xp5_ASAP7_75t_L g1793 ( 
.A1(n_1792),
.A2(n_1402),
.B(n_1406),
.C(n_1405),
.Y(n_1793)
);


endmodule