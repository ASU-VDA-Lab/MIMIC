module fake_jpeg_17243_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_20),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_56),
.B1(n_36),
.B2(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_30),
.B1(n_21),
.B2(n_26),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_58),
.B1(n_36),
.B2(n_37),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_82),
.Y(n_106)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_36),
.B1(n_33),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_84),
.B1(n_88),
.B2(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_39),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_39),
.C(n_35),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_35),
.C(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_39),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_48),
.B1(n_54),
.B2(n_53),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_99)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_26),
.B1(n_24),
.B2(n_37),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_54),
.B1(n_48),
.B2(n_3),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_37),
.B1(n_24),
.B2(n_27),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_110),
.C(n_87),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_23),
.B(n_20),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_120),
.Y(n_122)
);

OR2x4_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_23),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_113),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_111),
.B1(n_114),
.B2(n_92),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_35),
.B1(n_23),
.B2(n_20),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_35),
.B1(n_19),
.B2(n_3),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_35),
.B1(n_2),
.B2(n_4),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_35),
.B1(n_15),
.B2(n_6),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_92),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_136),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_67),
.B1(n_91),
.B2(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_98),
.B1(n_97),
.B2(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_75),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_100),
.B(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_158),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_126),
.C(n_129),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_101),
.B1(n_63),
.B2(n_70),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_132),
.B1(n_101),
.B2(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_99),
.B1(n_108),
.B2(n_104),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_128),
.B1(n_143),
.B2(n_135),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_120),
.B(n_74),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_8),
.Y(n_183)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_128),
.B1(n_122),
.B2(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_157),
.B1(n_155),
.B2(n_147),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_122),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_181),
.C(n_152),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_121),
.B1(n_125),
.B2(n_107),
.Y(n_182)
);

OAI322xp33_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_184),
.A3(n_185),
.B1(n_166),
.B2(n_156),
.C1(n_150),
.C2(n_182),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_145),
.C(n_60),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_153),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_176),
.B(n_164),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_146),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_152),
.C(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_150),
.C(n_157),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_170),
.B1(n_155),
.B2(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_165),
.B1(n_162),
.B2(n_88),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_188),
.C(n_191),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_185),
.B(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_183),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_177),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_199),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_188),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_205),
.C(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_192),
.C(n_64),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_60),
.C(n_73),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_225),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_14),
.C(n_10),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_220),
.B1(n_219),
.B2(n_11),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_229),
.Y(n_235)
);

OAI211xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_226),
.B(n_224),
.C(n_14),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_231),
.C(n_226),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_234),
.B(n_9),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_13),
.Y(n_238)
);


endmodule