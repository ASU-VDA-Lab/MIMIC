module fake_netlist_6_1015_n_1820 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1820);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1820;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1632;
wire n_1805;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g488 ( 
.A(n_333),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_412),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_178),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_434),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_165),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_249),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_392),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_406),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_243),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_196),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_255),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_9),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_158),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_304),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_1),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_371),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_430),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_139),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_471),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_59),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_270),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_79),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_22),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_193),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_476),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_259),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_264),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_157),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_87),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_283),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_300),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_451),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_403),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_443),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_159),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_311),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_59),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_384),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_204),
.Y(n_528)
);

CKINVDCx14_ASAP7_75t_R g529 ( 
.A(n_273),
.Y(n_529)
);

BUFx5_ASAP7_75t_L g530 ( 
.A(n_239),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_474),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_186),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_121),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_302),
.Y(n_534)
);

CKINVDCx6p67_ASAP7_75t_R g535 ( 
.A(n_37),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_428),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_271),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_71),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_315),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_185),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_452),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_375),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_212),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_223),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_246),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_366),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_344),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_8),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_312),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_195),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_341),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_365),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_385),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_120),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_118),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_51),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_103),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_469),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_203),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_288),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_388),
.Y(n_561)
);

BUFx5_ASAP7_75t_L g562 ( 
.A(n_240),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_133),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_138),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_303),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_290),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_34),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_429),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_111),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_446),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_276),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_138),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_101),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_374),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_331),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_89),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_97),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_199),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_450),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_219),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_437),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_285),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_350),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_442),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_78),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_461),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_345),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_192),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_182),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_232),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_351),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_468),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_338),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_143),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_414),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_181),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_404),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_295),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_334),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_449),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_487),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_116),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_417),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_453),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_68),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_372),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_420),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_64),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_370),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_379),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_151),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_433),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_386),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_235),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_306),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_75),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_431),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_11),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_90),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_152),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_445),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_117),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_320),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_211),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_256),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_71),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_263),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_74),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_214),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_145),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_150),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_201),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_29),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_358),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_151),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_407),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_132),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_346),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_143),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_280),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_179),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_464),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_377),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_359),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_207),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_357),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_118),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_164),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_31),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_241),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_102),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_480),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_66),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_335),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_7),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_463),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_459),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_269),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_36),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_427),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_161),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_153),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_382),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_67),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_230),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_129),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_210),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_298),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_141),
.Y(n_673)
);

CKINVDCx14_ASAP7_75t_R g674 ( 
.A(n_106),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_25),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_438),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_174),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_277),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_401),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_339),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_477),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_177),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_408),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_321),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_310),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_3),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_113),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_25),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_308),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_202),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_247),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_332),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_267),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_1),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_7),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_525),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_674),
.B(n_0),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_491),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_586),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_529),
.B(n_183),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_564),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_674),
.B(n_0),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_494),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_643),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_586),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_535),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_564),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_586),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_501),
.B(n_2),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_695),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_695),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_681),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_495),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_639),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_695),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_695),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_490),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_500),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_508),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_510),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_639),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_496),
.Y(n_724)
);

XNOR2xp5_ASAP7_75t_L g725 ( 
.A(n_653),
.B(n_492),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_533),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_498),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_530),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_538),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_554),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_653),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_556),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_503),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_563),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_506),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_548),
.B(n_2),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_504),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_506),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_517),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_574),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_597),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_652),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_509),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_513),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_606),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_612),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_584),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_514),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_548),
.B(n_3),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_499),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_584),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_663),
.B(n_4),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_519),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_521),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_530),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_522),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_632),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_523),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_532),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_581),
.B(n_4),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_634),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_635),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_502),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_5),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_667),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_536),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_537),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_663),
.B(n_5),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_512),
.B(n_6),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_505),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_641),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_511),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_688),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_694),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_652),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_601),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_516),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_698),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_753),
.B(n_529),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_703),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_714),
.B(n_520),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_710),
.B(n_547),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_764),
.B(n_547),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_R g791 ( 
.A(n_774),
.B(n_683),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_736),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_724),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_768),
.B(n_683),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_727),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_734),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_738),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_705),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_713),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_713),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_728),
.A2(n_589),
.B(n_515),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_704),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_745),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_746),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_R g805 ( 
.A(n_774),
.B(n_527),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_706),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_751),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_757),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_713),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_736),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

BUFx8_ASAP7_75t_L g812 ( 
.A(n_718),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_767),
.B(n_488),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_776),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_758),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_712),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_739),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_716),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_717),
.Y(n_820)
);

CKINVDCx6p67_ASAP7_75t_R g821 ( 
.A(n_739),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_719),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_760),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_728),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_750),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_507),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_763),
.B(n_553),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_759),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_720),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_776),
.B(n_782),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_721),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_737),
.B(n_488),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_726),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_729),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_759),
.B(n_681),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_730),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_697),
.B(n_681),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_732),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_790),
.B(n_782),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_790),
.B(n_770),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_802),
.B(n_740),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_825),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_800),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_789),
.B(n_702),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_833),
.B(n_822),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_789),
.B(n_794),
.Y(n_847)
);

AO21x2_ASAP7_75t_L g848 ( 
.A1(n_788),
.A2(n_700),
.B(n_773),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_783),
.B(n_786),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_800),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_834),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_837),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_800),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_794),
.B(n_828),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_838),
.B(n_771),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_784),
.B(n_769),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_825),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_829),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_829),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_839),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_838),
.B(n_827),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_832),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_819),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_838),
.B(n_696),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_813),
.B(n_744),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_791),
.B(n_515),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_814),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_791),
.B(n_780),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_838),
.B(n_489),
.Y(n_869)
);

INVx5_ASAP7_75t_L g870 ( 
.A(n_836),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_811),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_832),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_833),
.B(n_722),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_833),
.B(n_707),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_801),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_805),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_R g877 ( 
.A(n_831),
.B(n_805),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_824),
.B(n_600),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_787),
.B(n_733),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_831),
.B(n_707),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_811),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_832),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_810),
.B(n_578),
.Y(n_884)
);

AND2x2_ASAP7_75t_SL g885 ( 
.A(n_785),
.B(n_589),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_832),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_819),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_811),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_785),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_830),
.B(n_666),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_838),
.B(n_531),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_830),
.B(n_687),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_798),
.A2(n_666),
.B1(n_658),
.B2(n_591),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_835),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_806),
.B(n_591),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_793),
.B(n_658),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_799),
.B(n_642),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_835),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_817),
.B(n_735),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_835),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_799),
.B(n_539),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_811),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_835),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_795),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

BUFx8_ASAP7_75t_SL g907 ( 
.A(n_792),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_796),
.B(n_741),
.Y(n_908)
);

INVx4_ASAP7_75t_SL g909 ( 
.A(n_836),
.Y(n_909)
);

BUFx10_ASAP7_75t_L g910 ( 
.A(n_797),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_803),
.B(n_742),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_809),
.B(n_815),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_815),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_809),
.B(n_541),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_836),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_836),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_836),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_804),
.B(n_743),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_807),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_854),
.A2(n_816),
.B1(n_823),
.B2(n_808),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_854),
.B(n_672),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_918),
.B(n_812),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_847),
.B(n_672),
.Y(n_923)
);

OAI22xp33_ASAP7_75t_L g924 ( 
.A1(n_845),
.A2(n_601),
.B1(n_756),
.B2(n_752),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_843),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_918),
.B(n_812),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_892),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_847),
.B(n_493),
.Y(n_928)
);

INVxp33_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_SL g930 ( 
.A1(n_840),
.A2(n_755),
.B1(n_781),
.B2(n_750),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_845),
.A2(n_625),
.B1(n_604),
.B2(n_528),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_841),
.B(n_497),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_841),
.B(n_534),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_840),
.A2(n_542),
.B(n_546),
.C(n_540),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_918),
.B(n_812),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_903),
.B(n_550),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_890),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_846),
.B(n_851),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_856),
.B(n_543),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_903),
.B(n_558),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_865),
.B(n_518),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_842),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_885),
.B(n_559),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_885),
.B(n_865),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_852),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_908),
.B(n_524),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_848),
.B(n_561),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_876),
.B(n_821),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_848),
.B(n_566),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_846),
.B(n_862),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_905),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_846),
.B(n_570),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_906),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_911),
.B(n_908),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_875),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_899),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_893),
.A2(n_772),
.B1(n_583),
.B2(n_587),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_872),
.B(n_579),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_893),
.A2(n_598),
.B1(n_599),
.B2(n_594),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_868),
.B(n_544),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_899),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_882),
.B(n_602),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_890),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_899),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_874),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_886),
.B(n_611),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_880),
.B(n_747),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_873),
.B(n_896),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_L g971 ( 
.A(n_861),
.B(n_530),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_894),
.B(n_614),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_890),
.B(n_748),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_898),
.B(n_616),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_857),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_900),
.B(n_621),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_863),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_858),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_864),
.B(n_627),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_877),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_873),
.B(n_896),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_897),
.B(n_628),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_912),
.A2(n_649),
.B(n_636),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_901),
.B(n_650),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_869),
.A2(n_549),
.B1(n_551),
.B2(n_545),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_526),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_858),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_555),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_859),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_919),
.B(n_867),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_910),
.B(n_755),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_855),
.B(n_749),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_914),
.B(n_660),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_863),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_877),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_891),
.B(n_569),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_878),
.Y(n_997)
);

AND3x1_ASAP7_75t_L g998 ( 
.A(n_849),
.B(n_761),
.C(n_754),
.Y(n_998)
);

NAND2x1_ASAP7_75t_L g999 ( 
.A(n_917),
.B(n_681),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_910),
.B(n_552),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_887),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_895),
.A2(n_560),
.B1(n_568),
.B2(n_565),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_L g1003 ( 
.A(n_895),
.B(n_530),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_888),
.B(n_902),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_888),
.B(n_664),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_878),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_870),
.B(n_571),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_870),
.B(n_575),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_913),
.B(n_671),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_879),
.B(n_652),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_870),
.B(n_576),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_879),
.B(n_708),
.C(n_701),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_859),
.B(n_691),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_878),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_893),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_889),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_907),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_889),
.B(n_692),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_875),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_907),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_870),
.B(n_580),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_915),
.A2(n_585),
.B1(n_588),
.B2(n_582),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_895),
.A2(n_916),
.B1(n_915),
.B2(n_917),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_844),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_916),
.A2(n_766),
.B(n_775),
.C(n_765),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_844),
.A2(n_778),
.B(n_779),
.C(n_777),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_850),
.B(n_590),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_850),
.A2(n_593),
.B1(n_595),
.B2(n_592),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_853),
.B(n_596),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_603),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_883),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_SL g1032 ( 
.A1(n_881),
.A2(n_708),
.B1(n_715),
.B2(n_701),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_881),
.B(n_605),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_895),
.A2(n_562),
.B1(n_530),
.B2(n_572),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_904),
.B(n_607),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_895),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_904),
.B(n_577),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_904),
.A2(n_562),
.B1(n_530),
.B2(n_620),
.Y(n_1038)
);

INVxp33_ASAP7_75t_L g1039 ( 
.A(n_883),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_909),
.A2(n_562),
.B1(n_530),
.B2(n_622),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_909),
.B(n_608),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_871),
.B(n_623),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_871),
.B(n_624),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_955),
.B(n_715),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_925),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_938),
.B(n_909),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_944),
.B(n_613),
.C(n_610),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_927),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_980),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_997),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_977),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_995),
.B(n_946),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_952),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_1006),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1010),
.B(n_723),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_924),
.A2(n_731),
.B(n_723),
.C(n_818),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_923),
.A2(n_618),
.B(n_617),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_938),
.B(n_826),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_973),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_970),
.B(n_883),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_956),
.B(n_562),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_956),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_956),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_956),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_932),
.A2(n_562),
.B1(n_629),
.B2(n_573),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_994),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_1020),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_957),
.B(n_883),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_921),
.B(n_619),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_946),
.B(n_633),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_1017),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_1014),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_933),
.B(n_638),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_920),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1001),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_1012),
.B(n_1032),
.C(n_924),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_1024),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_964),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_975),
.Y(n_1079)
);

OR2x6_ASAP7_75t_SL g1080 ( 
.A(n_931),
.B(n_626),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_929),
.B(n_731),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1024),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_978),
.Y(n_1083)
);

BUFx10_ASAP7_75t_L g1084 ( 
.A(n_941),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_970),
.B(n_637),
.C(n_630),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_981),
.B(n_651),
.C(n_645),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_962),
.B(n_184),
.Y(n_1087)
);

AO221x1_ASAP7_75t_L g1088 ( 
.A1(n_1019),
.A2(n_678),
.B1(n_629),
.B2(n_573),
.C(n_659),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_973),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_981),
.B(n_640),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_987),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_941),
.B(n_996),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_991),
.B(n_573),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_945),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_996),
.B(n_928),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_942),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1036),
.Y(n_1097)
);

NOR2x1p5_ASAP7_75t_L g1098 ( 
.A(n_966),
.B(n_657),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1015),
.B(n_562),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_948),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_967),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_SL g1102 ( 
.A(n_930),
.B(n_668),
.C(n_665),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_939),
.B(n_670),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_SL g1105 ( 
.A(n_990),
.B(n_675),
.C(n_673),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_937),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_922),
.B(n_682),
.C(n_677),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_937),
.B(n_187),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1016),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_954),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_965),
.B(n_969),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_926),
.B(n_629),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_986),
.B(n_644),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_947),
.B(n_562),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_951),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_950),
.B(n_646),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_998),
.B(n_678),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1000),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_984),
.B(n_647),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_935),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_961),
.B(n_648),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_953),
.B(n_188),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1031),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1004),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_999),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_986),
.B(n_678),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_940),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_985),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_959),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_963),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1041),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_988),
.B(n_654),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_992),
.B(n_189),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_988),
.B(n_656),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_968),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_972),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_949),
.B(n_1043),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_982),
.B(n_661),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_974),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_976),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1042),
.B(n_662),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1037),
.B(n_669),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1042),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1009),
.Y(n_1145)
);

INVx4_ASAP7_75t_SL g1146 ( 
.A(n_960),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1037),
.B(n_676),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1043),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_971),
.B(n_679),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1039),
.B(n_680),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1013),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_943),
.B(n_684),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1025),
.B(n_190),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_934),
.A2(n_689),
.B(n_690),
.C(n_685),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1005),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1018),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_979),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_1026),
.B(n_6),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_993),
.Y(n_1159)
);

OR2x2_ASAP7_75t_SL g1160 ( 
.A(n_1033),
.B(n_8),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1027),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1028),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1029),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1023),
.B(n_1002),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_1003),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1030),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1023),
.B(n_693),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1035),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1007),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1022),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_983),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_958),
.B(n_191),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_958),
.A2(n_197),
.B1(n_198),
.B2(n_194),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_1040),
.B(n_9),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_960),
.B(n_200),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1008),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_SL g1177 ( 
.A(n_1011),
.B(n_10),
.C(n_11),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1021),
.B(n_205),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1038),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1038),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1040),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1034),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_952),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_1012),
.B(n_10),
.C(n_12),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_977),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_955),
.B(n_13),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_977),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_956),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_956),
.B(n_206),
.Y(n_1190)
);

CKINVDCx6p67_ASAP7_75t_R g1191 ( 
.A(n_1017),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_921),
.B(n_13),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_930),
.B(n_14),
.C(n_15),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_921),
.B(n_14),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_927),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_927),
.B(n_15),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_927),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_995),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_927),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_921),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_995),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_956),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_952),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_921),
.B(n_208),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_955),
.B(n_16),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1004),
.A2(n_486),
.B(n_213),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_927),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_921),
.B(n_209),
.Y(n_1208)
);

AND2x6_ASAP7_75t_SL g1209 ( 
.A(n_991),
.B(n_17),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_925),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_956),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_921),
.B(n_18),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_921),
.B(n_215),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_977),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_R g1215 ( 
.A(n_995),
.B(n_216),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_921),
.B(n_217),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_927),
.B(n_19),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_956),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_977),
.Y(n_1219)
);

BUFx4f_ASAP7_75t_SL g1220 ( 
.A(n_1017),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_980),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1114),
.A2(n_220),
.B(n_218),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1092),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1204),
.A2(n_222),
.B(n_221),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1052),
.B(n_20),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1049),
.B(n_21),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1062),
.Y(n_1227)
);

NOR4xp25_ASAP7_75t_L g1228 ( 
.A(n_1193),
.B(n_24),
.C(n_22),
.D(n_23),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1062),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1159),
.B(n_23),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1204),
.A2(n_225),
.B(n_224),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1208),
.A2(n_227),
.B(n_226),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1095),
.A2(n_229),
.B(n_228),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1208),
.A2(n_233),
.B(n_231),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1213),
.A2(n_236),
.B(n_234),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1213),
.A2(n_238),
.B(n_237),
.Y(n_1236)
);

AND3x4_ASAP7_75t_L g1237 ( 
.A(n_1058),
.B(n_26),
.C(n_27),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1197),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1099),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1124),
.B(n_26),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1115),
.B(n_1090),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1094),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1128),
.B(n_27),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1046),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1114),
.A2(n_1216),
.B(n_1060),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1110),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1216),
.A2(n_244),
.B(n_242),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1109),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1161),
.B(n_28),
.Y(n_1250)
);

NOR2xp67_ASAP7_75t_L g1251 ( 
.A(n_1053),
.B(n_1067),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1099),
.A2(n_1206),
.B(n_1082),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1192),
.A2(n_28),
.B(n_29),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_1081),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1049),
.B(n_30),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1163),
.B(n_30),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1077),
.A2(n_248),
.B(n_245),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1135),
.B(n_31),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1051),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1165),
.A2(n_251),
.B(n_250),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1070),
.B(n_32),
.Y(n_1261)
);

NOR2x1_ASAP7_75t_SL g1262 ( 
.A(n_1165),
.B(n_252),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1184),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1155),
.B(n_32),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1077),
.A2(n_254),
.B(n_253),
.Y(n_1265)
);

AND2x6_ASAP7_75t_L g1266 ( 
.A(n_1175),
.B(n_257),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1183),
.A2(n_1194),
.A3(n_1212),
.B(n_1181),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1131),
.B(n_33),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1066),
.Y(n_1269)
);

OAI22x1_ASAP7_75t_L g1270 ( 
.A1(n_1074),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1165),
.A2(n_260),
.B(n_258),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1082),
.A2(n_1123),
.B(n_1171),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1084),
.B(n_261),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1137),
.B(n_35),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1075),
.A2(n_265),
.B(n_262),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1164),
.A2(n_268),
.B(n_266),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1183),
.A2(n_38),
.A3(n_36),
.B(n_37),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1111),
.B(n_272),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1063),
.A2(n_275),
.B(n_274),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1157),
.B(n_38),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1116),
.A2(n_1167),
.B(n_1047),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1157),
.B(n_39),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1091),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1207),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1084),
.B(n_39),
.Y(n_1285)
);

OAI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1174),
.A2(n_40),
.B(n_41),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1048),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1186),
.A2(n_279),
.B(n_278),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1188),
.A2(n_282),
.B(n_281),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1182),
.A2(n_286),
.B(n_284),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1175),
.B(n_40),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1055),
.B(n_41),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1198),
.B(n_42),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1146),
.B(n_42),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1214),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1219),
.A2(n_289),
.B(n_287),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1044),
.B(n_43),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1045),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1195),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1187),
.A2(n_45),
.A3(n_43),
.B(n_44),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1205),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1091),
.Y(n_1302)
);

OA22x2_ASAP7_75t_L g1303 ( 
.A1(n_1112),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_1203),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1116),
.A2(n_49),
.A3(n_47),
.B(n_48),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1064),
.A2(n_292),
.B(n_291),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1146),
.B(n_49),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1138),
.B(n_50),
.Y(n_1308)
);

OA22x2_ASAP7_75t_L g1309 ( 
.A1(n_1112),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1167),
.A2(n_294),
.B(n_293),
.Y(n_1310)
);

AOI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1153),
.A2(n_52),
.B(n_53),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1064),
.A2(n_297),
.B(n_296),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1151),
.B(n_53),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1058),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1156),
.B(n_54),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1072),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1111),
.B(n_299),
.Y(n_1317)
);

INVx5_ASAP7_75t_L g1318 ( 
.A(n_1062),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1063),
.A2(n_305),
.B(n_301),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1078),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_309),
.B1(n_313),
.B2(n_307),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1047),
.A2(n_316),
.B(n_314),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1218),
.A2(n_318),
.B(n_317),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1127),
.B(n_54),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1130),
.B(n_55),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1202),
.A2(n_322),
.B(n_319),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1079),
.A2(n_324),
.B(n_323),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1218),
.A2(n_326),
.B(n_325),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1140),
.B(n_55),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1211),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1218),
.A2(n_328),
.B(n_327),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1142),
.B(n_56),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1083),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1104),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1071),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1210),
.Y(n_1336)
);

AOI21xp33_ASAP7_75t_L g1337 ( 
.A1(n_1113),
.A2(n_56),
.B(n_57),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1179),
.A2(n_330),
.B(n_329),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1201),
.B(n_58),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_SL g1340 ( 
.A(n_1211),
.B(n_58),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1180),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1341)
);

INVx3_ASAP7_75t_SL g1342 ( 
.A(n_1191),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1168),
.A2(n_1190),
.B(n_1176),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1143),
.A2(n_337),
.B(n_336),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1136),
.B(n_60),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1179),
.B(n_61),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1119),
.B(n_62),
.Y(n_1347)
);

AO21x1_ASAP7_75t_L g1348 ( 
.A1(n_1172),
.A2(n_63),
.B(n_64),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1119),
.B(n_65),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1068),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1200),
.A2(n_67),
.A3(n_65),
.B(n_66),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1169),
.A2(n_342),
.B(n_340),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1068),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1102),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1147),
.A2(n_347),
.B(n_343),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1056),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1189),
.A2(n_349),
.B(n_348),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1152),
.A2(n_353),
.B(n_352),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1069),
.A2(n_355),
.B(n_354),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1133),
.A2(n_360),
.B(n_356),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1073),
.B(n_72),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1144),
.B(n_361),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1046),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1166),
.B(n_73),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1211),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1122),
.A2(n_363),
.B(n_362),
.Y(n_1366)
);

AOI221x1_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.C(n_76),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1154),
.A2(n_367),
.B(n_364),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_R g1369 ( 
.A(n_1221),
.B(n_368),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1141),
.B(n_1145),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1141),
.B(n_77),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1096),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1122),
.A2(n_373),
.B(n_369),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1061),
.A2(n_378),
.B(n_376),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1057),
.A2(n_381),
.B(n_380),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1199),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1170),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1377)
);

BUFx2_ASAP7_75t_SL g1378 ( 
.A(n_1101),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1145),
.B(n_80),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1057),
.A2(n_1098),
.B(n_1173),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1149),
.A2(n_387),
.B(n_383),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1098),
.A2(n_391),
.B(n_389),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1189),
.A2(n_394),
.B(n_393),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1173),
.A2(n_396),
.B(n_395),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1087),
.A2(n_398),
.B(n_397),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1125),
.Y(n_1386)
);

INVx6_ASAP7_75t_SL g1387 ( 
.A(n_1112),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1144),
.B(n_399),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1097),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_1118),
.B(n_400),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1139),
.A2(n_1121),
.B(n_1087),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1150),
.A2(n_81),
.A3(n_82),
.B(n_83),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1153),
.A2(n_405),
.B(n_402),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1244),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1241),
.B(n_1076),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1244),
.B(n_1089),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1348),
.A2(n_1106),
.A3(n_1080),
.B(n_1088),
.Y(n_1397)
);

BUFx2_ASAP7_75t_R g1398 ( 
.A(n_1342),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1272),
.A2(n_1103),
.B(n_1196),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1266),
.B(n_1129),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1304),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1239),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1363),
.B(n_1108),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1239),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1284),
.B(n_1162),
.Y(n_1405)
);

BUFx8_ASAP7_75t_L g1406 ( 
.A(n_1316),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1227),
.B(n_1097),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1281),
.A2(n_1134),
.B(n_1178),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1242),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1372),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1252),
.A2(n_1217),
.B(n_1117),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1308),
.B(n_1185),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1297),
.A2(n_1065),
.B1(n_1120),
.B2(n_1093),
.C(n_1105),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1295),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1367),
.A2(n_1085),
.A3(n_1086),
.B(n_1177),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1295),
.Y(n_1416)
);

BUFx2_ASAP7_75t_R g1417 ( 
.A(n_1263),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1335),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1262),
.A2(n_1059),
.B(n_1160),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1327),
.A2(n_1125),
.B(n_1132),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1352),
.A2(n_1125),
.B(n_1132),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1245),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1225),
.B(n_1108),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_1107),
.B(n_1134),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_R g1425 ( 
.A(n_1335),
.B(n_1178),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1247),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1227),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1292),
.B(n_1093),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1266),
.A2(n_1215),
.B1(n_1132),
.B2(n_1093),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1376),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1378),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1266),
.A2(n_1158),
.B1(n_1097),
.B2(n_1054),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1251),
.B(n_1158),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1369),
.Y(n_1434)
);

AO21x1_ASAP7_75t_L g1435 ( 
.A1(n_1258),
.A2(n_1158),
.B(n_1209),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1259),
.Y(n_1436)
);

OAI211xp5_ASAP7_75t_L g1437 ( 
.A1(n_1354),
.A2(n_1209),
.B(n_1054),
.C(n_1050),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1343),
.A2(n_1126),
.B(n_1050),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1266),
.A2(n_1126),
.B1(n_1220),
.B2(n_83),
.Y(n_1439)
);

AOI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1332),
.A2(n_1126),
.B(n_81),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1389),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1370),
.B(n_82),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1306),
.A2(n_411),
.B(n_410),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1269),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1291),
.A2(n_1261),
.B1(n_1324),
.B2(n_1307),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1298),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1391),
.B(n_84),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1353),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1353),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1310),
.A2(n_415),
.B(n_413),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1238),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1249),
.Y(n_1452)
);

BUFx2_ASAP7_75t_R g1453 ( 
.A(n_1294),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1298),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1337),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_1349),
.B1(n_1347),
.B2(n_1386),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1363),
.B(n_485),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1237),
.A2(n_1364),
.B1(n_1377),
.B2(n_1361),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1262),
.A2(n_418),
.B(n_416),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1312),
.A2(n_484),
.B(n_483),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1281),
.A2(n_482),
.B(n_481),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1314),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1375),
.A2(n_479),
.B(n_478),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1293),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1314),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1303),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1326),
.A2(n_1265),
.B(n_1257),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1309),
.A2(n_1345),
.B1(n_1346),
.B2(n_1256),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1290),
.A2(n_473),
.B(n_472),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1333),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1278),
.B(n_470),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1275),
.A2(n_1289),
.B(n_1288),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1320),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1278),
.B(n_419),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1334),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1254),
.B(n_93),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1285),
.A2(n_1317),
.B1(n_1390),
.B2(n_1250),
.Y(n_1477)
);

AO31x2_ASAP7_75t_L g1478 ( 
.A1(n_1223),
.A2(n_94),
.A3(n_95),
.B(n_96),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1368),
.A2(n_466),
.B(n_465),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1246),
.A2(n_462),
.B(n_460),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1296),
.A2(n_458),
.B(n_457),
.Y(n_1481)
);

AO31x2_ASAP7_75t_L g1482 ( 
.A1(n_1341),
.A2(n_95),
.A3(n_96),
.B(n_97),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1389),
.B(n_1287),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1264),
.B(n_98),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1299),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1389),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1336),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1224),
.A2(n_456),
.B(n_454),
.Y(n_1488)
);

CKINVDCx8_ASAP7_75t_R g1489 ( 
.A(n_1227),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1283),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1229),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1231),
.A2(n_448),
.B(n_447),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1302),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1317),
.B(n_421),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1356),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1229),
.Y(n_1496)
);

AO32x2_ASAP7_75t_L g1497 ( 
.A1(n_1228),
.A2(n_99),
.A3(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1232),
.A2(n_444),
.B(n_441),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1339),
.B(n_103),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1240),
.B(n_104),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1243),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1286),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1267),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1234),
.A2(n_440),
.B(n_439),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1267),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1235),
.A2(n_1248),
.B(n_1236),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1267),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1382),
.A2(n_436),
.B(n_432),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_L g1509 ( 
.A(n_1230),
.B(n_426),
.Y(n_1509)
);

AOI21xp33_ASAP7_75t_R g1510 ( 
.A1(n_1268),
.A2(n_105),
.B(n_107),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1233),
.A2(n_425),
.B(n_424),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_R g1512 ( 
.A(n_1318),
.B(n_422),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1365),
.B(n_423),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1229),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1384),
.A2(n_108),
.B(n_109),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1280),
.A2(n_108),
.B(n_109),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1276),
.A2(n_110),
.B(n_111),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1274),
.A2(n_1313),
.B1(n_1315),
.B2(n_1371),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1393),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1379),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1365),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1318),
.B(n_112),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1387),
.Y(n_1524)
);

BUFx2_ASAP7_75t_R g1525 ( 
.A(n_1381),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1226),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1255),
.B(n_114),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1282),
.A2(n_114),
.B(n_115),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1301),
.B(n_115),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1393),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1338),
.A2(n_116),
.B(n_117),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1270),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1273),
.B(n_119),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1318),
.B(n_122),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1277),
.Y(n_1535)
);

BUFx10_ASAP7_75t_L g1536 ( 
.A(n_1387),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1321),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1395),
.B(n_1423),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1418),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1484),
.A2(n_1340),
.B1(n_1366),
.B2(n_1373),
.C(n_1362),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1523),
.B(n_1388),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1458),
.A2(n_1330),
.B1(n_1385),
.B2(n_1360),
.Y(n_1542)
);

BUFx4f_ASAP7_75t_SL g1543 ( 
.A(n_1406),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1439),
.B(n_1322),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1330),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1410),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1403),
.B(n_1330),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1447),
.A2(n_1344),
.B1(n_1355),
.B2(n_1358),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1451),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1516),
.A2(n_1359),
.B1(n_1383),
.B2(n_1374),
.C(n_1271),
.Y(n_1550)
);

AOI22x1_ASAP7_75t_L g1551 ( 
.A1(n_1515),
.A2(n_1260),
.B1(n_1279),
.B2(n_1323),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1435),
.A2(n_1322),
.B1(n_1222),
.B2(n_1319),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1477),
.A2(n_1328),
.B1(n_1331),
.B2(n_1222),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1418),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_SL g1555 ( 
.A(n_1398),
.B(n_1417),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1445),
.B(n_1468),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1418),
.B(n_1311),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1518),
.A2(n_1357),
.B1(n_1253),
.B2(n_1351),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1413),
.A2(n_1351),
.B(n_1305),
.C(n_1392),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1427),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1396),
.B(n_1300),
.Y(n_1561)
);

NAND2xp33_ASAP7_75t_SL g1562 ( 
.A(n_1401),
.B(n_1300),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1467),
.A2(n_1305),
.B(n_1277),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1396),
.B(n_1277),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1537),
.A2(n_1392),
.B1(n_1305),
.B2(n_125),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1412),
.B(n_1392),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1528),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1471),
.B(n_126),
.Y(n_1568)
);

AO31x2_ASAP7_75t_L g1569 ( 
.A1(n_1535),
.A2(n_127),
.A3(n_128),
.B(n_129),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1414),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1440),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1414),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1499),
.B(n_130),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1416),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1529),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1429),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1427),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1430),
.Y(n_1578)
);

OAI222xp33_ASAP7_75t_L g1579 ( 
.A1(n_1532),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.C1(n_137),
.C2(n_139),
.Y(n_1579)
);

AO32x2_ASAP7_75t_L g1580 ( 
.A1(n_1456),
.A2(n_136),
.A3(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_1580)
);

INVx4_ASAP7_75t_SL g1581 ( 
.A(n_1534),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1510),
.A2(n_1495),
.B1(n_1455),
.B2(n_1502),
.C(n_1466),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1489),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1485),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1433),
.A2(n_1526),
.B1(n_1500),
.B2(n_1520),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1471),
.B(n_1474),
.Y(n_1586)
);

AND2x6_ASAP7_75t_L g1587 ( 
.A(n_1402),
.B(n_140),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1464),
.B(n_1400),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1422),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1422),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1434),
.Y(n_1591)
);

AO31x2_ASAP7_75t_L g1592 ( 
.A1(n_1535),
.A2(n_142),
.A3(n_144),
.B(n_145),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1444),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1420),
.A2(n_142),
.B(n_144),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1409),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1527),
.B(n_146),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1405),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1474),
.B(n_147),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1426),
.B(n_148),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1486),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1433),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_R g1602 ( 
.A(n_1524),
.B(n_149),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1450),
.A2(n_181),
.B(n_154),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1444),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1436),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1494),
.B(n_153),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1494),
.B(n_154),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1428),
.B(n_155),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1402),
.B(n_155),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1419),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1452),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1454),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1470),
.B(n_160),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1533),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1431),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1536),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1469),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_1617)
);

OAI211xp5_ASAP7_75t_L g1618 ( 
.A1(n_1437),
.A2(n_166),
.B(n_167),
.C(n_168),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1457),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1476),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1473),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1522),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1469),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_1623)
);

AND2x6_ASAP7_75t_L g1624 ( 
.A(n_1404),
.B(n_172),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1531),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1425),
.B(n_176),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1487),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1493),
.B(n_176),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1450),
.A2(n_177),
.B(n_178),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1503),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1454),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1453),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1442),
.B(n_1475),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1475),
.B(n_179),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1407),
.B(n_180),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1448),
.A2(n_180),
.B1(n_1449),
.B2(n_1432),
.C(n_1446),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1490),
.B(n_1415),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1490),
.B(n_1415),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1538),
.B(n_1483),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1567),
.A2(n_1531),
.B1(n_1511),
.B2(n_1517),
.Y(n_1640)
);

AOI21xp33_ASAP7_75t_L g1641 ( 
.A1(n_1556),
.A2(n_1424),
.B(n_1511),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1582),
.A2(n_1424),
.B1(n_1509),
.B2(n_1534),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1581),
.B(n_1491),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1620),
.A2(n_1461),
.B1(n_1480),
.B2(n_1459),
.C(n_1505),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1546),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1597),
.A2(n_1457),
.B1(n_1513),
.B2(n_1462),
.Y(n_1646)
);

OAI211xp5_ASAP7_75t_L g1647 ( 
.A1(n_1601),
.A2(n_1497),
.B(n_1408),
.C(n_1512),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_L g1648 ( 
.A(n_1540),
.B(n_1399),
.C(n_1411),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1541),
.B(n_1397),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1576),
.A2(n_1465),
.B1(n_1394),
.B2(n_1463),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1585),
.A2(n_1394),
.B1(n_1521),
.B2(n_1441),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1636),
.A2(n_1463),
.B1(n_1507),
.B2(n_1505),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1591),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1544),
.A2(n_1622),
.B1(n_1618),
.B2(n_1624),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1581),
.B(n_1514),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1571),
.A2(n_1503),
.B1(n_1479),
.B2(n_1441),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1614),
.A2(n_1497),
.B(n_1479),
.C(n_1530),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1566),
.B(n_1397),
.Y(n_1658)
);

AO21x1_ASAP7_75t_L g1659 ( 
.A1(n_1562),
.A2(n_1530),
.B(n_1519),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1575),
.A2(n_1525),
.B1(n_1497),
.B2(n_1519),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1587),
.A2(n_1441),
.B1(n_1508),
.B2(n_1496),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1563),
.A2(n_1506),
.B(n_1472),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1586),
.A2(n_1438),
.B1(n_1496),
.B2(n_1481),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1635),
.A2(n_1496),
.B1(n_1482),
.B2(n_1478),
.Y(n_1664)
);

AOI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1542),
.A2(n_1548),
.B(n_1558),
.Y(n_1665)
);

OAI211xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1626),
.A2(n_1607),
.B(n_1606),
.C(n_1588),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1549),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1587),
.A2(n_1504),
.B1(n_1492),
.B2(n_1498),
.Y(n_1668)
);

AND2x6_ASAP7_75t_SL g1669 ( 
.A(n_1635),
.B(n_1482),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1617),
.A2(n_1478),
.B1(n_1421),
.B2(n_1443),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1608),
.B(n_1488),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1595),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1633),
.B(n_1460),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1579),
.A2(n_1565),
.B1(n_1623),
.B2(n_1559),
.C(n_1625),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1587),
.A2(n_1624),
.B1(n_1598),
.B2(n_1568),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1550),
.A2(n_1610),
.B1(n_1551),
.B2(n_1553),
.C(n_1552),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1587),
.A2(n_1624),
.B1(n_1598),
.B2(n_1568),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1573),
.B(n_1613),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1586),
.A2(n_1578),
.B1(n_1609),
.B2(n_1634),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1589),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1624),
.A2(n_1561),
.B1(n_1619),
.B2(n_1564),
.Y(n_1681)
);

AO31x2_ASAP7_75t_L g1682 ( 
.A1(n_1630),
.A2(n_1603),
.A3(n_1629),
.B(n_1637),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1555),
.A2(n_1632),
.B1(n_1545),
.B2(n_1543),
.Y(n_1683)
);

OAI21xp33_ASAP7_75t_L g1684 ( 
.A1(n_1599),
.A2(n_1628),
.B(n_1596),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_SL g1685 ( 
.A1(n_1638),
.A2(n_1590),
.B(n_1593),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1551),
.A2(n_1557),
.B1(n_1564),
.B2(n_1554),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1621),
.B(n_1627),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1584),
.A2(n_1616),
.B1(n_1615),
.B2(n_1611),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1605),
.A2(n_1583),
.B1(n_1547),
.B2(n_1600),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1583),
.A2(n_1547),
.B1(n_1539),
.B2(n_1604),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1583),
.A2(n_1539),
.B1(n_1631),
.B2(n_1612),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1570),
.A2(n_1572),
.B(n_1574),
.Y(n_1692)
);

INVx3_ASAP7_75t_SL g1693 ( 
.A(n_1577),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1630),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1594),
.A2(n_1560),
.B(n_1580),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1580),
.A2(n_1577),
.B1(n_1569),
.B2(n_1592),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1577),
.A2(n_1092),
.B1(n_946),
.B2(n_1458),
.C(n_930),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1580),
.A2(n_1297),
.B1(n_1567),
.B2(n_1102),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1658),
.B(n_1569),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1694),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1666),
.B(n_1592),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1662),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1680),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1649),
.B(n_1682),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1682),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1696),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1676),
.A2(n_1665),
.B(n_1648),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1645),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1639),
.B(n_1678),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1697),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1698),
.A2(n_1674),
.B1(n_1660),
.B2(n_1654),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1696),
.B(n_1697),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1641),
.B(n_1659),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1663),
.B(n_1671),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1660),
.A2(n_1699),
.B1(n_1684),
.B2(n_1679),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1679),
.B(n_1673),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1667),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1692),
.B(n_1664),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1640),
.B(n_1681),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1669),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1687),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1670),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1647),
.B(n_1657),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1686),
.B(n_1668),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1652),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1703),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1701),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1713),
.A2(n_1646),
.B1(n_1651),
.B2(n_1677),
.Y(n_1731)
);

OAI321xp33_ASAP7_75t_L g1732 ( 
.A1(n_1713),
.A2(n_1642),
.A3(n_1675),
.B1(n_1691),
.B2(n_1650),
.C(n_1644),
.Y(n_1732)
);

OAI321xp33_ASAP7_75t_L g1733 ( 
.A1(n_1726),
.A2(n_1661),
.A3(n_1656),
.B1(n_1690),
.B2(n_1688),
.C(n_1689),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1700),
.B(n_1714),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1693),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1710),
.B(n_1683),
.Y(n_1736)
);

AOI31xp33_ASAP7_75t_L g1737 ( 
.A1(n_1717),
.A2(n_1695),
.A3(n_1643),
.B(n_1655),
.Y(n_1737)
);

OAI31xp33_ASAP7_75t_L g1738 ( 
.A1(n_1709),
.A2(n_1643),
.A3(n_1653),
.B(n_1726),
.Y(n_1738)
);

AOI31xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1709),
.A2(n_1702),
.A3(n_1721),
.B(n_1719),
.Y(n_1739)
);

AO21x2_ASAP7_75t_L g1740 ( 
.A1(n_1707),
.A2(n_1715),
.B(n_1714),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

NOR4xp25_ASAP7_75t_SL g1742 ( 
.A(n_1728),
.B(n_1712),
.C(n_1723),
.D(n_1718),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1714),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1725),
.A2(n_1723),
.B1(n_1728),
.B2(n_1708),
.C(n_1715),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1704),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1710),
.B(n_1724),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1734),
.B(n_1705),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1730),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1745),
.B(n_1716),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1745),
.B(n_1716),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1740),
.B(n_1719),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1746),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1746),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1716),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1736),
.B(n_1711),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1743),
.B(n_1716),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1730),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1729),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1743),
.B(n_1723),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1730),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1723),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1729),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1735),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1762),
.B(n_1740),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1762),
.B(n_1740),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1754),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1756),
.B(n_1738),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1764),
.B(n_1720),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1761),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1764),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1765),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1769),
.A2(n_1739),
.B1(n_1738),
.B2(n_1744),
.C(n_1731),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1769),
.B(n_1760),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1760),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1773),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1776),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1774),
.B(n_1775),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1776),
.B(n_1764),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1775),
.A2(n_1732),
.B1(n_1733),
.B2(n_1725),
.C1(n_1722),
.C2(n_1766),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1782),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1731),
.C(n_1742),
.Y(n_1785)
);

AOI222xp33_ASAP7_75t_L g1786 ( 
.A1(n_1779),
.A2(n_1767),
.B1(n_1766),
.B2(n_1722),
.C1(n_1739),
.C2(n_1727),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1784),
.Y(n_1787)
);

XNOR2x2_ASAP7_75t_L g1788 ( 
.A(n_1785),
.B(n_1778),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1787),
.B(n_1781),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1789),
.A2(n_1788),
.B(n_1786),
.C(n_1783),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1790),
.Y(n_1791)
);

XNOR2xp5_ASAP7_75t_L g1792 ( 
.A(n_1790),
.B(n_1720),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1791),
.B(n_1767),
.Y(n_1793)
);

AOI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1792),
.A2(n_1752),
.B(n_1727),
.C(n_1735),
.Y(n_1794)
);

A2O1A1Ixp33_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1752),
.B(n_1737),
.C(n_1771),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1793),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1796),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1797),
.A2(n_1770),
.B1(n_1715),
.B2(n_1727),
.C(n_1722),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1795),
.Y(n_1800)
);

AO211x2_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1748),
.B(n_1747),
.C(n_1742),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1798),
.Y(n_1802)
);

XNOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1799),
.B(n_1721),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1798),
.Y(n_1804)
);

AO221x1_ASAP7_75t_L g1805 ( 
.A1(n_1798),
.A2(n_1763),
.B1(n_1759),
.B2(n_1729),
.C(n_1761),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1798),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1802),
.A2(n_1748),
.B(n_1750),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1804),
.A2(n_1763),
.B1(n_1759),
.B2(n_1749),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1806),
.A2(n_1763),
.B1(n_1759),
.B2(n_1749),
.Y(n_1809)
);

NOR2xp67_ASAP7_75t_L g1810 ( 
.A(n_1801),
.B(n_1763),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1803),
.A2(n_1750),
.B(n_1751),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1812),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1810),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1813),
.A2(n_1808),
.B1(n_1809),
.B2(n_1807),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1814),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1815),
.A2(n_1811),
.B1(n_1759),
.B2(n_1755),
.C(n_1757),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1817),
.A2(n_1816),
.B1(n_1757),
.B2(n_1755),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1706),
.B1(n_1749),
.B2(n_1758),
.C(n_1729),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1751),
.B(n_1706),
.C(n_1741),
.Y(n_1820)
);


endmodule