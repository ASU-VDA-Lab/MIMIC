module fake_jpeg_13032_n_414 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_414);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_44),
.B(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_66),
.Y(n_92)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_72),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_74),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_21),
.B1(n_25),
.B2(n_33),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_42),
.B1(n_28),
.B2(n_40),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_121),
.B1(n_72),
.B2(n_77),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_103),
.B1(n_117),
.B2(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_35),
.B1(n_28),
.B2(n_25),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_44),
.A2(n_40),
.B1(n_33),
.B2(n_26),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_119),
.B1(n_72),
.B2(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_118),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_50),
.A2(n_29),
.B1(n_23),
.B2(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_47),
.B(n_32),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_40),
.B1(n_33),
.B2(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_48),
.A2(n_36),
.B1(n_29),
.B2(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_52),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_121)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_142),
.B1(n_64),
.B2(n_81),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_74),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_74),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_55),
.B1(n_63),
.B2(n_75),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_165)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_72),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_143),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_67),
.B1(n_69),
.B2(n_46),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_77),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_58),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_53),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_71),
.C(n_78),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_104),
.C(n_85),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_100),
.B(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_26),
.B1(n_85),
.B2(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_26),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_160),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_181),
.B1(n_183),
.B2(n_185),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_114),
.B1(n_110),
.B2(n_89),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_89),
.B(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_128),
.B1(n_158),
.B2(n_125),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_68),
.B1(n_95),
.B2(n_93),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_128),
.A2(n_122),
.B1(n_93),
.B2(n_95),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_122),
.B1(n_98),
.B2(n_102),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_124),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_131),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_135),
.A2(n_122),
.B1(n_102),
.B2(n_84),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_131),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_138),
.B1(n_143),
.B2(n_146),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_102),
.B1(n_96),
.B2(n_83),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_196),
.Y(n_240)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_185),
.B1(n_180),
.B2(n_176),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_170),
.B(n_165),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_137),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_203),
.C(n_150),
.Y(n_244)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_153),
.C(n_137),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_127),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_207),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_187),
.B1(n_174),
.B2(n_164),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_184),
.B1(n_190),
.B2(n_175),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_171),
.B(n_132),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_215),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_147),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_217),
.B(n_169),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_134),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_145),
.B1(n_156),
.B2(n_140),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_220),
.B1(n_183),
.B2(n_173),
.Y(n_233)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_126),
.B1(n_133),
.B2(n_148),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_223),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_238),
.B1(n_239),
.B2(n_245),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_215),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_216),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_236),
.B1(n_242),
.B2(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_165),
.B1(n_186),
.B2(n_192),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_170),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_244),
.C(n_203),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_170),
.B1(n_167),
.B2(n_180),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_170),
.B1(n_176),
.B2(n_182),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_195),
.A2(n_178),
.B1(n_182),
.B2(n_124),
.Y(n_242)
);

AOI22x1_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_190),
.B1(n_114),
.B2(n_110),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_248),
.B(n_218),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_184),
.B1(n_162),
.B2(n_148),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_196),
.A2(n_184),
.B1(n_116),
.B2(n_83),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_149),
.B1(n_116),
.B2(n_161),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.C(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_201),
.C(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_256),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_214),
.C(n_198),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_262),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_211),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_260),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_217),
.C(n_200),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_263),
.C(n_270),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_208),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_209),
.C(n_212),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_264),
.B(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_268),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_235),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_234),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_235),
.B(n_243),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_221),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_219),
.B1(n_194),
.B2(n_202),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_227),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_166),
.B1(n_161),
.B2(n_157),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_166),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_91),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_91),
.B1(n_65),
.B2(n_123),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_31),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_239),
.C(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_31),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_279),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_233),
.B1(n_242),
.B2(n_247),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_284),
.A2(n_259),
.B1(n_272),
.B2(n_271),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_248),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_288),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_286),
.B(n_301),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_243),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_234),
.C(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_290),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_249),
.C(n_225),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_225),
.C(n_223),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_295),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_241),
.B1(n_250),
.B2(n_27),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_241),
.B1(n_250),
.B2(n_27),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_76),
.C(n_51),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_27),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_300),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_22),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_14),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_51),
.C(n_22),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_268),
.B(n_256),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_311),
.A2(n_301),
.B(n_2),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_327),
.B1(n_37),
.B2(n_3),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_277),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_320),
.B1(n_1),
.B2(n_2),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_288),
.B(n_305),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_5),
.B(n_6),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_291),
.A2(n_280),
.B1(n_279),
.B2(n_276),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_22),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_0),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_323),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_14),
.B(n_19),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_299),
.B(n_14),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_37),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_37),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_295),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_1),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_284),
.A3(n_290),
.B1(n_286),
.B2(n_300),
.C1(n_283),
.C2(n_281),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_330),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_333),
.A2(n_344),
.B1(n_314),
.B2(n_323),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_281),
.C(n_283),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_339),
.C(n_343),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_338),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_337),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_33),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_37),
.C(n_3),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_2),
.C(n_3),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_4),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_349),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_5),
.C(n_6),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_343),
.C(n_349),
.Y(n_359)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_334),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_357),
.A2(n_358),
.B(n_361),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_340),
.A2(n_317),
.B(n_316),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_362),
.Y(n_368)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_365),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_317),
.B(n_320),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_321),
.C(n_328),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_345),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_335),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_364),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_361),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_373),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_341),
.C(n_337),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_325),
.C(n_7),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_353),
.A2(n_318),
.B1(n_350),
.B2(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_375),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_351),
.A2(n_347),
.B1(n_325),
.B2(n_339),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_376),
.A2(n_363),
.B(n_362),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_319),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_379),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_319),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_368),
.B(n_354),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_384),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_382),
.A2(n_383),
.B(n_386),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_370),
.A2(n_359),
.B(n_363),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_379),
.B(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_364),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_388),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_6),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_369),
.B(n_372),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_376),
.B(n_377),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_399),
.B(n_8),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_367),
.C(n_7),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_397),
.Y(n_404)
);

NOR2x1p5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_7),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_9),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_8),
.B(n_9),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_380),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_401),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_8),
.C(n_9),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_404),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_405),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_406),
.A2(n_407),
.B(n_401),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_402),
.A2(n_393),
.B(n_398),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_410),
.Y(n_412)
);

OAI321xp33_ASAP7_75t_L g411 ( 
.A1(n_408),
.A2(n_400),
.A3(n_409),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_411)
);

AOI221xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_411),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_9),
.Y(n_414)
);


endmodule