module real_aes_7640_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_0), .A2(n_11), .B1(n_177), .B2(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_0), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_1), .Y(n_145) );
AOI21xp33_ASAP7_75t_L g294 ( .A1(n_2), .A2(n_217), .B(n_295), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g117 ( .A1(n_3), .A2(n_28), .B1(n_118), .B2(n_122), .C(n_127), .Y(n_117) );
INVx1_ASAP7_75t_L g202 ( .A(n_4), .Y(n_202) );
AND2x6_ASAP7_75t_L g222 ( .A(n_4), .B(n_200), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_4), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_5), .A2(n_216), .B(n_223), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_6), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g300 ( .A(n_7), .Y(n_300) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_8), .A2(n_22), .B1(n_91), .B2(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g214 ( .A(n_9), .Y(n_214) );
INVx1_ASAP7_75t_L g233 ( .A(n_10), .Y(n_233) );
INVx1_ASAP7_75t_L g178 ( .A(n_11), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_12), .A2(n_176), .B1(n_179), .B2(n_180), .Y(n_175) );
INVx1_ASAP7_75t_L g179 ( .A(n_12), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_12), .B(n_250), .Y(n_266) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_13), .A2(n_24), .B1(n_91), .B2(n_92), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_14), .B(n_217), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_15), .B(n_293), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_16), .A2(n_230), .B(n_232), .C(n_234), .Y(n_229) );
AOI22xp5_ASAP7_75t_SL g516 ( .A1(n_16), .A2(n_81), .B1(n_82), .B2(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_16), .Y(n_517) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_17), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_18), .B(n_265), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g137 ( .A1(n_19), .A2(n_26), .B1(n_138), .B2(n_142), .C(n_144), .Y(n_137) );
INVx1_ASAP7_75t_L g312 ( .A(n_20), .Y(n_312) );
INVx2_ASAP7_75t_L g220 ( .A(n_21), .Y(n_220) );
AOI222xp33_ASAP7_75t_L g157 ( .A1(n_23), .A2(n_29), .B1(n_33), .B2(n_158), .C1(n_160), .C2(n_166), .Y(n_157) );
OAI221xp5_ASAP7_75t_L g193 ( .A1(n_24), .A2(n_42), .B1(n_50), .B2(n_194), .C(n_195), .Y(n_193) );
INVxp67_ASAP7_75t_L g196 ( .A(n_24), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_25), .A2(n_222), .B(n_226), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g310 ( .A(n_27), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_30), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g131 ( .A(n_31), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_32), .Y(n_185) );
AOI221xp5_ASAP7_75t_L g84 ( .A1(n_34), .A2(n_52), .B1(n_85), .B2(n_102), .C(n_107), .Y(n_84) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_35), .A2(n_174), .B1(n_175), .B2(n_181), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_35), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_36), .A2(n_81), .B1(n_82), .B2(n_170), .Y(n_80) );
INVx1_ASAP7_75t_L g170 ( .A(n_36), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_37), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_38), .B(n_217), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_39), .A2(n_226), .B1(n_307), .B2(n_309), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_40), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_41), .Y(n_330) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_42), .A2(n_60), .B1(n_91), .B2(n_92), .Y(n_90) );
INVxp67_ASAP7_75t_L g197 ( .A(n_42), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_43), .A2(n_298), .B(n_299), .C(n_301), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_44), .Y(n_269) );
INVx1_ASAP7_75t_L g296 ( .A(n_45), .Y(n_296) );
INVx1_ASAP7_75t_L g200 ( .A(n_46), .Y(n_200) );
INVx1_ASAP7_75t_L g213 ( .A(n_47), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_48), .Y(n_194) );
AO22x1_ASAP7_75t_L g107 ( .A1(n_49), .A2(n_59), .B1(n_108), .B2(n_112), .Y(n_107) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_50), .A2(n_66), .B1(n_91), .B2(n_96), .Y(n_95) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_51), .A2(n_81), .B1(n_82), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_51), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_SL g320 ( .A1(n_53), .A2(n_250), .B(n_301), .C(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g322 ( .A(n_54), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_55), .Y(n_315) );
INVx1_ASAP7_75t_L g260 ( .A(n_56), .Y(n_260) );
INVx1_ASAP7_75t_L g188 ( .A(n_57), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_58), .A2(n_222), .B(n_226), .C(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_61), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g211 ( .A(n_62), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_63), .B(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_64), .A2(n_222), .B(n_226), .C(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g128 ( .A(n_65), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_67), .B(n_210), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_68), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_69), .A2(n_222), .B(n_226), .C(n_278), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_70), .Y(n_286) );
INVx1_ASAP7_75t_L g319 ( .A(n_71), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_72), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_73), .B(n_247), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_74), .Y(n_149) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_76), .B(n_238), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_77), .A2(n_217), .B(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_190), .B1(n_203), .B2(n_509), .C(n_515), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_171), .Y(n_79) );
INVx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AND4x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_117), .C(n_137), .D(n_157), .Y(n_83) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x6_ASAP7_75t_L g104 ( .A(n_88), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_L g159 ( .A(n_88), .B(n_154), .Y(n_159) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g111 ( .A(n_89), .B(n_95), .Y(n_111) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_90), .B(n_95), .Y(n_116) );
AND2x2_ASAP7_75t_L g125 ( .A(n_90), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g147 ( .A(n_90), .B(n_99), .Y(n_147) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g126 ( .A(n_95), .Y(n_126) );
INVx1_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
AND2x4_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g124 ( .A(n_97), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
OR2x2_ASAP7_75t_L g106 ( .A(n_98), .B(n_101), .Y(n_106) );
AND2x2_ASAP7_75t_L g121 ( .A(n_98), .B(n_101), .Y(n_121) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g154 ( .A(n_99), .B(n_101), .Y(n_154) );
INVx1_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
AND2x2_ASAP7_75t_L g164 ( .A(n_100), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx11_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g141 ( .A(n_105), .B(n_111), .Y(n_141) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x6_ASAP7_75t_L g143 ( .A(n_111), .B(n_121), .Y(n_143) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x6_ASAP7_75t_L g135 ( .A(n_116), .B(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx6_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_121), .B(n_125), .Y(n_130) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_131), .B2(n_132), .Y(n_127) );
BUFx2_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx6_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B1(n_149), .B2(n_150), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g168 ( .A(n_147), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
OR2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_165), .Y(n_169) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B1(n_182), .B2(n_183), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_175), .Y(n_181) );
INVx1_ASAP7_75t_L g180 ( .A(n_176), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_177), .A2(n_247), .B(n_333), .C(n_334), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_186), .B1(n_187), .B2(n_189), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_184), .Y(n_189) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
AND3x1_ASAP7_75t_SL g192 ( .A(n_193), .B(n_198), .C(n_201), .Y(n_192) );
INVxp67_ASAP7_75t_L g521 ( .A(n_193), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_SL g523 ( .A(n_198), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_198), .A2(n_526), .B(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g534 ( .A(n_198), .Y(n_534) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_199), .B(n_202), .Y(n_528) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_SL g533 ( .A(n_201), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
OR4x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_405), .C(n_464), .D(n_491), .Y(n_203) );
NAND3xp33_ASAP7_75t_SL g204 ( .A(n_205), .B(n_347), .C(n_372), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_271), .B(n_291), .C(n_324), .Y(n_205) );
AOI211xp5_ASAP7_75t_SL g495 ( .A1(n_206), .A2(n_496), .B(n_498), .C(n_501), .Y(n_495) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_240), .Y(n_206) );
INVx1_ASAP7_75t_L g370 ( .A(n_207), .Y(n_370) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g345 ( .A(n_208), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g377 ( .A(n_208), .Y(n_377) );
AND2x2_ASAP7_75t_L g432 ( .A(n_208), .B(n_401), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_208), .B(n_289), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_208), .B(n_290), .Y(n_490) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g351 ( .A(n_209), .Y(n_351) );
AND2x2_ASAP7_75t_L g394 ( .A(n_209), .B(n_258), .Y(n_394) );
AND2x2_ASAP7_75t_L g412 ( .A(n_209), .B(n_290), .Y(n_412) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_215), .B(n_237), .Y(n_209) );
INVx1_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
INVx2_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x2_ASAP7_75t_L g239 ( .A(n_211), .B(n_212), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_222), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_218), .B(n_222), .Y(n_261) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g514 ( .A(n_219), .Y(n_514) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
INVx1_ASAP7_75t_L g308 ( .A(n_220), .Y(n_308) );
INVx1_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
INVx3_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_221), .Y(n_250) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_221), .Y(n_265) );
INVx4_ASAP7_75t_SL g236 ( .A(n_222), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_229), .C(n_236), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_225), .A2(n_236), .B(n_296), .C(n_297), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_225), .A2(n_236), .B(n_319), .C(n_320), .Y(n_318) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
BUFx3_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_230), .B(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g309 ( .A1(n_231), .A2(n_310), .B1(n_311), .B2(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
OAI322xp33_ASAP7_75t_L g515 ( .A1(n_233), .A2(n_516), .A3(n_518), .B1(n_522), .B2(n_524), .C1(n_529), .C2(n_531), .Y(n_515) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g252 ( .A(n_235), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_236), .A2(n_261), .B1(n_306), .B2(n_313), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_236), .B(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g257 ( .A(n_238), .Y(n_257) );
OA21x2_ASAP7_75t_L g316 ( .A1(n_238), .A2(n_317), .B(n_323), .Y(n_316) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g254 ( .A(n_239), .Y(n_254) );
INVx4_ASAP7_75t_L g344 ( .A(n_240), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g399 ( .A1(n_240), .A2(n_400), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g480 ( .A(n_240), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_258), .Y(n_240) );
INVx1_ASAP7_75t_L g288 ( .A(n_241), .Y(n_288) );
AND2x2_ASAP7_75t_L g349 ( .A(n_241), .B(n_290), .Y(n_349) );
OR2x2_ASAP7_75t_L g378 ( .A(n_241), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g392 ( .A(n_241), .Y(n_392) );
INVx3_ASAP7_75t_L g401 ( .A(n_241), .Y(n_401) );
AND2x2_ASAP7_75t_L g411 ( .A(n_241), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g444 ( .A(n_241), .B(n_350), .Y(n_444) );
AND2x2_ASAP7_75t_L g468 ( .A(n_241), .B(n_424), .Y(n_468) );
OR2x6_ASAP7_75t_L g241 ( .A(n_242), .B(n_255), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g242 ( .A1(n_243), .A2(n_244), .B(n_253), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B(n_251), .Y(n_245) );
INVx5_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_248), .B(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_248), .B(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_251), .A2(n_264), .B(n_266), .Y(n_263) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g267 ( .A(n_253), .Y(n_267) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_254), .A2(n_305), .B(n_314), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_254), .B(n_315), .Y(n_314) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_254), .A2(n_329), .B(n_335), .Y(n_328) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx3_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
INVx2_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
AND2x2_ASAP7_75t_L g504 ( .A(n_258), .B(n_346), .Y(n_504) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_267), .B(n_268), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_262), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_261), .A2(n_330), .B(n_331), .Y(n_329) );
INVx4_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
INVx2_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_270), .B(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_270), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_287), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_273), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g424 ( .A(n_273), .B(n_412), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_273), .B(n_401), .Y(n_486) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g346 ( .A(n_274), .Y(n_346) );
AND2x2_ASAP7_75t_L g350 ( .A(n_274), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g391 ( .A(n_274), .B(n_392), .Y(n_391) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_285), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_284), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_282), .Y(n_278) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g301 ( .A(n_283), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_287), .B(n_387), .Y(n_409) );
INVx1_ASAP7_75t_L g448 ( .A(n_287), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_287), .B(n_375), .Y(n_492) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g355 ( .A(n_288), .B(n_350), .Y(n_355) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_290), .B(n_346), .Y(n_379) );
INVx1_ASAP7_75t_L g458 ( .A(n_290), .Y(n_458) );
AOI322xp5_ASAP7_75t_L g482 ( .A1(n_291), .A2(n_397), .A3(n_457), .B1(n_483), .B2(n_485), .C1(n_487), .C2(n_489), .Y(n_482) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_292), .B(n_303), .Y(n_291) );
AND2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_316), .Y(n_337) );
INVx1_ASAP7_75t_SL g340 ( .A(n_292), .Y(n_340) );
AND2x2_ASAP7_75t_L g342 ( .A(n_292), .B(n_304), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_292), .B(n_359), .Y(n_365) );
INVx2_ASAP7_75t_L g384 ( .A(n_292), .Y(n_384) );
AND2x2_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g435 ( .A(n_292), .B(n_359), .Y(n_435) );
BUFx2_ASAP7_75t_L g452 ( .A(n_292), .Y(n_452) );
AND2x2_ASAP7_75t_L g466 ( .A(n_292), .B(n_327), .Y(n_466) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_302), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_303), .B(n_354), .Y(n_381) );
AND2x2_ASAP7_75t_L g508 ( .A(n_303), .B(n_384), .Y(n_508) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_316), .Y(n_303) );
OR2x2_ASAP7_75t_L g353 ( .A(n_304), .B(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
AND2x2_ASAP7_75t_L g404 ( .A(n_304), .B(n_328), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_304), .B(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_304), .Y(n_488) );
INVx2_ASAP7_75t_L g334 ( .A(n_307), .Y(n_334) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g511 ( .A(n_311), .Y(n_511) );
AND2x2_ASAP7_75t_L g339 ( .A(n_316), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
BUFx2_ASAP7_75t_L g367 ( .A(n_316), .Y(n_367) );
AND2x2_ASAP7_75t_L g386 ( .A(n_316), .B(n_359), .Y(n_386) );
INVx3_ASAP7_75t_L g398 ( .A(n_316), .Y(n_398) );
OR2x2_ASAP7_75t_L g408 ( .A(n_316), .B(n_359), .Y(n_408) );
AOI31xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_338), .A3(n_341), .B(n_343), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_337), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_326), .B(n_360), .Y(n_371) );
OR2x2_ASAP7_75t_L g395 ( .A(n_326), .B(n_365), .Y(n_395) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_327), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g416 ( .A(n_327), .B(n_408), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_327), .B(n_398), .Y(n_426) );
AND2x2_ASAP7_75t_L g433 ( .A(n_327), .B(n_434), .Y(n_433) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_327), .B(n_397), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_327), .B(n_452), .Y(n_462) );
AND2x2_ASAP7_75t_L g474 ( .A(n_327), .B(n_359), .Y(n_474) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g354 ( .A(n_328), .Y(n_354) );
INVx1_ASAP7_75t_L g420 ( .A(n_337), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_337), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_339), .B(n_415), .Y(n_449) );
AND2x4_ASAP7_75t_L g360 ( .A(n_340), .B(n_361), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g439 ( .A(n_345), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_345), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g387 ( .A(n_346), .B(n_377), .Y(n_387) );
AND2x2_ASAP7_75t_L g481 ( .A(n_346), .B(n_351), .Y(n_481) );
INVx1_ASAP7_75t_L g506 ( .A(n_346), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_352), .B1(n_355), .B2(n_356), .C(n_362), .Y(n_347) );
CKINVDCx14_ASAP7_75t_R g368 ( .A(n_348), .Y(n_368) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_349), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_352), .B(n_403), .Y(n_422) );
INVx3_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g471 ( .A(n_353), .B(n_367), .Y(n_471) );
AND2x2_ASAP7_75t_L g385 ( .A(n_354), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_354), .B(n_398), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g485 ( .A(n_354), .B(n_455), .C(n_486), .Y(n_485) );
AOI211xp5_ASAP7_75t_SL g418 ( .A1(n_355), .A2(n_419), .B(n_421), .C(n_429), .Y(n_418) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_357), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_358), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_358), .B(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g500 ( .A(n_360), .B(n_474), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_368), .B1(n_369), .B2(n_371), .Y(n_362) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_366), .B(n_415), .Y(n_446) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_369), .A2(n_461), .B1(n_492), .B2(n_499), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_380), .B1(n_382), .B2(n_387), .C(n_388), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_378), .A2(n_389), .B1(n_395), .B2(n_396), .C(n_399), .Y(n_388) );
INVx1_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_SL g403 ( .A(n_384), .Y(n_403) );
OR2x2_ASAP7_75t_L g476 ( .A(n_384), .B(n_408), .Y(n_476) );
AND2x2_ASAP7_75t_L g478 ( .A(n_384), .B(n_386), .Y(n_478) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
AOI21xp33_ASAP7_75t_SL g447 ( .A1(n_390), .A2(n_448), .B(n_449), .Y(n_447) );
OR2x2_ASAP7_75t_L g454 ( .A(n_390), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g428 ( .A(n_391), .B(n_412), .Y(n_428) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp33_ASAP7_75t_SL g445 ( .A(n_396), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_397), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_398), .B(n_434), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_401), .A2(n_414), .B(n_416), .C(n_417), .Y(n_413) );
NAND2x1_ASAP7_75t_SL g438 ( .A(n_401), .B(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_402), .A2(n_451), .B1(n_453), .B2(n_456), .Y(n_450) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_404), .B(n_494), .Y(n_493) );
NAND5xp2_ASAP7_75t_L g405 ( .A(n_406), .B(n_418), .C(n_436), .D(n_450), .E(n_459), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_413), .Y(n_406) );
INVx1_ASAP7_75t_L g463 ( .A(n_409), .Y(n_463) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_411), .A2(n_430), .B1(n_470), .B2(n_472), .C(n_475), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_412), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_415), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_415), .B(n_481), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_427), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g503 ( .A(n_432), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B1(n_444), .B2(n_445), .C(n_447), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g487 ( .A(n_442), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g494 ( .A(n_452), .Y(n_494) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B(n_463), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI211xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B(n_469), .C(n_482), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_467), .A2(n_492), .B(n_493), .C(n_495), .Y(n_491) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_471), .B(n_473), .Y(n_472) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_505), .B(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g527 ( .A(n_510), .Y(n_527) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_513), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
endmodule