module fake_jpeg_2623_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_29),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_66),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_38),
.B1(n_47),
.B2(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_50),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_50),
.C(n_38),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_58),
.B(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_41),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_53),
.B1(n_55),
.B2(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_67),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_107),
.B1(n_108),
.B2(n_5),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_4),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_111),
.C(n_113),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_16),
.B1(n_35),
.B2(n_31),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_14),
.B1(n_28),
.B2(n_27),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_36),
.C(n_24),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_4),
.Y(n_113)
);

XNOR2x1_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_22),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_118),
.B(n_119),
.Y(n_123)
);

NOR4xp25_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_17),
.C(n_12),
.D(n_19),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_122),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_109),
.B1(n_99),
.B2(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.C(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_107),
.B1(n_112),
.B2(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_117),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_124),
.B1(n_115),
.B2(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_123),
.B(n_9),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_8),
.Y(n_134)
);


endmodule