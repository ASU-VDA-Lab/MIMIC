module real_jpeg_22329_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_304, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_304;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_300;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_299;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_0),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_1),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_1),
.A2(n_37),
.B1(n_48),
.B2(n_50),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_2),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_144),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_144),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_2),
.A2(n_27),
.B1(n_36),
.B2(n_144),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_3),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_27),
.B1(n_36),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_4),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_116),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_48),
.B1(n_50),
.B2(n_116),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_116),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_50),
.B(n_60),
.C(n_130),
.D(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_5),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_47),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_83),
.B(n_149),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_33),
.B(n_44),
.C(n_182),
.D(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_5),
.B(n_33),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_118),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_32),
.B(n_34),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_5),
.A2(n_27),
.B1(n_36),
.B2(n_166),
.Y(n_241)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_7),
.B(n_150),
.Y(n_149)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_27),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_11),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_93),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_93),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_93),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_12),
.A2(n_27),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_12),
.A2(n_39),
.B1(n_48),
.B2(n_50),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_12),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_206)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_15),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_95),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_26),
.A2(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_26),
.A2(n_31),
.B1(n_115),
.B2(n_250),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_27),
.A2(n_29),
.B(n_166),
.C(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_31),
.A2(n_35),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_31),
.A2(n_91),
.B(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_45),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_43),
.A2(n_54),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_43),
.A2(n_238),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_44),
.A2(n_47),
.B1(n_74),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_44),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_45),
.B(n_50),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_46),
.A2(n_48),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_54),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_54),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_54),
.A2(n_202),
.B(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_67),
.B1(n_77),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_67),
.B1(n_88),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_59),
.A2(n_67),
.B1(n_143),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_59),
.A2(n_180),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_59),
.A2(n_67),
.B1(n_110),
.B2(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_63),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_60),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_61),
.B(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_64),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_65),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_67),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_67),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_67),
.A2(n_145),
.B(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_90),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_81),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_82),
.A2(n_87),
.B1(n_89),
.B2(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_86),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_83),
.A2(n_85),
.B1(n_192),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_83),
.A2(n_85),
.B1(n_206),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_83),
.A2(n_106),
.B1(n_107),
.B2(n_228),
.Y(n_257)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_155),
.B(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_85),
.B(n_166),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_87),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_94),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_96),
.Y(n_290)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_102),
.A2(n_103),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.C(n_113),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_104),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_105),
.B(n_109),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_107),
.A2(n_164),
.B(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_111),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_112),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_117),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_278),
.A3(n_291),
.B1(n_297),
.B2(n_302),
.C(n_304),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_244),
.C(n_274),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_218),
.B(n_243),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_195),
.B(n_217),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_174),
.B(n_194),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_151),
.B(n_173),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_142),
.C(n_147),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_161),
.B(n_172),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_159),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_167),
.B(n_171),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_187),
.B2(n_193),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_186),
.C(n_193),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_183),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_213),
.C(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_210),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_207),
.C(n_208),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_231),
.C(n_232),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_227),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_256),
.C(n_259),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_272),
.B2(n_273),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_264),
.C(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_269),
.C(n_271),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);


endmodule