module real_jpeg_5197_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_0),
.A2(n_47),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_0),
.A2(n_47),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_0),
.A2(n_47),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_103),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_103),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_2),
.A2(n_103),
.B1(n_165),
.B2(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_3),
.A2(n_258),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_3),
.A2(n_303),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_3),
.A2(n_303),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_3),
.A2(n_303),
.B1(n_411),
.B2(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_4),
.B(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_4),
.A2(n_267),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_4),
.B(n_204),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_4),
.B(n_377),
.C(n_379),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g381 ( 
.A1(n_4),
.A2(n_382),
.B1(n_383),
.B2(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_4),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_4),
.B(n_101),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_4),
.A2(n_153),
.B1(n_322),
.B2(n_428),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_5),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_5),
.A2(n_288),
.B1(n_298),
.B2(n_314),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_5),
.A2(n_298),
.B1(n_385),
.B2(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_5),
.A2(n_298),
.B1(n_417),
.B2(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_7),
.A2(n_78),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_7),
.A2(n_54),
.B1(n_78),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_78),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_8),
.A2(n_139),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_8),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_8),
.A2(n_243),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_8),
.A2(n_243),
.B1(n_405),
.B2(n_408),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_8),
.A2(n_243),
.B1(n_385),
.B2(n_468),
.Y(n_467)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_10),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_10),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_10),
.Y(n_345)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_11),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_14),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_14),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_14),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_14),
.Y(n_269)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_14),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_67),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_15),
.A2(n_67),
.B1(n_132),
.B2(n_139),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_15),
.A2(n_67),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_210),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_208),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_187),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_27),
.B(n_187),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_27),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_27),
.B(n_212),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_108),
.CI(n_151),
.CON(n_27),
.SN(n_27)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_28),
.A2(n_29),
.B(n_71),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_71),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_50),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_30),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_43),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_31),
.A2(n_43),
.B(n_51),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_31),
.A2(n_51),
.B1(n_62),
.B2(n_237),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_31),
.B(n_382),
.Y(n_426)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_32),
.B(n_63),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_32),
.A2(n_52),
.B1(n_174),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_32),
.A2(n_52),
.B1(n_381),
.B2(n_388),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_32),
.A2(n_52),
.B1(n_388),
.B2(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_32),
.A2(n_52),
.B1(n_398),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_36),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_38),
.Y(n_170)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_43),
.A2(n_51),
.B(n_179),
.Y(n_307)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_45),
.Y(n_461)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_46),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_46),
.Y(n_384)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_48),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_49),
.Y(n_387)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_49),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_49),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_62),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_51),
.A2(n_173),
.B(n_179),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_51),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_53)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_54),
.Y(n_375)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_60),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_61),
.Y(n_399)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_70),
.B1(n_85),
.B2(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_70),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_83),
.B1(n_101),
.B2(n_102),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_73),
.A2(n_84),
.B(n_201),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g449 ( 
.A1(n_74),
.A2(n_450),
.A3(n_453),
.B1(n_456),
.B2(n_457),
.Y(n_449)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_75),
.A2(n_382),
.B(n_456),
.Y(n_465)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_76),
.Y(n_293)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_102),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_83),
.B(n_115),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_83),
.A2(n_196),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_83),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_83),
.A2(n_101),
.B1(n_350),
.B2(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_84),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_84),
.A2(n_313),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_84),
.A2(n_313),
.B1(n_316),
.B2(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_86),
.Y(n_459)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_89)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_92),
.Y(n_263)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_92),
.Y(n_315)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_94),
.Y(n_455)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_122),
.B2(n_150),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_120),
.B2(n_121),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_111),
.A2(n_121),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_112),
.B(n_121),
.C(n_122),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_114),
.A2(n_197),
.B(n_316),
.Y(n_334)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_118),
.B(n_382),
.Y(n_456)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_122),
.A2(n_150),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_130),
.B(n_136),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_123),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_123),
.A2(n_141),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_123),
.A2(n_141),
.B1(n_242),
.B2(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_125),
.Y(n_314)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_129),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_181),
.B(n_186),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_140),
.A2(n_204),
.B1(n_295),
.B2(n_301),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_141),
.A2(n_242),
.B(n_245),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_171),
.B(n_180),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_152),
.A2(n_180),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_152),
.A2(n_172),
.B1(n_215),
.B2(n_359),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_161),
.B(n_163),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_153),
.A2(n_271),
.B1(n_279),
.B2(n_283),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_153),
.A2(n_283),
.B(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_153),
.A2(n_230),
.B(n_404),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_153),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_153),
.A2(n_322),
.B1(n_416),
.B2(n_428),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_153),
.A2(n_163),
.B(n_320),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_156),
.Y(n_278)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_156),
.Y(n_411)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_156),
.Y(n_417)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_160),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_160),
.Y(n_437)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_169),
.Y(n_430)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_170),
.Y(n_407)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_170),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_172),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_181),
.B(n_204),
.Y(n_245)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_185),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_202),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_248),
.B(n_499),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_218),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_213),
.B(n_217),
.CI(n_218),
.CON(n_367),
.SN(n_367)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_240),
.C(n_246),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_219),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_234),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_220),
.A2(n_234),
.B1(n_235),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_220),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_230),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_222),
.A2(n_272),
.B(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_361)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_368),
.B(n_493),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_353),
.C(n_365),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_338),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_251),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_326),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_252),
.B(n_326),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_306),
.C(n_318),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_253),
.B(n_352),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_285),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_286),
.C(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_270),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_255),
.B(n_270),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_258),
.A3(n_260),
.B1(n_262),
.B2(n_266),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_284),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.Y(n_285)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_318),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.C(n_312),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_307),
.B(n_308),
.CI(n_312),
.CON(n_340),
.SN(n_340)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_325),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_329),
.C(n_331),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_337),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_336),
.C(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_351),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_339),
.B(n_351),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.C(n_342),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_340),
.B(n_491),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_340),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_341),
.B(n_342),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.C(n_348),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_343),
.A2(n_344),
.B1(n_346),
.B2(n_347),
.Y(n_478)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_348),
.B(n_478),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

A2O1A1O1Ixp25_ASAP7_75t_L g493 ( 
.A1(n_353),
.A2(n_365),
.B(n_494),
.C(n_497),
.D(n_498),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_364),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_354),
.B(n_364),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_358),
.C(n_363),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_360),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_366),
.B(n_367),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_367),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_488),
.B(n_492),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_473),
.B(n_487),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_445),
.B(n_472),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_412),
.B(n_444),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_393),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_373),
.B(n_393),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_380),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_380),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_403),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_402),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_395),
.B(n_402),
.C(n_403),
.Y(n_446)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_397),
.Y(n_402)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_424),
.B(n_443),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_423),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_423),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_431),
.B(n_442),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_426),
.B(n_427),
.Y(n_442)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_438),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_447),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_463),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_464),
.C(n_466),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_462),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_462),
.Y(n_481)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx11_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_475),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_482),
.C(n_485),
.Y(n_489)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_481),
.A2(n_482),
.B1(n_485),
.B2(n_486),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_490),
.Y(n_492)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);


endmodule