module fake_netlist_1_8062_n_1641 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1641);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1641;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1557;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_1607;
wire n_906;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx3_ASAP7_75t_L g374 ( .A(n_109), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_225), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_53), .B(n_19), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_4), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_237), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_372), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_139), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_110), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_338), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_291), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_269), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_214), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_238), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_130), .Y(n_389) );
CKINVDCx16_ASAP7_75t_R g390 ( .A(n_326), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_308), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_50), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_306), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_194), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_149), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_244), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_279), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_286), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_96), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_92), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_213), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_209), .Y(n_404) );
INVxp33_ASAP7_75t_L g405 ( .A(n_79), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_216), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_31), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_165), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_249), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_163), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_6), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_162), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_197), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_228), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_72), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_45), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_203), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_219), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_200), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_180), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_132), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_103), .Y(n_423) );
INVxp33_ASAP7_75t_SL g424 ( .A(n_204), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_359), .B(n_141), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_217), .B(n_163), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_192), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_310), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_92), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_226), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_284), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_116), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_161), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_119), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_320), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_31), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_100), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_256), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_158), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_311), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_154), .B(n_361), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_281), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_307), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_202), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_247), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_230), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_131), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_93), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_39), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_370), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_37), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_51), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_229), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_154), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_111), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_332), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_350), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_343), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_260), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_1), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_241), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_98), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_137), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_294), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_49), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_137), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_171), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_24), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_14), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_14), .Y(n_470) );
BUFx8_ASAP7_75t_SL g471 ( .A(n_150), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_61), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_302), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_47), .B(n_173), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_158), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_336), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_246), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_73), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_147), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_29), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_367), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_280), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_37), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_252), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_352), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_181), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_354), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_56), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_236), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_285), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_297), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_48), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_19), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_59), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_364), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_259), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_132), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_41), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_29), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_314), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_13), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_171), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g503 ( .A(n_282), .B(n_334), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_122), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_165), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_255), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_234), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_342), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_330), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_184), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_239), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_139), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_199), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_106), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_108), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_257), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_347), .Y(n_517) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_180), .B(n_210), .Y(n_518) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_290), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_201), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_198), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_6), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_298), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_48), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_161), .B(n_121), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_181), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_56), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_316), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_258), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_254), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_55), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_251), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_245), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_250), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_10), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_309), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_149), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_301), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_54), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_344), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_3), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_33), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_117), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_221), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_119), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_128), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_104), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_329), .Y(n_548) );
INVxp33_ASAP7_75t_SL g549 ( .A(n_304), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_315), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_188), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_337), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_266), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_106), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_12), .Y(n_555) );
INVxp33_ASAP7_75t_SL g556 ( .A(n_99), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_270), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_2), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_220), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_30), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_287), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_125), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_325), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_235), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_159), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_76), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_351), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_423), .A2(n_3), .B1(n_0), .B2(n_1), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_413), .B(n_0), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_395), .B(n_4), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_374), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_560), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_405), .B(n_5), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_523), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_374), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_374), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_523), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_405), .B(n_5), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_502), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_500), .B(n_7), .Y(n_581) );
OAI22x1_ASAP7_75t_SL g582 ( .A1(n_377), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_502), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_415), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_415), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_416), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_416), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_447), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_463), .B(n_8), .Y(n_591) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_406), .A2(n_187), .B(n_186), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_447), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_406), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_409), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_556), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_463), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_409), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_414), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_414), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_556), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_601) );
INVx6_ASAP7_75t_L g602 ( .A(n_388), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_480), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_512), .Y(n_604) );
AND2x6_ASAP7_75t_L g605 ( .A(n_461), .B(n_189), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_552), .B(n_15), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_461), .Y(n_607) );
INVx6_ASAP7_75t_L g608 ( .A(n_390), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_484), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_480), .B(n_15), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_597), .B(n_442), .Y(n_611) );
BUFx10_ASAP7_75t_L g612 ( .A(n_602), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_595), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_602), .B(n_464), .Y(n_614) );
OR2x6_ASAP7_75t_L g615 ( .A(n_573), .B(n_452), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_575), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_575), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_591), .B(n_384), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_591), .B(n_380), .C(n_375), .Y(n_619) );
INVx6_ASAP7_75t_L g620 ( .A(n_591), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_573), .A2(n_381), .B1(n_392), .B2(n_389), .Y(n_621) );
NAND2xp33_ASAP7_75t_L g622 ( .A(n_605), .B(n_378), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_610), .B(n_384), .Y(n_623) );
INVx5_ASAP7_75t_L g624 ( .A(n_605), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_572), .B(n_436), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_610), .B(n_385), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_592), .Y(n_627) );
NAND2xp33_ASAP7_75t_L g628 ( .A(n_605), .B(n_379), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_579), .A2(n_610), .B1(n_591), .B2(n_581), .Y(n_629) );
INVx4_ASAP7_75t_L g630 ( .A(n_610), .Y(n_630) );
INVx5_ASAP7_75t_L g631 ( .A(n_605), .Y(n_631) );
AND2x6_ASAP7_75t_L g632 ( .A(n_579), .B(n_383), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_602), .B(n_420), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_575), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_595), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_595), .Y(n_637) );
OR2x6_ASAP7_75t_L g638 ( .A(n_579), .B(n_452), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_595), .Y(n_639) );
INVx4_ASAP7_75t_L g640 ( .A(n_605), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_595), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_581), .B(n_519), .Y(n_643) );
BUFx4f_ASAP7_75t_L g644 ( .A(n_605), .Y(n_644) );
INVx8_ASAP7_75t_L g645 ( .A(n_605), .Y(n_645) );
NAND2xp33_ASAP7_75t_L g646 ( .A(n_605), .B(n_417), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_603), .Y(n_647) );
OR2x6_ASAP7_75t_L g648 ( .A(n_568), .B(n_474), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_615), .B(n_570), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_643), .B(n_602), .Y(n_650) );
INVx8_ASAP7_75t_L g651 ( .A(n_615), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_616), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_647), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_647), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_643), .B(n_608), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_633), .B(n_608), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_627), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_615), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_647), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_641), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_630), .B(n_376), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_611), .B(n_608), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_616), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_632), .B(n_608), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_644), .B(n_640), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_615), .B(n_570), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_632), .A2(n_598), .B1(n_599), .B2(n_594), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_634), .Y(n_668) );
NOR2x2_ASAP7_75t_L g669 ( .A(n_615), .B(n_582), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_632), .B(n_606), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_638), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_638), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_632), .B(n_606), .Y(n_673) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_625), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_634), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_638), .Y(n_676) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_630), .B(n_569), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_644), .B(n_387), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_634), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_632), .A2(n_598), .B1(n_599), .B2(n_594), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_634), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_630), .B(n_596), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_616), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g684 ( .A(n_645), .B(n_605), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_627), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_629), .A2(n_431), .B1(n_446), .B2(n_428), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_644), .A2(n_592), .B(n_576), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_632), .B(n_571), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_638), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_617), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_638), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_644), .B(n_393), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_632), .B(n_571), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_630), .B(n_576), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_614), .B(n_538), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_618), .B(n_596), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_623), .B(n_577), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_625), .B(n_469), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_626), .B(n_601), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_620), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_635), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_635), .Y(n_703) );
BUFx8_ASAP7_75t_L g704 ( .A(n_627), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_620), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_648), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_640), .B(n_394), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_621), .A2(n_431), .B1(n_446), .B2(n_428), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_640), .B(n_398), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_612), .B(n_412), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_620), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_619), .B(n_577), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_620), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_613), .Y(n_714) );
OR2x6_ASAP7_75t_L g715 ( .A(n_648), .B(n_568), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_612), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_648), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_619), .A2(n_592), .B(n_583), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_613), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_648), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_612), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_648), .A2(n_612), .B1(n_628), .B2(n_622), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_624), .B(n_510), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_627), .Y(n_724) );
BUFx6f_ASAP7_75t_SL g725 ( .A(n_627), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_645), .B(n_580), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_624), .B(n_399), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_645), .B(n_424), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_642), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_724), .A2(n_646), .B(n_645), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_649), .B(n_382), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_705), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_674), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_651), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_651), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_660), .B(n_471), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_712), .A2(n_526), .B(n_554), .C(n_525), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_695), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_658), .B(n_624), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_649), .B(n_401), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_687), .A2(n_631), .B(n_624), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_708), .B(n_401), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_671), .B(n_624), .Y(n_743) );
INVxp67_ASAP7_75t_L g744 ( .A(n_686), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_711), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_697), .A2(n_476), .B1(n_487), .B2(n_473), .Y(n_746) );
BUFx3_ASAP7_75t_L g747 ( .A(n_682), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_672), .B(n_631), .Y(n_748) );
NOR3xp33_ASAP7_75t_SL g749 ( .A(n_717), .B(n_411), .C(n_407), .Y(n_749) );
NAND2x1p5_ASAP7_75t_L g750 ( .A(n_689), .B(n_631), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_701), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_661), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_715), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_649), .B(n_407), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_666), .B(n_411), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_691), .B(n_631), .Y(n_756) );
O2A1O1Ixp5_ASAP7_75t_L g757 ( .A1(n_718), .A2(n_603), .B(n_567), .C(n_391), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_676), .B(n_545), .C(n_439), .Y(n_758) );
AO32x1_ASAP7_75t_L g759 ( .A1(n_723), .A2(n_413), .A3(n_598), .B1(n_599), .B2(n_594), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_713), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_666), .B(n_486), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_665), .A2(n_637), .B(n_636), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_726), .A2(n_637), .B(n_636), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_715), .A2(n_487), .B1(n_507), .B2(n_476), .Y(n_764) );
O2A1O1Ixp33_ASAP7_75t_SL g765 ( .A1(n_707), .A2(n_400), .B(n_404), .C(n_403), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_666), .B(n_486), .Y(n_766) );
NOR3xp33_ASAP7_75t_SL g767 ( .A(n_669), .B(n_504), .C(n_497), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_710), .B(n_497), .Y(n_768) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_657), .Y(n_769) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_669), .B(n_504), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_713), .Y(n_771) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_657), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_670), .B(n_505), .Y(n_773) );
INVx3_ASAP7_75t_L g774 ( .A(n_701), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_716), .B(n_385), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_682), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_700), .A2(n_396), .B(n_408), .C(n_402), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_650), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_701), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_715), .A2(n_507), .B1(n_607), .B2(n_537), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_667), .A2(n_607), .B1(n_429), .B2(n_555), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_673), .B(n_386), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_696), .B(n_505), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_690), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_697), .B(n_514), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_667), .A2(n_429), .B1(n_555), .B2(n_537), .Y(n_786) );
AOI22x1_ASAP7_75t_L g787 ( .A1(n_677), .A2(n_639), .B1(n_600), .B2(n_609), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_692), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_696), .B(n_514), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_668), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_700), .B(n_424), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_655), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_722), .B(n_680), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_704), .Y(n_794) );
O2A1O1Ixp33_ASAP7_75t_L g795 ( .A1(n_698), .A2(n_421), .B(n_422), .C(n_410), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_706), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_680), .A2(n_549), .B1(n_432), .B2(n_434), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_702), .A2(n_558), .B(n_501), .C(n_437), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_697), .A2(n_549), .B1(n_501), .B2(n_519), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_703), .A2(n_449), .B(n_451), .C(n_433), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_688), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_720), .A2(n_542), .B1(n_543), .B2(n_515), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_709), .A2(n_419), .B(n_418), .Y(n_803) );
O2A1O1Ixp5_ASAP7_75t_SL g804 ( .A1(n_678), .A2(n_585), .B(n_587), .C(n_584), .Y(n_804) );
BUFx12f_ASAP7_75t_L g805 ( .A(n_704), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_694), .A2(n_460), .B(n_462), .C(n_454), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_662), .B(n_515), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_704), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_675), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_656), .B(n_542), .Y(n_810) );
AOI21xp33_ASAP7_75t_L g811 ( .A1(n_728), .A2(n_546), .B(n_543), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_728), .B(n_546), .Y(n_812) );
BUFx3_ASAP7_75t_L g813 ( .A(n_675), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_664), .B(n_547), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_679), .Y(n_815) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_657), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_653), .A2(n_466), .B1(n_467), .B2(n_465), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_721), .B(n_547), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g819 ( .A(n_652), .B(n_386), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_679), .Y(n_820) );
INVx5_ASAP7_75t_L g821 ( .A(n_657), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_653), .A2(n_470), .B1(n_472), .B2(n_468), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_681), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_681), .B(n_566), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_654), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_684), .A2(n_438), .B(n_435), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_678), .A2(n_566), .B1(n_455), .B2(n_478), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_663), .B(n_488), .Y(n_828) );
O2A1O1Ixp33_ASAP7_75t_L g829 ( .A1(n_693), .A2(n_493), .B(n_494), .C(n_492), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_683), .B(n_397), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_693), .A2(n_499), .B(n_522), .C(n_498), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_659), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_659), .A2(n_450), .B(n_440), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_725), .B(n_479), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_685), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_725), .B(n_483), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_L g837 ( .A1(n_727), .A2(n_524), .B(n_535), .C(n_527), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_685), .A2(n_539), .B1(n_562), .B2(n_541), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_729), .A2(n_459), .B(n_456), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_727), .A2(n_565), .B1(n_512), .B2(n_584), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_714), .A2(n_475), .B1(n_531), .B2(n_448), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_719), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_719), .B(n_397), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_674), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_724), .A2(n_490), .B(n_482), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_649), .B(n_489), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_660), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_699), .B(n_585), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_697), .A2(n_495), .B1(n_506), .B2(n_489), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_715), .A2(n_588), .B1(n_590), .B2(n_587), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_674), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_660), .B(n_481), .Y(n_852) );
NOR2xp67_ASAP7_75t_L g853 ( .A(n_660), .B(n_495), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g854 ( .A1(n_687), .A2(n_496), .B(n_491), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_781), .A2(n_441), .B1(n_425), .B2(n_448), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_764), .A2(n_780), .B1(n_781), .B2(n_786), .Y(n_856) );
NAND3xp33_ASAP7_75t_L g857 ( .A(n_758), .B(n_609), .C(n_600), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_746), .B(n_520), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_828), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_786), .B(n_590), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_764), .A2(n_511), .B1(n_513), .B2(n_508), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_741), .A2(n_517), .B(n_516), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_828), .Y(n_863) );
INVx2_ASAP7_75t_SL g864 ( .A(n_805), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_737), .A2(n_604), .B(n_593), .C(n_528), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_848), .Y(n_866) );
OAI21x1_ASAP7_75t_L g867 ( .A1(n_741), .A2(n_551), .B(n_509), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_794), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_730), .A2(n_533), .B(n_530), .Y(n_869) );
BUFx2_ASAP7_75t_SL g870 ( .A(n_808), .Y(n_870) );
INVx4_ASAP7_75t_L g871 ( .A(n_821), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_780), .Y(n_872) );
OAI21xp5_ASAP7_75t_L g873 ( .A1(n_757), .A2(n_536), .B(n_534), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_763), .A2(n_559), .B(n_553), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_744), .A2(n_448), .B1(n_531), .B2(n_475), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_854), .A2(n_563), .B(n_561), .Y(n_876) );
INVx6_ASAP7_75t_L g877 ( .A(n_753), .Y(n_877) );
A2O1A1Ixp33_ASAP7_75t_L g878 ( .A1(n_777), .A2(n_518), .B(n_426), .C(n_564), .Y(n_878) );
AO32x2_ASAP7_75t_L g879 ( .A1(n_850), .A2(n_600), .A3(n_609), .B1(n_595), .B2(n_604), .Y(n_879) );
AO31x2_ASAP7_75t_L g880 ( .A1(n_798), .A2(n_578), .A3(n_586), .B(n_574), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_733), .A2(n_511), .B1(n_513), .B2(n_508), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_784), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_795), .A2(n_503), .B(n_551), .C(n_593), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_788), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_854), .A2(n_544), .B(n_540), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_787), .A2(n_578), .B(n_574), .Y(n_886) );
BUFx2_ASAP7_75t_R g887 ( .A(n_770), .Y(n_887) );
O2A1O1Ixp33_ASAP7_75t_SL g888 ( .A1(n_793), .A2(n_589), .B(n_586), .C(n_191), .Y(n_888) );
BUFx5_ASAP7_75t_L g889 ( .A(n_835), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_752), .Y(n_890) );
A2O1A1Ixp33_ASAP7_75t_L g891 ( .A1(n_829), .A2(n_609), .B(n_600), .C(n_531), .Y(n_891) );
A2O1A1Ixp33_ASAP7_75t_L g892 ( .A1(n_831), .A2(n_600), .B(n_609), .C(n_475), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_L g893 ( .A1(n_800), .A2(n_589), .B(n_18), .C(n_16), .Y(n_893) );
NOR2xp33_ASAP7_75t_SL g894 ( .A(n_844), .B(n_540), .Y(n_894) );
AO31x2_ASAP7_75t_L g895 ( .A1(n_838), .A2(n_609), .A3(n_18), .B(n_16), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_790), .Y(n_896) );
OAI21xp5_ASAP7_75t_L g897 ( .A1(n_804), .A2(n_548), .B(n_544), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_742), .B(n_548), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_762), .A2(n_430), .B(n_427), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_851), .A2(n_444), .B1(n_445), .B2(n_443), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_738), .A2(n_457), .B1(n_458), .B2(n_453), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_785), .B(n_17), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_776), .Y(n_903) );
O2A1O1Ixp33_ASAP7_75t_L g904 ( .A1(n_797), .A2(n_21), .B(n_17), .C(n_20), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_845), .A2(n_485), .B(n_477), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_791), .A2(n_529), .B1(n_532), .B2(n_521), .Y(n_906) );
INVx1_ASAP7_75t_SL g907 ( .A(n_842), .Y(n_907) );
BUFx3_ASAP7_75t_L g908 ( .A(n_747), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_810), .B(n_557), .C(n_550), .Y(n_909) );
CKINVDCx16_ASAP7_75t_R g910 ( .A(n_796), .Y(n_910) );
BUFx12f_ASAP7_75t_L g911 ( .A(n_734), .Y(n_911) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_769), .Y(n_912) );
OAI21xp5_ASAP7_75t_SL g913 ( .A1(n_736), .A2(n_799), .B(n_849), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_778), .B(n_20), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_768), .B(n_21), .Y(n_915) );
INVx2_ASAP7_75t_SL g916 ( .A(n_735), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_792), .B(n_22), .Y(n_917) );
AO31x2_ASAP7_75t_L g918 ( .A1(n_838), .A2(n_26), .A3(n_23), .B(n_25), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_735), .B(n_25), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_809), .Y(n_920) );
O2A1O1Ixp33_ASAP7_75t_L g921 ( .A1(n_797), .A2(n_28), .B(n_26), .C(n_27), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_820), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_837), .A2(n_32), .B(n_27), .C(n_30), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g924 ( .A1(n_812), .A2(n_33), .B(n_34), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_749), .B(n_34), .C(n_35), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_731), .B(n_35), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_815), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_732), .Y(n_928) );
AND2x4_ASAP7_75t_L g929 ( .A(n_853), .B(n_36), .Y(n_929) );
O2A1O1Ixp33_ASAP7_75t_L g930 ( .A1(n_806), .A2(n_39), .B(n_36), .C(n_38), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_802), .B(n_38), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_769), .A2(n_193), .B(n_190), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_740), .B(n_754), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_745), .Y(n_934) );
AOI221x1_ASAP7_75t_L g935 ( .A1(n_826), .A2(n_42), .B1(n_40), .B2(n_41), .C(n_43), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_772), .A2(n_196), .B(n_195), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_823), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_767), .Y(n_938) );
O2A1O1Ixp33_ASAP7_75t_L g939 ( .A1(n_783), .A2(n_43), .B(n_40), .C(n_42), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_789), .B(n_44), .Y(n_940) );
BUFx12f_ASAP7_75t_L g941 ( .A(n_750), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_751), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_755), .B(n_44), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_761), .B(n_45), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_766), .B(n_46), .Y(n_945) );
AO31x2_ASAP7_75t_L g946 ( .A1(n_817), .A2(n_49), .A3(n_46), .B(n_47), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_817), .Y(n_947) );
OAI222xp33_ASAP7_75t_L g948 ( .A1(n_822), .A2(n_50), .B1(n_51), .B2(n_52), .C1(n_53), .C2(n_54), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_801), .A2(n_206), .B(n_205), .Y(n_949) );
AO32x2_ASAP7_75t_L g950 ( .A1(n_822), .A2(n_52), .A3(n_55), .B1(n_57), .B2(n_58), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_811), .B(n_57), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_846), .A2(n_60), .B1(n_58), .B2(n_59), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_833), .A2(n_62), .B(n_60), .C(n_61), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_852), .B(n_62), .Y(n_954) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_816), .Y(n_955) );
CKINVDCx12_ASAP7_75t_R g956 ( .A(n_760), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_825), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_807), .B(n_63), .Y(n_958) );
NOR2x1_ASAP7_75t_R g959 ( .A(n_775), .B(n_63), .Y(n_959) );
AOI21xp5_ASAP7_75t_L g960 ( .A1(n_816), .A2(n_208), .B(n_207), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g961 ( .A(n_818), .B(n_64), .Y(n_961) );
AOI21xp5_ASAP7_75t_L g962 ( .A1(n_843), .A2(n_212), .B(n_211), .Y(n_962) );
INVx3_ASAP7_75t_L g963 ( .A(n_751), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_813), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_771), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_774), .Y(n_966) );
AND2x2_ASAP7_75t_SL g967 ( .A(n_834), .B(n_64), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_814), .A2(n_67), .B1(n_65), .B2(n_66), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_773), .B(n_65), .Y(n_969) );
A2O1A1Ixp33_ASAP7_75t_L g970 ( .A1(n_839), .A2(n_68), .B(n_66), .C(n_67), .Y(n_970) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_821), .Y(n_971) );
NOR2x1_ASAP7_75t_R g972 ( .A(n_821), .B(n_68), .Y(n_972) );
BUFx8_ASAP7_75t_L g973 ( .A(n_832), .Y(n_973) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_827), .A2(n_71), .B1(n_69), .B2(n_70), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_824), .A2(n_71), .B1(n_69), .B2(n_70), .Y(n_975) );
INVx2_ASAP7_75t_SL g976 ( .A(n_819), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_782), .A2(n_76), .B1(n_74), .B2(n_75), .Y(n_977) );
NAND2x1p5_ASAP7_75t_L g978 ( .A(n_821), .B(n_77), .Y(n_978) );
OAI21xp5_ASAP7_75t_SL g979 ( .A1(n_836), .A2(n_77), .B(n_78), .Y(n_979) );
AO31x2_ASAP7_75t_L g980 ( .A1(n_759), .A2(n_80), .A3(n_78), .B(n_79), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_840), .A2(n_80), .B1(n_81), .B2(n_82), .C(n_83), .Y(n_981) );
AO31x2_ASAP7_75t_L g982 ( .A1(n_759), .A2(n_83), .A3(n_81), .B(n_82), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_779), .Y(n_983) );
AOI21xp33_ASAP7_75t_L g984 ( .A1(n_830), .A2(n_84), .B(n_85), .Y(n_984) );
OAI21xp5_ASAP7_75t_L g985 ( .A1(n_803), .A2(n_218), .B(n_215), .Y(n_985) );
BUFx2_ASAP7_75t_L g986 ( .A(n_750), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_841), .B(n_86), .Y(n_987) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_765), .B(n_86), .C(n_87), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_759), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_739), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_743), .A2(n_88), .B1(n_90), .B2(n_91), .Y(n_991) );
AOI21xp5_ASAP7_75t_L g992 ( .A1(n_748), .A2(n_223), .B(n_222), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_756), .A2(n_227), .B(n_224), .Y(n_993) );
A2O1A1Ixp33_ASAP7_75t_L g994 ( .A1(n_777), .A2(n_90), .B(n_91), .C(n_93), .Y(n_994) );
OR2x6_ASAP7_75t_L g995 ( .A(n_805), .B(n_94), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_781), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_744), .B(n_95), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_784), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_744), .B(n_97), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_828), .Y(n_1000) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_741), .A2(n_232), .B(n_231), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_781), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_1002) );
A2O1A1Ixp33_ASAP7_75t_L g1003 ( .A1(n_777), .A2(n_101), .B(n_102), .C(n_103), .Y(n_1003) );
O2A1O1Ixp33_ASAP7_75t_L g1004 ( .A1(n_737), .A2(n_101), .B(n_102), .C(n_104), .Y(n_1004) );
OAI21xp5_ASAP7_75t_L g1005 ( .A1(n_757), .A2(n_240), .B(n_233), .Y(n_1005) );
AND2x2_ASAP7_75t_SL g1006 ( .A(n_808), .B(n_105), .Y(n_1006) );
INVx3_ASAP7_75t_L g1007 ( .A(n_805), .Y(n_1007) );
INVx3_ASAP7_75t_L g1008 ( .A(n_805), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_747), .B(n_105), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_828), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_847), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_856), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_866), .B(n_107), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_1011), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_855), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_1015) );
A2O1A1Ixp33_ASAP7_75t_L g1016 ( .A1(n_940), .A2(n_112), .B(n_113), .C(n_114), .Y(n_1016) );
NOR2xp67_ASAP7_75t_SL g1017 ( .A(n_941), .B(n_114), .Y(n_1017) );
AOI21xp33_ASAP7_75t_L g1018 ( .A1(n_865), .A2(n_115), .B(n_116), .Y(n_1018) );
OAI21xp33_ASAP7_75t_L g1019 ( .A1(n_954), .A2(n_115), .B(n_117), .Y(n_1019) );
OAI21xp5_ASAP7_75t_L g1020 ( .A1(n_933), .A2(n_118), .B(n_120), .Y(n_1020) );
AOI21xp5_ASAP7_75t_L g1021 ( .A1(n_869), .A2(n_243), .B(n_242), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_882), .Y(n_1022) );
BUFx4f_ASAP7_75t_SL g1023 ( .A(n_1007), .Y(n_1023) );
INVx4_ASAP7_75t_SL g1024 ( .A(n_995), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1006), .B(n_120), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_884), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_967), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_1027) );
OAI22xp5_ASAP7_75t_SL g1028 ( .A1(n_995), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1028) );
OR2x6_ASAP7_75t_L g1029 ( .A(n_870), .B(n_124), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_998), .Y(n_1030) );
INVx1_ASAP7_75t_SL g1031 ( .A(n_907), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_986), .B(n_126), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_927), .Y(n_1033) );
AOI21xp33_ASAP7_75t_L g1034 ( .A1(n_913), .A2(n_127), .B(n_128), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_937), .Y(n_1035) );
AOI21xp33_ASAP7_75t_L g1036 ( .A1(n_915), .A2(n_127), .B(n_129), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_957), .Y(n_1037) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_989), .A2(n_253), .B(n_248), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_910), .B(n_129), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_947), .A2(n_131), .B1(n_133), .B2(n_134), .Y(n_1040) );
NAND2x1p5_ASAP7_75t_L g1041 ( .A(n_1007), .B(n_133), .Y(n_1041) );
AOI21xp5_ASAP7_75t_L g1042 ( .A1(n_969), .A2(n_292), .B(n_369), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g1043 ( .A1(n_876), .A2(n_289), .B(n_368), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_883), .A2(n_134), .B(n_135), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g1045 ( .A1(n_898), .A2(n_135), .B1(n_136), .B2(n_138), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_927), .Y(n_1046) );
A2O1A1Ixp33_ASAP7_75t_L g1047 ( .A1(n_958), .A2(n_136), .B(n_138), .C(n_140), .Y(n_1047) );
AO21x2_ASAP7_75t_L g1048 ( .A1(n_897), .A2(n_295), .B(n_366), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_860), .A2(n_140), .B1(n_141), .B2(n_142), .Y(n_1049) );
A2O1A1Ixp33_ASAP7_75t_L g1050 ( .A1(n_961), .A2(n_142), .B(n_143), .C(n_144), .Y(n_1050) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_894), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_1051) );
A2O1A1Ixp33_ASAP7_75t_L g1052 ( .A1(n_1004), .A2(n_145), .B(n_146), .C(n_147), .Y(n_1052) );
INVx6_ASAP7_75t_L g1053 ( .A(n_973), .Y(n_1053) );
AOI21xp5_ASAP7_75t_L g1054 ( .A1(n_874), .A2(n_299), .B(n_365), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_896), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_951), .A2(n_858), .B1(n_931), .B2(n_902), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_868), .B(n_146), .Y(n_1057) );
OAI22x1_ASAP7_75t_L g1058 ( .A1(n_1009), .A2(n_148), .B1(n_150), .B2(n_151), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_859), .B(n_148), .Y(n_1059) );
OAI21xp5_ASAP7_75t_L g1060 ( .A1(n_997), .A2(n_152), .B(n_153), .Y(n_1060) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_973), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_887), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_911), .Y(n_1063) );
CKINVDCx12_ASAP7_75t_R g1064 ( .A(n_972), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_861), .A2(n_153), .B1(n_155), .B2(n_156), .Y(n_1065) );
OA21x2_ASAP7_75t_L g1066 ( .A1(n_886), .A2(n_300), .B(n_362), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_920), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_871), .B(n_155), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1069 ( .A1(n_873), .A2(n_943), .B(n_926), .Y(n_1069) );
NAND2x1p5_ASAP7_75t_L g1070 ( .A(n_1008), .B(n_156), .Y(n_1070) );
BUFx5_ASAP7_75t_L g1071 ( .A(n_928), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_863), .B(n_157), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_862), .A2(n_303), .B(n_360), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_890), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_919), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_871), .B(n_157), .Y(n_1076) );
A2O1A1Ixp33_ASAP7_75t_L g1077 ( .A1(n_893), .A2(n_159), .B(n_160), .C(n_162), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_919), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1000), .B(n_160), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_1008), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_934), .Y(n_1081) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_996), .A2(n_164), .B1(n_166), .B2(n_167), .C(n_168), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_979), .A2(n_164), .B1(n_166), .B2(n_167), .C(n_168), .Y(n_1083) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_1009), .A2(n_169), .B1(n_170), .B2(n_172), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_903), .B(n_169), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_945), .A2(n_170), .B1(n_172), .B2(n_173), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_1010), .A2(n_174), .B1(n_175), .B2(n_176), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_908), .B(n_174), .Y(n_1088) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_938), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_971), .B(n_175), .Y(n_1090) );
OA21x2_ASAP7_75t_L g1091 ( .A1(n_949), .A2(n_313), .B(n_358), .Y(n_1091) );
AO21x2_ASAP7_75t_L g1092 ( .A1(n_891), .A2(n_312), .B(n_356), .Y(n_1092) );
AO31x2_ASAP7_75t_L g1093 ( .A1(n_935), .A2(n_176), .A3(n_177), .B(n_178), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_971), .B(n_916), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_978), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_944), .B(n_177), .Y(n_1096) );
AOI21xp5_ASAP7_75t_L g1097 ( .A1(n_962), .A2(n_317), .B(n_355), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_922), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_971), .B(n_178), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_999), .A2(n_318), .B(n_349), .Y(n_1100) );
A2O1A1Ixp33_ASAP7_75t_L g1101 ( .A1(n_904), .A2(n_179), .B(n_182), .C(n_183), .Y(n_1101) );
OA21x2_ASAP7_75t_L g1102 ( .A1(n_985), .A2(n_305), .B(n_348), .Y(n_1102) );
OAI22xp5_ASAP7_75t_SL g1103 ( .A1(n_956), .A2(n_179), .B1(n_182), .B2(n_183), .Y(n_1103) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_881), .A2(n_185), .B1(n_261), .B2(n_262), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_968), .A2(n_185), .B1(n_263), .B2(n_264), .Y(n_1105) );
NAND3x1_ASAP7_75t_L g1106 ( .A(n_988), .B(n_265), .C(n_267), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_1001), .A2(n_268), .B(n_271), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_914), .B(n_272), .Y(n_1108) );
OAI21xp5_ASAP7_75t_L g1109 ( .A1(n_878), .A2(n_273), .B(n_274), .Y(n_1109) );
OAI21x1_ASAP7_75t_L g1110 ( .A1(n_932), .A2(n_275), .B(n_276), .Y(n_1110) );
OAI21xp5_ASAP7_75t_L g1111 ( .A1(n_885), .A2(n_917), .B(n_857), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_976), .B(n_371), .Y(n_1112) );
OAI21x1_ASAP7_75t_L g1113 ( .A1(n_936), .A2(n_277), .B(n_278), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_1002), .A2(n_283), .B1(n_288), .B2(n_293), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_877), .A2(n_296), .B1(n_319), .B2(n_321), .Y(n_1115) );
OR2x6_ASAP7_75t_L g1116 ( .A(n_864), .B(n_322), .Y(n_1116) );
BUFx4f_ASAP7_75t_SL g1117 ( .A(n_929), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1118 ( .A(n_877), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_906), .B(n_964), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_965), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_899), .A2(n_323), .B(n_324), .Y(n_1121) );
AOI21xp33_ASAP7_75t_L g1122 ( .A1(n_959), .A2(n_327), .B(n_328), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_946), .Y(n_1123) );
AO21x2_ASAP7_75t_L g1124 ( .A1(n_892), .A2(n_331), .B(n_333), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_946), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_946), .Y(n_1126) );
A2O1A1Ixp33_ASAP7_75t_L g1127 ( .A1(n_921), .A2(n_339), .B(n_340), .C(n_341), .Y(n_1127) );
AOI322xp5_ASAP7_75t_L g1128 ( .A1(n_974), .A2(n_345), .A3(n_346), .B1(n_929), .B2(n_981), .C1(n_924), .C2(n_991), .Y(n_1128) );
BUFx6f_ASAP7_75t_L g1129 ( .A(n_912), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_925), .A2(n_984), .B1(n_952), .B2(n_987), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1131 ( .A1(n_994), .A2(n_1003), .B1(n_923), .B2(n_977), .C(n_930), .Y(n_1131) );
OA21x2_ASAP7_75t_L g1132 ( .A1(n_875), .A2(n_960), .B(n_953), .Y(n_1132) );
OR2x6_ASAP7_75t_L g1133 ( .A(n_939), .B(n_975), .Y(n_1133) );
INVx4_ASAP7_75t_SL g1134 ( .A(n_918), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g1135 ( .A(n_955), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_901), .B(n_983), .Y(n_1136) );
NAND2xp5_ASAP7_75t_SL g1137 ( .A(n_889), .B(n_900), .Y(n_1137) );
OAI21xp5_ASAP7_75t_L g1138 ( .A1(n_905), .A2(n_909), .B(n_970), .Y(n_1138) );
INVx3_ASAP7_75t_L g1139 ( .A(n_942), .Y(n_1139) );
NAND2x1_ASAP7_75t_L g1140 ( .A(n_942), .B(n_963), .Y(n_1140) );
AOI21xp33_ASAP7_75t_L g1141 ( .A1(n_966), .A2(n_963), .B(n_990), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_918), .B(n_895), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_918), .B(n_895), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_880), .Y(n_1144) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_889), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_992), .B(n_993), .Y(n_1146) );
AOI222xp33_ASAP7_75t_L g1147 ( .A1(n_948), .A2(n_950), .B1(n_895), .B2(n_980), .C1(n_982), .C2(n_879), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_950), .Y(n_1148) );
OAI21xp33_ASAP7_75t_SL g1149 ( .A1(n_950), .A2(n_879), .B(n_980), .Y(n_1149) );
OAI21x1_ASAP7_75t_L g1150 ( .A1(n_879), .A2(n_889), .B(n_980), .Y(n_1150) );
AOI21xp5_ASAP7_75t_L g1151 ( .A1(n_889), .A2(n_854), .B(n_888), .Y(n_1151) );
A2O1A1Ixp33_ASAP7_75t_L g1152 ( .A1(n_982), .A2(n_940), .B(n_958), .C(n_961), .Y(n_1152) );
INVx2_ASAP7_75t_L g1153 ( .A(n_982), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_889), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_910), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_856), .B(n_715), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_856), .A2(n_674), .B1(n_764), .B2(n_686), .Y(n_1157) );
AO21x2_ASAP7_75t_L g1158 ( .A1(n_989), .A2(n_1005), .B(n_854), .Y(n_1158) );
OA21x2_ASAP7_75t_L g1159 ( .A1(n_989), .A2(n_867), .B(n_1005), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_856), .A2(n_781), .B1(n_780), .B2(n_764), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_856), .B(n_715), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1162 ( .A1(n_933), .A2(n_757), .B(n_876), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_884), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_884), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_927), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1074), .Y(n_1166) );
INVxp67_ASAP7_75t_R g1167 ( .A(n_1028), .Y(n_1167) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_1053), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1157), .B(n_1160), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1156), .B(n_1161), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1046), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1026), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1163), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1164), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1165), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1035), .B(n_1037), .Y(n_1176) );
BUFx6f_ASAP7_75t_L g1177 ( .A(n_1129), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1022), .B(n_1033), .Y(n_1178) );
OR2x6_ASAP7_75t_L g1179 ( .A(n_1116), .B(n_1029), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1055), .B(n_1067), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1098), .B(n_1030), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1117), .A2(n_1116), .B1(n_1027), .B2(n_1083), .Y(n_1182) );
OR2x2_ASAP7_75t_SL g1183 ( .A(n_1053), .B(n_1142), .Y(n_1183) );
INVxp67_ASAP7_75t_L g1184 ( .A(n_1014), .Y(n_1184) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_1032), .Y(n_1185) );
AO21x2_ASAP7_75t_L g1186 ( .A1(n_1152), .A2(n_1125), .B(n_1123), .Y(n_1186) );
A2O1A1Ixp33_ASAP7_75t_L g1187 ( .A1(n_1128), .A2(n_1020), .B(n_1034), .C(n_1101), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1032), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1081), .Y(n_1189) );
AO21x2_ASAP7_75t_L g1190 ( .A1(n_1126), .A2(n_1151), .B(n_1153), .Y(n_1190) );
AO21x2_ASAP7_75t_L g1191 ( .A1(n_1126), .A2(n_1144), .B(n_1158), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1013), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1120), .Y(n_1193) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_1069), .A2(n_1131), .B(n_1162), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1068), .B(n_1076), .Y(n_1195) );
INVx3_ASAP7_75t_L g1196 ( .A(n_1071), .Y(n_1196) );
INVx3_ASAP7_75t_L g1197 ( .A(n_1071), .Y(n_1197) );
BUFx6f_ASAP7_75t_L g1198 ( .A(n_1129), .Y(n_1198) );
OAI21xp5_ASAP7_75t_L g1199 ( .A1(n_1052), .A2(n_1130), .B(n_1138), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1075), .B(n_1078), .Y(n_1200) );
AO21x2_ASAP7_75t_L g1201 ( .A1(n_1144), .A2(n_1158), .B(n_1148), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1029), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1076), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1071), .Y(n_1204) );
INVx1_ASAP7_75t_SL g1205 ( .A(n_1063), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1085), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1059), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1072), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1079), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1090), .B(n_1099), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1129), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1095), .B(n_1136), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1058), .Y(n_1213) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_1154), .B(n_1094), .Y(n_1214) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1135), .Y(n_1215) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1135), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1154), .B(n_1094), .Y(n_1217) );
BUFx2_ASAP7_75t_L g1218 ( .A(n_1024), .Y(n_1218) );
INVx4_ASAP7_75t_L g1219 ( .A(n_1024), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1090), .B(n_1099), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1159), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_1084), .A2(n_1065), .B1(n_1045), .B2(n_1086), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1060), .B(n_1134), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1134), .B(n_1025), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1041), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1070), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1227 ( .A1(n_1064), .A2(n_1057), .B1(n_1061), .B2(n_1012), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1044), .B(n_1093), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1031), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_1145), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1093), .B(n_1139), .Y(n_1231) );
OAI21xp5_ASAP7_75t_L g1232 ( .A1(n_1077), .A2(n_1018), .B(n_1111), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1096), .B(n_1119), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1049), .Y(n_1234) );
AOI33xp33_ASAP7_75t_L g1235 ( .A1(n_1088), .A2(n_1040), .A3(n_1087), .B1(n_1051), .B2(n_1082), .B3(n_1105), .Y(n_1235) );
INVx3_ASAP7_75t_L g1236 ( .A(n_1140), .Y(n_1236) );
OAI21xp5_ASAP7_75t_L g1237 ( .A1(n_1127), .A2(n_1109), .B(n_1050), .Y(n_1237) );
OAI21xp5_ASAP7_75t_L g1238 ( .A1(n_1047), .A2(n_1016), .B(n_1019), .Y(n_1238) );
INVx3_ASAP7_75t_L g1239 ( .A(n_1139), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1088), .Y(n_1240) );
HB1xp67_ASAP7_75t_L g1241 ( .A(n_1080), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1015), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1066), .Y(n_1243) );
INVxp67_ASAP7_75t_L g1244 ( .A(n_1017), .Y(n_1244) );
OR2x6_ASAP7_75t_L g1245 ( .A(n_1133), .B(n_1137), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1118), .B(n_1036), .Y(n_1246) );
BUFx2_ASAP7_75t_L g1247 ( .A(n_1155), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1093), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1103), .Y(n_1249) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1066), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1147), .B(n_1133), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1039), .B(n_1023), .Y(n_1252) );
INVx3_ASAP7_75t_SL g1253 ( .A(n_1062), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1112), .Y(n_1254) );
AND2x4_ASAP7_75t_L g1255 ( .A(n_1146), .B(n_1092), .Y(n_1255) );
OAI221xp5_ASAP7_75t_SL g1256 ( .A1(n_1149), .A2(n_1104), .B1(n_1115), .B2(n_1043), .C(n_1108), .Y(n_1256) );
BUFx3_ASAP7_75t_L g1257 ( .A(n_1089), .Y(n_1257) );
INVx1_ASAP7_75t_SL g1258 ( .A(n_1122), .Y(n_1258) );
BUFx3_ASAP7_75t_L g1259 ( .A(n_1110), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1106), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1113), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1132), .B(n_1048), .Y(n_1262) );
AO21x2_ASAP7_75t_L g1263 ( .A1(n_1048), .A2(n_1038), .B(n_1141), .Y(n_1263) );
OAI211xp5_ASAP7_75t_L g1264 ( .A1(n_1100), .A2(n_1042), .B(n_1021), .C(n_1054), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1132), .B(n_1124), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1114), .B(n_1121), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1124), .B(n_1073), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1107), .A2(n_913), .B1(n_1056), .B2(n_1157), .C(n_979), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1097), .B(n_1156), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1157), .B(n_872), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1046), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1160), .B(n_1156), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1074), .Y(n_1273) );
OA21x2_ASAP7_75t_L g1274 ( .A1(n_1143), .A2(n_1150), .B(n_1125), .Y(n_1274) );
OR2x6_ASAP7_75t_L g1275 ( .A(n_1116), .B(n_978), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1156), .B(n_1161), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1157), .B(n_872), .Y(n_1277) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_1053), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1160), .B(n_1156), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1160), .A2(n_1156), .B1(n_1161), .B2(n_715), .Y(n_1280) );
OA21x2_ASAP7_75t_L g1281 ( .A1(n_1143), .A2(n_1150), .B(n_1125), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1074), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_1160), .A2(n_1156), .B1(n_1161), .B2(n_715), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1074), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1156), .B(n_1161), .Y(n_1285) );
INVx2_ASAP7_75t_SL g1286 ( .A(n_1053), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1156), .B(n_1161), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1156), .B(n_1161), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1074), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_1117), .Y(n_1290) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1046), .B(n_1165), .Y(n_1291) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_1014), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_1014), .Y(n_1293) );
AOI21xp5_ASAP7_75t_SL g1294 ( .A1(n_1091), .A2(n_1102), .B(n_972), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1074), .Y(n_1295) );
OA21x2_ASAP7_75t_L g1296 ( .A1(n_1143), .A2(n_1150), .B(n_1125), .Y(n_1296) );
OR2x6_ASAP7_75t_L g1297 ( .A(n_1116), .B(n_978), .Y(n_1297) );
OA21x2_ASAP7_75t_L g1298 ( .A1(n_1143), .A2(n_1150), .B(n_1125), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1276), .B(n_1285), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1171), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1276), .B(n_1285), .Y(n_1301) );
BUFx3_ASAP7_75t_L g1302 ( .A(n_1290), .Y(n_1302) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1171), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1287), .B(n_1288), .Y(n_1304) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1175), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_1169), .A2(n_1179), .B1(n_1280), .B2(n_1283), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1287), .B(n_1288), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1271), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_1169), .A2(n_1268), .B1(n_1249), .B2(n_1179), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1291), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1311 ( .A(n_1293), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1272), .B(n_1279), .Y(n_1312) );
BUFx3_ASAP7_75t_L g1313 ( .A(n_1168), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1272), .B(n_1279), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1251), .B(n_1178), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1251), .B(n_1178), .Y(n_1316) );
INVxp67_ASAP7_75t_SL g1317 ( .A(n_1230), .Y(n_1317) );
NAND2x1p5_ASAP7_75t_SL g1318 ( .A(n_1223), .B(n_1265), .Y(n_1318) );
AND2x4_ASAP7_75t_L g1319 ( .A(n_1255), .B(n_1231), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1176), .B(n_1181), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1176), .B(n_1181), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1170), .B(n_1180), .Y(n_1322) );
INVxp67_ASAP7_75t_L g1323 ( .A(n_1292), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1180), .B(n_1231), .Y(n_1324) );
INVx1_ASAP7_75t_SL g1325 ( .A(n_1205), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1326 ( .A(n_1244), .B(n_1179), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1269), .B(n_1186), .Y(n_1327) );
OAI21xp5_ASAP7_75t_L g1328 ( .A1(n_1187), .A2(n_1222), .B(n_1199), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1186), .B(n_1228), .Y(n_1329) );
NAND2x1_ASAP7_75t_L g1330 ( .A(n_1196), .B(n_1197), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1183), .B(n_1212), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1332 ( .A(n_1255), .B(n_1196), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1228), .B(n_1166), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1183), .B(n_1212), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_1179), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1172), .B(n_1173), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1248), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1174), .B(n_1273), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1201), .Y(n_1339) );
BUFx2_ASAP7_75t_L g1340 ( .A(n_1197), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1282), .B(n_1284), .Y(n_1341) );
AND2x2_ASAP7_75t_SL g1342 ( .A(n_1195), .B(n_1223), .Y(n_1342) );
NAND2x1p5_ASAP7_75t_SL g1343 ( .A(n_1195), .B(n_1265), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1289), .B(n_1295), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_1182), .A2(n_1234), .B1(n_1213), .B2(n_1297), .Y(n_1345) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1221), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1189), .B(n_1224), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1270), .B(n_1277), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1206), .B(n_1233), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1224), .B(n_1201), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1233), .B(n_1192), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1201), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1191), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1191), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1191), .Y(n_1355) );
INVx5_ASAP7_75t_L g1356 ( .A(n_1275), .Y(n_1356) );
INVx1_ASAP7_75t_SL g1357 ( .A(n_1241), .Y(n_1357) );
BUFx2_ASAP7_75t_L g1358 ( .A(n_1275), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1194), .B(n_1193), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1184), .B(n_1185), .Y(n_1360) );
INVx3_ASAP7_75t_L g1361 ( .A(n_1177), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1204), .B(n_1274), .Y(n_1362) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1246), .B(n_1227), .C(n_1260), .Y(n_1363) );
BUFx3_ASAP7_75t_L g1364 ( .A(n_1168), .Y(n_1364) );
INVxp67_ASAP7_75t_SL g1365 ( .A(n_1210), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1274), .B(n_1281), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1281), .B(n_1296), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1281), .B(n_1296), .Y(n_1368) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_1214), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1188), .B(n_1229), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1371 ( .A(n_1275), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1296), .B(n_1298), .Y(n_1372) );
BUFx2_ASAP7_75t_L g1373 ( .A(n_1275), .Y(n_1373) );
INVx3_ASAP7_75t_L g1374 ( .A(n_1177), .Y(n_1374) );
BUFx2_ASAP7_75t_L g1375 ( .A(n_1297), .Y(n_1375) );
BUFx3_ASAP7_75t_L g1376 ( .A(n_1278), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1214), .B(n_1217), .Y(n_1377) );
BUFx2_ASAP7_75t_L g1378 ( .A(n_1297), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1214), .B(n_1217), .Y(n_1379) );
AND2x4_ASAP7_75t_L g1380 ( .A(n_1245), .B(n_1190), .Y(n_1380) );
BUFx2_ASAP7_75t_L g1381 ( .A(n_1297), .Y(n_1381) );
BUFx2_ASAP7_75t_L g1382 ( .A(n_1198), .Y(n_1382) );
NOR2x1_ASAP7_75t_L g1383 ( .A(n_1294), .B(n_1236), .Y(n_1383) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_1319), .B(n_1245), .Y(n_1384) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1346), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1324), .B(n_1262), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1324), .B(n_1262), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1320), .B(n_1240), .Y(n_1388) );
AOI21xp33_ASAP7_75t_SL g1389 ( .A1(n_1343), .A2(n_1253), .B(n_1286), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1336), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1336), .Y(n_1391) );
NAND2x1p5_ASAP7_75t_L g1392 ( .A(n_1356), .B(n_1219), .Y(n_1392) );
NAND2xp5_ASAP7_75t_SL g1393 ( .A(n_1356), .B(n_1219), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1333), .B(n_1245), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1329), .B(n_1245), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1329), .B(n_1210), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g1397 ( .A(n_1323), .Y(n_1397) );
INVx3_ASAP7_75t_L g1398 ( .A(n_1330), .Y(n_1398) );
BUFx2_ASAP7_75t_L g1399 ( .A(n_1317), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1341), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1327), .B(n_1220), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1320), .B(n_1200), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1321), .B(n_1202), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1337), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1327), .B(n_1220), .Y(n_1405) );
INVx6_ASAP7_75t_L g1406 ( .A(n_1356), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1348), .B(n_1203), .Y(n_1407) );
AND2x4_ASAP7_75t_L g1408 ( .A(n_1319), .B(n_1236), .Y(n_1408) );
NAND2x1p5_ASAP7_75t_L g1409 ( .A(n_1356), .B(n_1219), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1321), .B(n_1242), .Y(n_1410) );
AND2x4_ASAP7_75t_L g1411 ( .A(n_1319), .B(n_1236), .Y(n_1411) );
INVx1_ASAP7_75t_SL g1412 ( .A(n_1357), .Y(n_1412) );
INVxp67_ASAP7_75t_L g1413 ( .A(n_1311), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1337), .Y(n_1414) );
AOI22xp33_ASAP7_75t_SL g1415 ( .A1(n_1356), .A2(n_1218), .B1(n_1225), .B2(n_1226), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1312), .B(n_1209), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1312), .B(n_1208), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1314), .B(n_1207), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1300), .Y(n_1419) );
NAND2xp5_ASAP7_75t_SL g1420 ( .A(n_1356), .B(n_1286), .Y(n_1420) );
HB1xp67_ASAP7_75t_L g1421 ( .A(n_1370), .Y(n_1421) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_1319), .B(n_1259), .Y(n_1422) );
AND2x2_ASAP7_75t_SL g1423 ( .A(n_1342), .B(n_1235), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1314), .B(n_1232), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1350), .B(n_1211), .Y(n_1425) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1315), .B(n_1211), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1341), .Y(n_1427) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_1325), .B(n_1252), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_1328), .A2(n_1238), .B1(n_1266), .B2(n_1237), .Y(n_1429) );
AND2x4_ASAP7_75t_L g1430 ( .A(n_1332), .B(n_1259), .Y(n_1430) );
NAND2x1p5_ASAP7_75t_L g1431 ( .A(n_1358), .B(n_1198), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1300), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1322), .B(n_1239), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1308), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1350), .B(n_1216), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_1315), .B(n_1216), .Y(n_1436) );
AND2x4_ASAP7_75t_SL g1437 ( .A(n_1371), .B(n_1239), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1322), .B(n_1254), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1316), .B(n_1215), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1316), .B(n_1215), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1343), .B(n_1267), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1344), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1344), .Y(n_1443) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1302), .B(n_1247), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1299), .B(n_1243), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1299), .B(n_1235), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1301), .B(n_1250), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1301), .B(n_1250), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1338), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1304), .B(n_1261), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1304), .B(n_1263), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1307), .B(n_1263), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1307), .B(n_1278), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1310), .B(n_1263), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1308), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1390), .B(n_1391), .Y(n_1456) );
INVx1_ASAP7_75t_SL g1457 ( .A(n_1412), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1399), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1386), .B(n_1362), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1400), .B(n_1359), .Y(n_1460) );
INVxp67_ASAP7_75t_L g1461 ( .A(n_1397), .Y(n_1461) );
A2O1A1Ixp33_ASAP7_75t_L g1462 ( .A1(n_1423), .A2(n_1331), .B(n_1334), .C(n_1381), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1386), .B(n_1362), .Y(n_1463) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1404), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1427), .Y(n_1465) );
AOI22xp5_ASAP7_75t_L g1466 ( .A1(n_1423), .A2(n_1345), .B1(n_1306), .B2(n_1167), .Y(n_1466) );
NAND2x1p5_ASAP7_75t_L g1467 ( .A(n_1393), .B(n_1358), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1387), .B(n_1366), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1387), .B(n_1366), .Y(n_1469) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1416), .B(n_1331), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1442), .Y(n_1471) );
INVx2_ASAP7_75t_SL g1472 ( .A(n_1406), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1451), .B(n_1367), .Y(n_1473) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1424), .B(n_1318), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1424), .B(n_1318), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1451), .B(n_1367), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1443), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1452), .B(n_1368), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1404), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1452), .B(n_1368), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1450), .B(n_1372), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1450), .B(n_1372), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1401), .B(n_1380), .Y(n_1483) );
INVx2_ASAP7_75t_L g1484 ( .A(n_1414), .Y(n_1484) );
INVx2_ASAP7_75t_L g1485 ( .A(n_1414), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1419), .Y(n_1486) );
BUFx2_ASAP7_75t_L g1487 ( .A(n_1392), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1417), .B(n_1318), .Y(n_1488) );
INVx2_ASAP7_75t_L g1489 ( .A(n_1385), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1419), .Y(n_1490) );
AND2x4_ASAP7_75t_L g1491 ( .A(n_1408), .B(n_1380), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1492 ( .A(n_1417), .B(n_1347), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1401), .B(n_1380), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1405), .B(n_1380), .Y(n_1494) );
AOI22xp5_ASAP7_75t_L g1495 ( .A1(n_1429), .A2(n_1306), .B1(n_1309), .B2(n_1363), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1410), .B(n_1349), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1432), .Y(n_1497) );
AND2x4_ASAP7_75t_L g1498 ( .A(n_1408), .B(n_1332), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1405), .B(n_1353), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1449), .B(n_1351), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1432), .Y(n_1501) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_1418), .B(n_1303), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1434), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1434), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1421), .B(n_1335), .Y(n_1505) );
AND2x2_ASAP7_75t_SL g1506 ( .A(n_1384), .B(n_1342), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1418), .B(n_1303), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_1402), .B(n_1305), .Y(n_1508) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1455), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1446), .B(n_1396), .Y(n_1510) );
OAI21xp33_ASAP7_75t_L g1511 ( .A1(n_1441), .A2(n_1360), .B(n_1326), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1445), .B(n_1447), .Y(n_1512) );
NOR2x1_ASAP7_75t_L g1513 ( .A(n_1444), .B(n_1302), .Y(n_1513) );
INVx1_ASAP7_75t_SL g1514 ( .A(n_1457), .Y(n_1514) );
OAI32xp33_ASAP7_75t_L g1515 ( .A1(n_1488), .A2(n_1409), .A3(n_1392), .B1(n_1441), .B2(n_1413), .Y(n_1515) );
NAND2xp5_ASAP7_75t_SL g1516 ( .A(n_1506), .B(n_1389), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1473), .B(n_1476), .Y(n_1517) );
A2O1A1Ixp33_ASAP7_75t_L g1518 ( .A1(n_1506), .A2(n_1373), .B(n_1375), .C(n_1378), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1456), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1466), .A2(n_1342), .B1(n_1381), .B2(n_1378), .Y(n_1520) );
INVxp67_ASAP7_75t_L g1521 ( .A(n_1513), .Y(n_1521) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1489), .Y(n_1522) );
AOI22xp5_ASAP7_75t_L g1523 ( .A1(n_1495), .A2(n_1375), .B1(n_1373), .B2(n_1395), .Y(n_1523) );
OR2x2_ASAP7_75t_L g1524 ( .A(n_1492), .B(n_1445), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1473), .B(n_1447), .Y(n_1525) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_1511), .B(n_1403), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_1512), .B(n_1448), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1470), .Y(n_1528) );
INVx2_ASAP7_75t_L g1529 ( .A(n_1464), .Y(n_1529) );
INVx1_ASAP7_75t_SL g1530 ( .A(n_1512), .Y(n_1530) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1464), .Y(n_1531) );
AND2x4_ASAP7_75t_SL g1532 ( .A(n_1498), .B(n_1408), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1533 ( .A(n_1461), .Y(n_1533) );
NOR2x1_ASAP7_75t_L g1534 ( .A(n_1487), .B(n_1420), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1479), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1476), .B(n_1448), .Y(n_1536) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1465), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1478), .B(n_1425), .Y(n_1538) );
NAND2xp5_ASAP7_75t_SL g1539 ( .A(n_1462), .B(n_1398), .Y(n_1539) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1484), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1510), .B(n_1439), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1471), .Y(n_1542) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1477), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1486), .Y(n_1544) );
NOR2xp33_ASAP7_75t_L g1545 ( .A(n_1505), .B(n_1453), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1546 ( .A(n_1499), .B(n_1439), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1547 ( .A(n_1468), .B(n_1426), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1499), .B(n_1440), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1478), .B(n_1425), .Y(n_1549) );
NAND2x1_ASAP7_75t_SL g1550 ( .A(n_1491), .B(n_1253), .Y(n_1550) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1468), .B(n_1426), .Y(n_1551) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1529), .Y(n_1552) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1529), .Y(n_1553) );
INVx1_ASAP7_75t_SL g1554 ( .A(n_1514), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1526), .B(n_1480), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1517), .B(n_1480), .Y(n_1556) );
HB1xp67_ASAP7_75t_L g1557 ( .A(n_1530), .Y(n_1557) );
O2A1O1Ixp33_ASAP7_75t_L g1558 ( .A1(n_1539), .A2(n_1462), .B(n_1428), .C(n_1500), .Y(n_1558) );
AOI222xp33_ASAP7_75t_SL g1559 ( .A1(n_1520), .A2(n_1458), .B1(n_1501), .B2(n_1509), .C1(n_1504), .C2(n_1503), .Y(n_1559) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1535), .Y(n_1560) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1544), .Y(n_1561) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1537), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1542), .Y(n_1563) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1533), .B(n_1496), .Y(n_1564) );
HB1xp67_ASAP7_75t_L g1565 ( .A(n_1521), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1531), .Y(n_1566) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1543), .Y(n_1567) );
INVxp67_ASAP7_75t_SL g1568 ( .A(n_1534), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1517), .B(n_1481), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1519), .B(n_1481), .Y(n_1570) );
OR2x2_ASAP7_75t_L g1571 ( .A(n_1547), .B(n_1469), .Y(n_1571) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1531), .Y(n_1572) );
A2O1A1Ixp33_ASAP7_75t_L g1573 ( .A1(n_1550), .A2(n_1474), .B(n_1475), .C(n_1472), .Y(n_1573) );
AOI21xp5_ASAP7_75t_L g1574 ( .A1(n_1516), .A2(n_1467), .B(n_1409), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1528), .B(n_1482), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1551), .Y(n_1576) );
NAND3xp33_ASAP7_75t_L g1577 ( .A(n_1539), .B(n_1339), .C(n_1352), .Y(n_1577) );
OAI21xp5_ASAP7_75t_L g1578 ( .A1(n_1518), .A2(n_1415), .B(n_1467), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1540), .Y(n_1579) );
AOI21xp5_ASAP7_75t_L g1580 ( .A1(n_1573), .A2(n_1516), .B(n_1518), .Y(n_1580) );
OAI21xp5_ASAP7_75t_L g1581 ( .A1(n_1573), .A2(n_1515), .B(n_1523), .Y(n_1581) );
AOI21xp5_ASAP7_75t_SL g1582 ( .A1(n_1558), .A2(n_1409), .B(n_1392), .Y(n_1582) );
OAI22xp5_ASAP7_75t_L g1583 ( .A1(n_1574), .A2(n_1532), .B1(n_1533), .B2(n_1527), .Y(n_1583) );
AOI321xp33_ASAP7_75t_L g1584 ( .A1(n_1568), .A2(n_1545), .A3(n_1365), .B1(n_1395), .B2(n_1460), .C(n_1433), .Y(n_1584) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_1571), .A2(n_1532), .B1(n_1524), .B2(n_1541), .Y(n_1585) );
A2O1A1Ixp33_ASAP7_75t_L g1586 ( .A1(n_1578), .A2(n_1525), .B(n_1536), .C(n_1549), .Y(n_1586) );
NAND2xp5_ASAP7_75t_SL g1587 ( .A(n_1577), .B(n_1525), .Y(n_1587) );
INVxp67_ASAP7_75t_L g1588 ( .A(n_1565), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1560), .Y(n_1589) );
OAI22xp5_ASAP7_75t_L g1590 ( .A1(n_1571), .A2(n_1548), .B1(n_1546), .B2(n_1536), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1556), .B(n_1538), .Y(n_1591) );
INVx1_ASAP7_75t_SL g1592 ( .A(n_1554), .Y(n_1592) );
OAI21xp33_ASAP7_75t_L g1593 ( .A1(n_1555), .A2(n_1549), .B(n_1538), .Y(n_1593) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1561), .Y(n_1594) );
OA22x2_ASAP7_75t_L g1595 ( .A1(n_1557), .A2(n_1498), .B1(n_1491), .B2(n_1384), .Y(n_1595) );
AOI222xp33_ASAP7_75t_L g1596 ( .A1(n_1564), .A2(n_1438), .B1(n_1469), .B2(n_1482), .C1(n_1388), .C2(n_1459), .Y(n_1596) );
AOI21xp5_ASAP7_75t_L g1597 ( .A1(n_1570), .A2(n_1498), .B(n_1491), .Y(n_1597) );
AOI32xp33_ASAP7_75t_L g1598 ( .A1(n_1556), .A2(n_1459), .A3(n_1463), .B1(n_1483), .B2(n_1493), .Y(n_1598) );
AOI221xp5_ASAP7_75t_L g1599 ( .A1(n_1580), .A2(n_1563), .B1(n_1562), .B2(n_1567), .C(n_1576), .Y(n_1599) );
OAI221xp5_ASAP7_75t_L g1600 ( .A1(n_1581), .A2(n_1575), .B1(n_1569), .B2(n_1572), .C(n_1579), .Y(n_1600) );
O2A1O1Ixp33_ASAP7_75t_L g1601 ( .A1(n_1588), .A2(n_1364), .B(n_1376), .C(n_1313), .Y(n_1601) );
NOR4xp25_ASAP7_75t_L g1602 ( .A(n_1592), .B(n_1256), .C(n_1559), .D(n_1566), .Y(n_1602) );
OAI22xp33_ASAP7_75t_L g1603 ( .A1(n_1595), .A2(n_1406), .B1(n_1507), .B2(n_1502), .Y(n_1603) );
AOI211xp5_ASAP7_75t_SL g1604 ( .A1(n_1582), .A2(n_1294), .B(n_1266), .C(n_1407), .Y(n_1604) );
O2A1O1Ixp33_ASAP7_75t_SL g1605 ( .A1(n_1586), .A2(n_1579), .B(n_1572), .C(n_1566), .Y(n_1605) );
OAI321xp33_ASAP7_75t_L g1606 ( .A1(n_1583), .A2(n_1553), .A3(n_1407), .B1(n_1436), .B2(n_1494), .C(n_1431), .Y(n_1606) );
BUFx12f_ASAP7_75t_L g1607 ( .A(n_1591), .Y(n_1607) );
NOR2x1_ASAP7_75t_L g1608 ( .A(n_1587), .B(n_1313), .Y(n_1608) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_1584), .A2(n_1552), .B1(n_1364), .B2(n_1376), .C(n_1383), .Y(n_1609) );
OAI311xp33_ASAP7_75t_L g1610 ( .A1(n_1596), .A2(n_1436), .A3(n_1508), .B1(n_1440), .C1(n_1394), .Y(n_1610) );
OAI221xp5_ASAP7_75t_L g1611 ( .A1(n_1595), .A2(n_1540), .B1(n_1497), .B2(n_1490), .C(n_1522), .Y(n_1611) );
AOI221x1_ASAP7_75t_L g1612 ( .A1(n_1585), .A2(n_1398), .B1(n_1353), .B2(n_1354), .C(n_1355), .Y(n_1612) );
NAND4xp25_ASAP7_75t_L g1613 ( .A(n_1604), .B(n_1598), .C(n_1593), .D(n_1257), .Y(n_1613) );
XNOR2xp5_ASAP7_75t_L g1614 ( .A(n_1602), .B(n_1590), .Y(n_1614) );
OAI211xp5_ASAP7_75t_SL g1615 ( .A1(n_1599), .A2(n_1597), .B(n_1594), .C(n_1589), .Y(n_1615) );
NOR2x1p5_ASAP7_75t_L g1616 ( .A(n_1607), .B(n_1257), .Y(n_1616) );
NAND4xp25_ASAP7_75t_L g1617 ( .A(n_1612), .B(n_1384), .C(n_1411), .D(n_1258), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1608), .Y(n_1618) );
NOR3xp33_ASAP7_75t_L g1619 ( .A(n_1606), .B(n_1264), .C(n_1398), .Y(n_1619) );
AOI211xp5_ASAP7_75t_L g1620 ( .A1(n_1603), .A2(n_1411), .B(n_1422), .C(n_1430), .Y(n_1620) );
NAND4xp75_ASAP7_75t_L g1621 ( .A(n_1618), .B(n_1610), .C(n_1600), .D(n_1605), .Y(n_1621) );
NAND3xp33_ASAP7_75t_L g1622 ( .A(n_1614), .B(n_1619), .C(n_1615), .Y(n_1622) );
NAND4xp25_ASAP7_75t_L g1623 ( .A(n_1613), .B(n_1601), .C(n_1611), .D(n_1609), .Y(n_1623) );
NOR3xp33_ASAP7_75t_L g1624 ( .A(n_1617), .B(n_1339), .C(n_1352), .Y(n_1624) );
AOI22x1_ASAP7_75t_L g1625 ( .A1(n_1616), .A2(n_1431), .B1(n_1411), .B2(n_1340), .Y(n_1625) );
NOR3xp33_ASAP7_75t_L g1626 ( .A(n_1620), .B(n_1361), .C(n_1374), .Y(n_1626) );
INVx2_ASAP7_75t_L g1627 ( .A(n_1625), .Y(n_1627) );
NOR2xp67_ASAP7_75t_L g1628 ( .A(n_1623), .B(n_1485), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1622), .B(n_1485), .Y(n_1629) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1621), .Y(n_1630) );
OA22x2_ASAP7_75t_L g1631 ( .A1(n_1630), .A2(n_1624), .B1(n_1626), .B2(n_1437), .Y(n_1631) );
XOR2xp5_ASAP7_75t_L g1632 ( .A(n_1629), .B(n_1431), .Y(n_1632) );
XNOR2x1_ASAP7_75t_L g1633 ( .A(n_1628), .B(n_1267), .Y(n_1633) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1632), .Y(n_1634) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1631), .Y(n_1635) );
AOI222xp33_ASAP7_75t_SL g1636 ( .A1(n_1634), .A2(n_1627), .B1(n_1633), .B2(n_1382), .C1(n_1361), .C2(n_1374), .Y(n_1636) );
OAI21xp33_ASAP7_75t_SL g1637 ( .A1(n_1635), .A2(n_1369), .B(n_1454), .Y(n_1637) );
AOI31xp33_ASAP7_75t_L g1638 ( .A1(n_1637), .A2(n_1379), .A3(n_1377), .B(n_1422), .Y(n_1638) );
AOI22xp33_ASAP7_75t_L g1639 ( .A1(n_1636), .A2(n_1406), .B1(n_1430), .B2(n_1422), .Y(n_1639) );
XNOR2x1_ASAP7_75t_L g1640 ( .A(n_1638), .B(n_1430), .Y(n_1640) );
AOI22xp33_ASAP7_75t_SL g1641 ( .A1(n_1640), .A2(n_1639), .B1(n_1377), .B2(n_1435), .Y(n_1641) );
endmodule