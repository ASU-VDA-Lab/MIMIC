module real_aes_16950_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_119;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g877 ( .A(n_0), .B(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_1), .A2(n_34), .B1(n_132), .B2(n_224), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_2), .A2(n_10), .B1(n_529), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g878 ( .A(n_3), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_4), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_5), .A2(n_11), .B1(n_530), .B2(n_566), .Y(n_565) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_6), .B(n_816), .Y(n_815) );
OR2x2_ASAP7_75t_L g825 ( .A(n_7), .B(n_31), .Y(n_825) );
BUFx2_ASAP7_75t_L g871 ( .A(n_7), .Y(n_871) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_8), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_9), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_12), .B(n_147), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_13), .A2(n_101), .B1(n_177), .B2(n_529), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_14), .A2(n_30), .B1(n_547), .B2(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_15), .B(n_147), .Y(n_544) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_16), .A2(n_47), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_17), .B(n_228), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_18), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_19), .A2(n_38), .B1(n_184), .B2(n_199), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_20), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_21), .A2(n_44), .B1(n_199), .B2(n_529), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_22), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_23), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_24), .B(n_207), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_25), .Y(n_536) );
XNOR2x1_ASAP7_75t_L g816 ( .A(n_26), .B(n_39), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_27), .B(n_125), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_28), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_29), .Y(n_176) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_31), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_32), .A2(n_84), .B1(n_132), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_33), .A2(n_37), .B1(n_132), .B2(n_532), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_35), .A2(n_50), .B1(n_529), .B2(n_584), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_36), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_40), .B(n_147), .Y(n_195) );
INVx2_ASAP7_75t_L g820 ( .A(n_41), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_42), .B(n_180), .Y(n_222) );
BUFx3_ASAP7_75t_L g823 ( .A(n_43), .Y(n_823) );
INVx1_ASAP7_75t_L g837 ( .A(n_43), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_45), .B(n_166), .Y(n_230) );
XOR2x2_ASAP7_75t_L g114 ( .A(n_46), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_46), .A2(n_842), .B1(n_843), .B2(n_846), .Y(n_841) );
INVx1_ASAP7_75t_L g846 ( .A(n_46), .Y(n_846) );
AND2x2_ASAP7_75t_L g258 ( .A(n_48), .B(n_166), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_49), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_51), .B(n_207), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_52), .B(n_184), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_53), .A2(n_70), .B1(n_184), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_54), .A2(n_73), .B1(n_132), .B2(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_55), .B(n_288), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_56), .A2(n_136), .B(n_145), .C(n_251), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_57), .A2(n_98), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g128 ( .A(n_58), .Y(n_128) );
AND2x4_ASAP7_75t_L g150 ( .A(n_59), .B(n_151), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_60), .A2(n_61), .B1(n_199), .B2(n_211), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_62), .A2(n_81), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_62), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_63), .B(n_125), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_64), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_65), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_66), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g151 ( .A(n_67), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_68), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_69), .B(n_125), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_71), .B(n_132), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_72), .B(n_180), .C(n_224), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_74), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_75), .B(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g138 ( .A(n_76), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_77), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_78), .B(n_147), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_79), .B(n_141), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_80), .A2(n_97), .B1(n_145), .B2(n_199), .Y(n_516) );
INVx1_ASAP7_75t_L g845 ( .A(n_81), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_82), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_83), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_85), .A2(n_91), .B1(n_206), .B2(n_207), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_86), .A2(n_105), .B1(n_866), .B2(n_879), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_87), .B(n_147), .Y(n_179) );
NAND2xp33_ASAP7_75t_SL g164 ( .A(n_88), .B(n_135), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_89), .B(n_178), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_90), .B(n_125), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_92), .Y(n_569) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_93), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g828 ( .A(n_94), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g548 ( .A(n_95), .B(n_147), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g134 ( .A(n_96), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_99), .B(n_166), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g160 ( .A(n_100), .B(n_135), .C(n_159), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_102), .B(n_132), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_103), .B(n_207), .Y(n_286) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_817), .B(n_826), .Y(n_105) );
XOR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_814), .Y(n_106) );
AOI21x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_114), .B(n_503), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g503 ( .A(n_109), .B(n_504), .Y(n_503) );
INVx8_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx12f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g864 ( .A(n_112), .B(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g838 ( .A(n_113), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_115), .A2(n_840), .B1(n_841), .B2(n_847), .Y(n_839) );
INVx2_ASAP7_75t_L g847 ( .A(n_115), .Y(n_847) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_435), .Y(n_115) );
NAND4xp25_ASAP7_75t_L g116 ( .A(n_117), .B(n_310), .C(n_350), .D(n_399), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_118), .B(n_259), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_169), .B1(n_231), .B2(n_240), .Y(n_118) );
INVx1_ASAP7_75t_L g431 ( .A(n_119), .Y(n_431) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_120), .B(n_278), .Y(n_347) );
AND2x2_ASAP7_75t_L g378 ( .A(n_120), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_152), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_121), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g302 ( .A(n_121), .Y(n_302) );
AND2x2_ASAP7_75t_L g477 ( .A(n_121), .B(n_345), .Y(n_477) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g242 ( .A(n_122), .Y(n_242) );
AND2x2_ASAP7_75t_L g330 ( .A(n_122), .B(n_292), .Y(n_330) );
AND2x2_ASAP7_75t_L g374 ( .A(n_122), .B(n_279), .Y(n_374) );
OR2x2_ASAP7_75t_L g392 ( .A(n_122), .B(n_393), .Y(n_392) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g296 ( .A(n_123), .B(n_279), .Y(n_296) );
BUFx2_ASAP7_75t_L g353 ( .A(n_123), .Y(n_353) );
OR2x2_ASAP7_75t_L g361 ( .A(n_123), .B(n_319), .Y(n_361) );
INVx1_ASAP7_75t_L g416 ( .A(n_123), .Y(n_416) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx2_ASAP7_75t_L g556 ( .A(n_125), .Y(n_556) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_SL g148 ( .A(n_126), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_SL g155 ( .A(n_126), .Y(n_155) );
INVx2_ASAP7_75t_L g191 ( .A(n_126), .Y(n_191) );
BUFx3_ASAP7_75t_L g512 ( .A(n_126), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_126), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g540 ( .A(n_126), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_126), .B(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_126), .B(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_139), .B(n_148), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_134), .B(n_136), .Y(n_130) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_132), .A2(n_199), .B1(n_256), .B2(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g530 ( .A(n_132), .Y(n_530) );
INVx4_ASAP7_75t_L g532 ( .A(n_132), .Y(n_532) );
INVx1_ASAP7_75t_L g584 ( .A(n_132), .Y(n_584) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_133), .Y(n_135) );
INVx1_ASAP7_75t_L g145 ( .A(n_133), .Y(n_145) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx1_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx1_ASAP7_75t_L g208 ( .A(n_133), .Y(n_208) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
INVx2_ASAP7_75t_L g253 ( .A(n_133), .Y(n_253) );
INVx2_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx1_ASAP7_75t_L g547 ( .A(n_135), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_136), .A2(n_162), .B(n_164), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_136), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_136), .A2(n_283), .B(n_284), .Y(n_282) );
BUFx4f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g143 ( .A(n_138), .Y(n_143) );
INVx1_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
BUFx8_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B1(n_144), .B2(n_146), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_141), .A2(n_182), .B(n_183), .Y(n_181) );
INVx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g213 ( .A(n_143), .Y(n_213) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_147), .A2(n_158), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g228 ( .A(n_147), .Y(n_228) );
INVx3_ASAP7_75t_L g529 ( .A(n_147), .Y(n_529) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_149), .A2(n_157), .B(n_161), .Y(n_156) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_149), .A2(n_175), .B(n_181), .Y(n_174) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_149), .A2(n_193), .B(n_196), .Y(n_192) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_149), .A2(n_221), .B(n_225), .Y(n_220) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_149), .A2(n_282), .B(n_285), .Y(n_281) );
BUFx10_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx10_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
INVx1_ASAP7_75t_L g519 ( .A(n_150), .Y(n_519) );
AND2x2_ASAP7_75t_L g243 ( .A(n_152), .B(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g355 ( .A(n_152), .B(n_332), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_152), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g393 ( .A(n_153), .Y(n_393) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_153), .Y(n_398) );
AND2x2_ASAP7_75t_L g415 ( .A(n_153), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g305 ( .A(n_154), .B(n_245), .Y(n_305) );
INVx1_ASAP7_75t_L g319 ( .A(n_154), .Y(n_319) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_165), .Y(n_154) );
INVx1_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
INVx1_ASAP7_75t_L g517 ( .A(n_159), .Y(n_517) );
INVx1_ASAP7_75t_SL g533 ( .A(n_159), .Y(n_533) );
INVx1_ASAP7_75t_L g575 ( .A(n_163), .Y(n_575) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_167), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_167), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g214 ( .A(n_168), .Y(n_214) );
INVx2_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
NAND2x1_ASAP7_75t_L g169 ( .A(n_170), .B(n_186), .Y(n_169) );
AND2x4_ASAP7_75t_L g480 ( .A(n_170), .B(n_408), .Y(n_480) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_171), .Y(n_239) );
BUFx3_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
INVx1_ASAP7_75t_L g340 ( .A(n_171), .Y(n_340) );
AND2x2_ASAP7_75t_L g343 ( .A(n_171), .B(n_189), .Y(n_343) );
AND2x2_ASAP7_75t_L g368 ( .A(n_171), .B(n_219), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_171), .Y(n_371) );
AND2x2_ASAP7_75t_L g403 ( .A(n_171), .B(n_268), .Y(n_403) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_269) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_173), .A2(n_281), .B(n_290), .Y(n_280) );
OAI21xp33_ASAP7_75t_SL g308 ( .A1(n_173), .A2(n_281), .B(n_290), .Y(n_308) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .C(n_180), .Y(n_175) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_197), .B(n_198), .Y(n_196) );
INVx6_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g542 ( .A1(n_180), .A2(n_532), .B(n_543), .C(n_544), .Y(n_542) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_201), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g312 ( .A(n_188), .B(n_298), .Y(n_312) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g338 ( .A(n_190), .B(n_325), .Y(n_338) );
AND2x2_ASAP7_75t_L g367 ( .A(n_190), .B(n_203), .Y(n_367) );
OR2x2_ASAP7_75t_L g463 ( .A(n_190), .B(n_203), .Y(n_463) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_200), .Y(n_190) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_191), .A2(n_220), .B(n_230), .Y(n_219) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_192), .B(n_200), .Y(n_237) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_191), .A2(n_220), .B(n_230), .Y(n_268) );
INVx2_ASAP7_75t_L g206 ( .A(n_199), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_199), .A2(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g342 ( .A(n_201), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g491 ( .A(n_201), .Y(n_491) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_202), .Y(n_233) );
OR2x2_ASAP7_75t_L g425 ( .A(n_202), .B(n_235), .Y(n_425) );
INVx1_ASAP7_75t_L g447 ( .A(n_202), .Y(n_447) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_219), .Y(n_202) );
AND2x2_ASAP7_75t_L g263 ( .A(n_203), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_268), .Y(n_298) );
INVx1_ASAP7_75t_L g325 ( .A(n_203), .Y(n_325) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_203), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_203), .B(n_219), .Y(n_412) );
AO31x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_214), .A3(n_215), .B(n_216), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_209), .B1(n_210), .B2(n_212), .Y(n_204) );
INVx1_ASAP7_75t_L g566 ( .A(n_207), .Y(n_566) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_209), .A2(n_514), .B1(n_516), .B2(n_517), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_209), .A2(n_528), .B1(n_531), .B2(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_209), .A2(n_546), .B(n_548), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_209), .A2(n_212), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_209), .A2(n_533), .B1(n_565), .B2(n_567), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_209), .A2(n_212), .B1(n_574), .B2(n_576), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_209), .A2(n_212), .B1(n_583), .B2(n_585), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_209), .A2(n_212), .B1(n_599), .B2(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g577 ( .A(n_211), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_212), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g289 ( .A(n_213), .Y(n_289) );
INVx2_ASAP7_75t_L g247 ( .A(n_214), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_214), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_SL g568 ( .A(n_214), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_215), .A2(n_553), .A3(n_556), .B(n_557), .Y(n_552) );
AO31x2_ASAP7_75t_L g563 ( .A1(n_215), .A2(n_526), .A3(n_564), .B(n_568), .Y(n_563) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_215), .A2(n_512), .A3(n_573), .B(n_578), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx2_ASAP7_75t_L g526 ( .A(n_218), .Y(n_526) );
AND2x2_ASAP7_75t_L g349 ( .A(n_219), .B(n_269), .Y(n_349) );
INVx2_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_229), .Y(n_225) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR3x1_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .C(n_238), .Y(n_232) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_235), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g297 ( .A(n_235), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g348 ( .A(n_235), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g388 ( .A(n_235), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_235), .B(n_411), .Y(n_443) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_236), .B(n_324), .Y(n_384) );
AND2x2_ASAP7_75t_L g408 ( .A(n_236), .B(n_268), .Y(n_408) );
BUFx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
BUFx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g419 ( .A(n_239), .B(n_298), .Y(n_419) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_242), .B(n_305), .Y(n_484) );
AND2x4_ASAP7_75t_L g476 ( .A(n_243), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_243), .B(n_296), .Y(n_490) );
INVx2_ASAP7_75t_L g292 ( .A(n_244), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_244), .Y(n_295) );
INVx2_ASAP7_75t_L g380 ( .A(n_244), .Y(n_380) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g364 ( .A(n_245), .Y(n_364) );
AOI21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B(n_258), .Y(n_245) );
NOR2xp67_ASAP7_75t_SL g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g581 ( .A(n_247), .Y(n_581) );
INVx1_ASAP7_75t_L g534 ( .A(n_248), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_SL g515 ( .A(n_253), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_299), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_275), .B1(n_293), .B2(n_297), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_270), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g327 ( .A(n_263), .B(n_274), .Y(n_327) );
AND2x2_ASAP7_75t_L g487 ( .A(n_263), .B(n_368), .Y(n_487) );
BUFx2_ASAP7_75t_L g358 ( .A(n_264), .Y(n_358) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g357 ( .A(n_267), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g272 ( .A(n_268), .Y(n_272) );
INVx1_ASAP7_75t_L g324 ( .A(n_268), .Y(n_324) );
INVx1_ASAP7_75t_L g449 ( .A(n_269), .Y(n_449) );
AOI31xp33_ASAP7_75t_L g467 ( .A1(n_270), .A2(n_468), .A3(n_469), .B(n_470), .Y(n_467) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_272), .B(n_367), .Y(n_466) );
INVx2_ASAP7_75t_L g494 ( .A(n_272), .Y(n_494) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_273), .Y(n_309) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_274), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g452 ( .A(n_274), .B(n_412), .Y(n_452) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_291), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g363 ( .A(n_279), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_289), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx1_ASAP7_75t_L g356 ( .A(n_295), .Y(n_356) );
INVx1_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g397 ( .A(n_296), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g453 ( .A(n_296), .B(n_380), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_297), .A2(n_370), .B(n_372), .Y(n_369) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_309), .Y(n_299) );
NAND3x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .C(n_306), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g471 ( .A(n_302), .B(n_391), .Y(n_471) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2x1_ASAP7_75t_SL g424 ( .A(n_304), .B(n_336), .Y(n_424) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g344 ( .A(n_305), .B(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_306), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_306), .B(n_415), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_306), .B(n_415), .Y(n_488) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g391 ( .A(n_308), .B(n_364), .Y(n_391) );
AND2x2_ASAP7_75t_L g311 ( .A(n_309), .B(n_312), .Y(n_311) );
AOI221x1_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_313), .B1(n_320), .B2(n_329), .C(n_333), .Y(n_310) );
AOI32xp33_ASAP7_75t_L g492 ( .A1(n_312), .A2(n_493), .A3(n_498), .B1(n_499), .B2(n_501), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_317), .B(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_319), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
OR2x2_ASAP7_75t_L g448 ( .A(n_319), .B(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_326), .C(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g370 ( .A(n_323), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g387 ( .A(n_323), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_326), .A2(n_423), .B1(n_425), .B2(n_426), .Y(n_422) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g500 ( .A(n_330), .Y(n_500) );
INVx2_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .B(n_341), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g469 ( .A(n_338), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_339), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_346), .B2(n_348), .Y(n_341) );
AND2x4_ASAP7_75t_L g438 ( .A(n_344), .B(n_353), .Y(n_438) );
INVx1_ASAP7_75t_L g497 ( .A(n_345), .Y(n_497) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g376 ( .A(n_349), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_349), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_349), .B(n_377), .Y(n_468) );
AOI211x1_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_357), .B(n_359), .C(n_385), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR3x2_ASAP7_75t_L g460 ( .A(n_353), .B(n_355), .C(n_356), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_354), .A2(n_376), .B1(n_378), .B2(n_381), .Y(n_375) );
NOR2x1p5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_356), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_355), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_493) );
INVx2_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_365), .B(n_369), .C(n_375), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_367), .B(n_371), .Y(n_382) );
INVx1_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_367), .B(n_474), .Y(n_482) );
OAI32xp33_ASAP7_75t_L g457 ( .A1(n_368), .A2(n_413), .A3(n_458), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g474 ( .A(n_368), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_368), .B(n_388), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_371), .B(n_405), .Y(n_440) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g418 ( .A(n_377), .B(n_403), .Y(n_418) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g427 ( .A(n_380), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g395 ( .A(n_383), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B1(n_394), .B2(n_396), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g414 ( .A(n_391), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_391), .B(n_398), .Y(n_502) );
INVx1_ASAP7_75t_SL g428 ( .A(n_392), .Y(n_428) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_422), .C(n_429), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_413), .B(n_417), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_406), .Y(n_401) );
INVxp67_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .C(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g421 ( .A(n_415), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_423), .A2(n_474), .B1(n_475), .B2(n_478), .C(n_479), .Y(n_473) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI32xp33_ASAP7_75t_L g429 ( .A1(n_426), .A2(n_430), .A3(n_431), .B1(n_432), .B2(n_434), .Y(n_429) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_432), .A2(n_442), .B1(n_443), .B2(n_444), .C(n_450), .Y(n_441) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_454), .C(n_472), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B(n_441), .Y(n_436) );
AOI211x1_ASAP7_75t_L g454 ( .A1(n_437), .A2(n_455), .B(n_457), .C(n_464), .Y(n_454) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2x1_ASAP7_75t_SL g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g456 ( .A(n_447), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AO21x1_ASAP7_75t_L g464 ( .A1(n_453), .A2(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g498 ( .A(n_469), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_485), .Y(n_472) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI21xp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_481), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g495 ( .A(n_494), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND4xp75_ASAP7_75t_L g504 ( .A(n_505), .B(n_654), .C(n_730), .D(n_782), .Y(n_504) );
AND3x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_627), .C(n_640), .Y(n_505) );
AOI221x1_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_559), .B1(n_588), .B2(n_592), .C(n_604), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_507), .A2(n_628), .B(n_630), .C(n_631), .Y(n_627) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_522), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g591 ( .A(n_511), .Y(n_591) );
BUFx2_ASAP7_75t_L g609 ( .A(n_511), .Y(n_609) );
OR2x2_ASAP7_75t_L g651 ( .A(n_511), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g658 ( .A(n_511), .B(n_525), .Y(n_658) );
AND2x4_ASAP7_75t_L g693 ( .A(n_511), .B(n_524), .Y(n_693) );
OR2x2_ASAP7_75t_L g736 ( .A(n_511), .B(n_552), .Y(n_736) );
AO31x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .A3(n_518), .B(n_520), .Y(n_511) );
AO31x2_ASAP7_75t_L g580 ( .A1(n_518), .A2(n_581), .A3(n_582), .B(n_586), .Y(n_580) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_SL g549 ( .A(n_519), .Y(n_549) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_537), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_524), .B(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_524), .Y(n_623) );
INVx2_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
INVx3_ASAP7_75t_L g663 ( .A(n_524), .Y(n_663) );
AND2x2_ASAP7_75t_L g781 ( .A(n_524), .B(n_610), .Y(n_781) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g646 ( .A(n_525), .Y(n_646) );
AO31x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .A3(n_534), .B(n_535), .Y(n_525) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_534), .A2(n_581), .A3(n_598), .B(n_601), .Y(n_597) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g666 ( .A(n_538), .Y(n_666) );
INVx1_ASAP7_75t_L g793 ( .A(n_538), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
AND2x2_ASAP7_75t_L g589 ( .A(n_539), .B(n_552), .Y(n_589) );
INVx1_ASAP7_75t_L g652 ( .A(n_539), .Y(n_652) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_550), .Y(n_539) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_540), .A2(n_541), .B(n_550), .Y(n_611) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B(n_549), .Y(n_541) );
INVx2_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
AND2x2_ASAP7_75t_L g659 ( .A(n_551), .B(n_610), .Y(n_659) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_552), .Y(n_681) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_561), .A2(n_653), .B1(n_657), .B2(n_660), .Y(n_656) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_570), .Y(n_561) );
INVx1_ASAP7_75t_L g674 ( .A(n_562), .Y(n_674) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g594 ( .A(n_563), .B(n_572), .Y(n_594) );
AND2x2_ASAP7_75t_L g625 ( .A(n_563), .B(n_580), .Y(n_625) );
INVx4_ASAP7_75t_SL g636 ( .A(n_563), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_563), .B(n_670), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_563), .B(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g707 ( .A(n_571), .B(n_685), .Y(n_707) );
OR2x2_ASAP7_75t_L g740 ( .A(n_571), .B(n_722), .Y(n_740) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_580), .Y(n_571) );
INVx2_ASAP7_75t_L g614 ( .A(n_572), .Y(n_614) );
INVx1_ASAP7_75t_L g619 ( .A(n_572), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_572), .B(n_596), .Y(n_626) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
INVx1_ASAP7_75t_L g670 ( .A(n_572), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_572), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g603 ( .A(n_580), .Y(n_603) );
AND2x4_ASAP7_75t_L g613 ( .A(n_580), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g639 ( .A(n_580), .Y(n_639) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_580), .Y(n_716) );
INVx1_ASAP7_75t_L g809 ( .A(n_580), .Y(n_809) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_589), .B(n_662), .Y(n_729) );
AND2x2_ASAP7_75t_L g742 ( .A(n_589), .B(n_658), .Y(n_742) );
AND2x2_ASAP7_75t_L g812 ( .A(n_589), .B(n_663), .Y(n_812) );
AND2x4_ASAP7_75t_L g647 ( .A(n_591), .B(n_610), .Y(n_647) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g714 ( .A(n_594), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g728 ( .A(n_594), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_594), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g630 ( .A(n_595), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_595), .B(n_668), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_595), .A2(n_725), .B(n_728), .C(n_729), .Y(n_724) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_603), .Y(n_595) );
AND2x2_ASAP7_75t_L g695 ( .A(n_596), .B(n_636), .Y(n_695) );
INVx3_ASAP7_75t_L g722 ( .A(n_596), .Y(n_722) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g617 ( .A(n_597), .Y(n_617) );
AND2x4_ASAP7_75t_L g643 ( .A(n_597), .B(n_603), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_603), .B(n_636), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_612), .B1(n_620), .B2(n_624), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g761 ( .A(n_606), .Y(n_761) );
AND2x4_ASAP7_75t_L g672 ( .A(n_607), .B(n_652), .Y(n_672) );
INVx1_ASAP7_75t_L g692 ( .A(n_607), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_609), .A2(n_665), .B1(n_675), .B2(n_677), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_609), .B(n_666), .Y(n_723) );
NAND2x1_ASAP7_75t_L g780 ( .A(n_609), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g795 ( .A(n_609), .Y(n_795) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g734 ( .A(n_611), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g653 ( .A(n_613), .B(n_635), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_613), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_613), .B(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_613), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_613), .B(n_676), .Y(n_775) );
AND2x4_ASAP7_75t_L g798 ( .A(n_613), .B(n_726), .Y(n_798) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx3_ASAP7_75t_L g676 ( .A(n_616), .Y(n_676) );
AND2x2_ASAP7_75t_L g688 ( .A(n_616), .B(n_681), .Y(n_688) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g638 ( .A(n_617), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g686 ( .A(n_617), .Y(n_686) );
INVx1_ASAP7_75t_L g629 ( .A(n_618), .Y(n_629) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g786 ( .A(n_619), .B(n_636), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g712 ( .A(n_621), .B(n_693), .Y(n_712) );
INVx2_ASAP7_75t_L g753 ( .A(n_621), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_621), .B(n_647), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_622), .B(n_672), .Y(n_802) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_625), .B(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_L g697 ( .A(n_625), .B(n_642), .Y(n_697) );
INVx1_ASAP7_75t_L g789 ( .A(n_625), .Y(n_789) );
AND2x2_ASAP7_75t_L g788 ( .A(n_626), .B(n_715), .Y(n_788) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_630), .A2(n_760), .B1(n_762), .B2(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_L g668 ( .A(n_636), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g704 ( .A(n_636), .Y(n_704) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_636), .Y(n_710) );
INVx2_ASAP7_75t_L g727 ( .A(n_636), .Y(n_727) );
OR2x2_ASAP7_75t_L g748 ( .A(n_636), .B(n_711), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_636), .B(n_706), .Y(n_758) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g725 ( .A(n_638), .B(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_638), .Y(n_779) );
INVx1_ASAP7_75t_L g706 ( .A(n_639), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B(n_648), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_643), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g711 ( .A(n_643), .Y(n_711) );
AND2x2_ASAP7_75t_L g785 ( .A(n_643), .B(n_786), .Y(n_785) );
AOI211x1_ASAP7_75t_SL g713 ( .A1(n_644), .A2(n_714), .B(n_717), .C(n_724), .Y(n_713) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g770 ( .A(n_646), .B(n_647), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_647), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_647), .Y(n_763) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g678 ( .A(n_650), .Y(n_678) );
NOR2x1p5_ASAP7_75t_L g735 ( .A(n_650), .B(n_736), .Y(n_735) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_651), .B(n_680), .Y(n_679) );
NOR2xp67_ASAP7_75t_SL g752 ( .A(n_651), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g813 ( .A(n_653), .B(n_721), .Y(n_813) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_698), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_664), .C(n_682), .Y(n_655) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_658), .Y(n_689) );
AND2x2_ASAP7_75t_L g696 ( .A(n_658), .B(n_692), .Y(n_696) );
AND2x4_ASAP7_75t_SL g810 ( .A(n_658), .B(n_672), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_661), .A2(n_703), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g792 ( .A(n_663), .B(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_671), .B2(n_673), .Y(n_665) );
NAND2x1_ASAP7_75t_L g741 ( .A(n_668), .B(n_721), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_668), .B(n_715), .Y(n_751) );
INVx1_ASAP7_75t_L g778 ( .A(n_668), .Y(n_778) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_671), .A2(n_797), .B(n_800), .Y(n_796) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_672), .A2(n_684), .B(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g757 ( .A(n_676), .Y(n_757) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g701 ( .A(n_679), .Y(n_701) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_689), .B1(n_690), .B2(n_694), .C1(n_696), .C2(n_697), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_684), .A2(n_718), .B(n_723), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_685), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g799 ( .A(n_685), .Y(n_799) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_686), .Y(n_805) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
AND2x2_ASAP7_75t_L g769 ( .A(n_691), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g762 ( .A(n_692), .B(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_713), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_708), .B2(n_712), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g719 ( .A(n_705), .Y(n_719) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g747 ( .A(n_722), .B(n_739), .Y(n_747) );
OR2x2_ASAP7_75t_L g807 ( .A(n_722), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND5xp2_ASAP7_75t_L g783 ( .A(n_728), .B(n_775), .C(n_784), .D(n_787), .E(n_789), .Y(n_783) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_766), .Y(n_730) );
NAND2xp67_ASAP7_75t_SL g731 ( .A(n_732), .B(n_749), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_737), .B1(n_742), .B2(n_743), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_740), .C(n_741), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g772 ( .A(n_741), .Y(n_772) );
NAND3xp33_ASAP7_75t_SL g743 ( .A(n_744), .B(n_747), .C(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g765 ( .A(n_746), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_SL g777 ( .A1(n_747), .A2(n_778), .B(n_779), .C(n_780), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_754), .B2(n_755), .C(n_759), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_756), .B(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g773 ( .A(n_760), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_771), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g776 ( .A(n_770), .Y(n_776) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_774), .C(n_777), .Y(n_771) );
AOI211x1_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_790), .B(n_796), .C(n_811), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2x1_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B1(n_806), .B2(n_810), .Y(n_800) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx12f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x6_ASAP7_75t_SL g818 ( .A(n_819), .B(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx3_ASAP7_75t_L g832 ( .A(n_820), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_820), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2x1_ASAP7_75t_L g865 ( .A(n_823), .B(n_825), .Y(n_865) );
AND3x2_ASAP7_75t_L g835 ( .A(n_824), .B(n_836), .C(n_838), .Y(n_835) );
AND2x6_ASAP7_75t_SL g851 ( .A(n_824), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_833), .B(n_848), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
OAI31xp33_ASAP7_75t_SL g849 ( .A1(n_828), .A2(n_839), .A3(n_850), .B(n_854), .Y(n_849) );
AOI21xp33_ASAP7_75t_SL g848 ( .A1(n_829), .A2(n_849), .B(n_858), .Y(n_848) );
INVx2_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
BUFx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx8_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_839), .Y(n_833) );
INVx4_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR3xp33_ASAP7_75t_L g875 ( .A(n_836), .B(n_838), .C(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g853 ( .A(n_837), .Y(n_853) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx5_ASAP7_75t_L g857 ( .A(n_851), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_854), .A2(n_859), .B(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
INVx5_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
BUFx10_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx6_ASAP7_75t_L g879 ( .A(n_867), .Y(n_879) );
INVx8_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OR2x6_ASAP7_75t_L g868 ( .A(n_869), .B(n_874), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVxp33_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
endmodule