module real_jpeg_1082_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_54),
.B1(n_56),
.B2(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_39),
.B1(n_54),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_4),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_4),
.B(n_30),
.C(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_33),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_4),
.B(n_54),
.C(n_66),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_4),
.B(n_104),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_4),
.B(n_45),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_4),
.B(n_46),
.C(n_48),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_4),
.B(n_69),
.Y(n_247)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_28),
.B1(n_54),
.B2(n_56),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_172)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_117),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_82),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_82),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_76),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_72),
.B2(n_75),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_129),
.C(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_20),
.A2(n_21),
.B1(n_129),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_20),
.A2(n_21),
.B1(n_93),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_21),
.B(n_93),
.C(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_33),
.B2(n_38),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_30),
.Y(n_32)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_25),
.B(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_35),
.B(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_38),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_59),
.B1(n_60),
.B2(n_71),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_72),
.C(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_71),
.B1(n_77),
.B2(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_57),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_91),
.B(n_108),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_44),
.A2(n_52),
.B1(n_110),
.B2(n_134),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_44),
.A2(n_52),
.B1(n_110),
.B2(n_134),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_44),
.A2(n_52),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_57),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_45)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_48),
.B(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI22x1_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_54),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_69),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_64),
.A2(n_68),
.B(n_81),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_80),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_75),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_72),
.A2(n_75),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_72),
.A2(n_75),
.B1(n_156),
.B2(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_149),
.C(n_156),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_75),
.B(n_129),
.C(n_182),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_96),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_89),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_93),
.B(n_190),
.C(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_93),
.A2(n_174),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_111),
.B(n_112),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_98),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_107),
.B1(n_111),
.B2(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_101),
.B(n_153),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_103),
.A2(n_104),
.B1(n_153),
.B2(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_136),
.B(n_152),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_105),
.A2(n_152),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_137),
.B(n_270),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_119),
.B(n_122),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_145),
.B1(n_182),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_129),
.A2(n_145),
.B1(n_154),
.B2(n_155),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_129),
.B(n_154),
.C(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_131),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_132),
.A2(n_133),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_132),
.A2(n_133),
.B1(n_220),
.B2(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_133),
.B(n_215),
.C(n_220),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_133),
.B(n_171),
.C(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_160),
.B(n_269),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_157),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_141),
.B(n_157),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_148),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_142),
.B(n_146),
.Y(n_267)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_148),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_150),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_154),
.A2(n_155),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_154),
.B(n_241),
.Y(n_249)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_264),
.B(n_268),
.Y(n_160)
);

OAI211xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_193),
.B(n_207),
.C(n_208),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_183),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_175),
.B2(n_176),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_178),
.C(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_171),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_171),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_235),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_189),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_191),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_209),
.C(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_199),
.C(n_205),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21x1_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_226),
.B(n_263),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_214),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_257),
.B(n_262),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_251),
.B(n_256),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_243),
.B(n_250),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_237),
.B(n_242),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_234),
.B(n_236),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_261),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);


endmodule