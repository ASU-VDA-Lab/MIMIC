module fake_jpeg_21512_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_53),
.Y(n_68)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_56),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_37),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_34),
.C(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_67),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_35),
.B1(n_55),
.B2(n_42),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_37),
.B1(n_32),
.B2(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_65),
.Y(n_106)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_39),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_70),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_38),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_16),
.B1(n_32),
.B2(n_21),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_80),
.B1(n_41),
.B2(n_48),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_31),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_28),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_32),
.B1(n_39),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_33),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_84),
.Y(n_110)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_34),
.Y(n_128)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_69),
.B1(n_70),
.B2(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_33),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_57),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_17),
.B1(n_19),
.B2(n_18),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_130),
.B(n_34),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_61),
.B1(n_78),
.B2(n_102),
.Y(n_164)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_117),
.Y(n_153)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_68),
.B(n_69),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_34),
.B(n_24),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_57),
.A3(n_70),
.B1(n_17),
.B2(n_64),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_20),
.C(n_24),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_122),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_34),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_34),
.B(n_36),
.C(n_39),
.Y(n_130)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_66),
.B1(n_77),
.B2(n_75),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_101),
.B1(n_75),
.B2(n_85),
.Y(n_138)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_157),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_144),
.B1(n_34),
.B2(n_29),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_92),
.B1(n_105),
.B2(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_92),
.B1(n_84),
.B2(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_155),
.B1(n_162),
.B2(n_29),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_24),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_148),
.B(n_161),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_109),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_90),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_71),
.C(n_82),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_111),
.C(n_134),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_61),
.B1(n_78),
.B2(n_58),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_166),
.C(n_0),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_132),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_20),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_102),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_111),
.B1(n_125),
.B2(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_90),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_155),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_175),
.Y(n_210)
);

BUFx4f_ASAP7_75t_SL g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_162),
.B(n_141),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_179),
.B(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_185),
.Y(n_205)
);

CKINVDCx10_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_158),
.C(n_160),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_120),
.C(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_131),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_130),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_193),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_117),
.B(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_29),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_30),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_0),
.B(n_30),
.Y(n_218)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_204),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_157),
.B1(n_153),
.B2(n_26),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_189),
.Y(n_228)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_10),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_11),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_11),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_220),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_168),
.B1(n_195),
.B2(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_11),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_197),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_9),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_236),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_176),
.B(n_179),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_230),
.B(n_214),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_184),
.C(n_180),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_191),
.C(n_197),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_170),
.C(n_182),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_208),
.B1(n_209),
.B2(n_207),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_177),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_177),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_203),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_205),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_225),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_226),
.C(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_219),
.B(n_198),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_235),
.B(n_221),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_191),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_218),
.B1(n_170),
.B2(n_199),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_238),
.C(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_224),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_254),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_262),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_228),
.B1(n_208),
.B2(n_215),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_199),
.C(n_215),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_251),
.C(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_252),
.C(n_199),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_251),
.CI(n_254),
.CON(n_270),
.SN(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_278),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_203),
.C(n_250),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_265),
.B1(n_264),
.B2(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_273),
.C(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_204),
.C(n_26),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_276),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_259),
.B(n_1),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_9),
.B(n_1),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_278),
.C(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_25),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_290),
.B(n_291),
.Y(n_294)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_288),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_295),
.A3(n_294),
.B1(n_292),
.B2(n_23),
.C1(n_22),
.C2(n_7),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_6),
.C(n_2),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_7),
.B(n_3),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_4),
.A3(n_6),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_0),
.Y(n_300)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_4),
.B1(n_6),
.B2(n_12),
.C(n_13),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_4),
.B(n_0),
.Y(n_302)
);


endmodule