module fake_jpeg_12046_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_18),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_57),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_26),
.B1(n_24),
.B2(n_38),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_80),
.C(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_85),
.B1(n_28),
.B2(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_74),
.Y(n_99)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_19),
.B(n_36),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_25),
.B(n_34),
.C(n_36),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_37),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_22),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_28),
.B1(n_31),
.B2(n_21),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_55),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_44),
.B1(n_17),
.B2(n_25),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_39),
.B(n_22),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_32),
.B(n_86),
.C(n_55),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_110),
.A2(n_111),
.B1(n_123),
.B2(n_103),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_64),
.A2(n_47),
.B1(n_53),
.B2(n_52),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_95),
.B1(n_44),
.B2(n_59),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_130),
.Y(n_150)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_135),
.Y(n_139)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_87),
.C(n_59),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_44),
.B1(n_53),
.B2(n_52),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_59),
.B1(n_43),
.B2(n_53),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_33),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_134),
.Y(n_159)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_63),
.B(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_20),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_79),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_118),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_73),
.B(n_80),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_166),
.B(n_119),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_160),
.B1(n_165),
.B2(n_167),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_105),
.B(n_61),
.CI(n_82),
.CON(n_146),
.SN(n_146)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_124),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_170),
.B1(n_122),
.B2(n_69),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_52),
.B1(n_41),
.B2(n_51),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_92),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_19),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_103),
.B(n_51),
.C(n_81),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_131),
.C(n_108),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_109),
.A2(n_32),
.B(n_34),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_110),
.B1(n_132),
.B2(n_127),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_124),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_70),
.B1(n_51),
.B2(n_69),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_175),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_151),
.B(n_157),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_185),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_192),
.B1(n_194),
.B2(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_180),
.A2(n_29),
.B(n_30),
.Y(n_224)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_164),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_184),
.C(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_128),
.C(n_129),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_137),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_121),
.B1(n_125),
.B2(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_193),
.B1(n_197),
.B2(n_199),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_202),
.B1(n_204),
.B2(n_155),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_106),
.C(n_100),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_149),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_113),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_125),
.B1(n_121),
.B2(n_20),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_117),
.B1(n_81),
.B2(n_65),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_20),
.B1(n_31),
.B2(n_28),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_43),
.B1(n_93),
.B2(n_76),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_141),
.A2(n_168),
.B1(n_146),
.B2(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_101),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_29),
.C(n_9),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_141),
.A2(n_93),
.B1(n_76),
.B2(n_43),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_120),
.B1(n_115),
.B2(n_114),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_147),
.B1(n_29),
.B2(n_30),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_115),
.B(n_116),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_29),
.B(n_1),
.Y(n_230)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_114),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_86),
.C(n_30),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_29),
.C(n_2),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_166),
.B1(n_152),
.B2(n_142),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_209),
.A2(n_213),
.B(n_221),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_229),
.Y(n_241)
);

AO21x2_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_151),
.B(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_211),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_160),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_232),
.C(n_205),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_138),
.B1(n_158),
.B2(n_86),
.Y(n_213)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_224),
.B(n_225),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_147),
.A3(n_157),
.B1(n_158),
.B2(n_30),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_233),
.B1(n_234),
.B2(n_0),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_180),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_195),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_231),
.B(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_29),
.B(n_1),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_178),
.B1(n_176),
.B2(n_172),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_172),
.A2(n_187),
.B1(n_175),
.B2(n_197),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_182),
.B(n_179),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_184),
.C(n_181),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_242),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_196),
.B1(n_189),
.B2(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_255),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_211),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_260),
.Y(n_262)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_186),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_256),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_10),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_202),
.B1(n_199),
.B2(n_10),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_230),
.B(n_231),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_9),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_206),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_202),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_219),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_244),
.B1(n_246),
.B2(n_245),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_7),
.C(n_14),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_234),
.B1(n_233),
.B2(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_211),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_278),
.B1(n_246),
.B2(n_211),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_224),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_272),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_232),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_213),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.C(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_208),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_211),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_283),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_245),
.B1(n_248),
.B2(n_243),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_288),
.B1(n_280),
.B2(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_238),
.C(n_243),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_294),
.C(n_295),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_245),
.B1(n_238),
.B2(n_242),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_237),
.B(n_209),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_275),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_237),
.B(n_225),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_268),
.B1(n_278),
.B2(n_281),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_240),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_208),
.C(n_209),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_298),
.B(n_305),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_276),
.C(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_303),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_217),
.B1(n_262),
.B2(n_229),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_266),
.C(n_262),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_288),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_292),
.B1(n_294),
.B2(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_295),
.C(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_302),
.B(n_307),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_315),
.B(n_0),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_286),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_296),
.B(n_270),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_283),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_222),
.B1(n_7),
.B2(n_11),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_299),
.B(n_309),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_325),
.B(n_3),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_310),
.C(n_306),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_328),
.B1(n_5),
.B2(n_3),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_326),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_311),
.A2(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_317),
.C(n_315),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_331),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_318),
.B(n_13),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_0),
.C(n_2),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_332),
.A2(n_335),
.B(n_328),
.Y(n_337)
);

NAND4xp25_ASAP7_75t_SL g338 ( 
.A(n_333),
.B(n_334),
.C(n_329),
.D(n_4),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_334),
.C(n_4),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_3),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_340),
.B(n_4),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_4),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_5),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_5),
.Y(n_345)
);


endmodule