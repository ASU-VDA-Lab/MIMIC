module real_aes_7382_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g191 ( .A1(n_0), .A2(n_192), .B(n_193), .C(n_197), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_1), .B(n_187), .Y(n_198) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_3), .B(n_152), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_4), .A2(n_133), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_138), .B(n_143), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_6), .A2(n_133), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_7), .B(n_187), .Y(n_484) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_8), .A2(n_166), .B(n_216), .Y(n_215) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_10), .A2(n_138), .B(n_143), .C(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g539 ( .A(n_11), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_39), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_13), .B(n_196), .Y(n_516) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_15), .B(n_152), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_16), .A2(n_153), .B(n_524), .C(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_17), .B(n_187), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_18), .B(n_180), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_19), .A2(n_143), .B(n_174), .C(n_179), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_20), .A2(n_195), .B(n_210), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_21), .B(n_196), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_22), .A2(n_75), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_22), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_23), .B(n_196), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_24), .Y(n_465) );
INVx1_ASAP7_75t_L g490 ( .A(n_25), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_26), .A2(n_143), .B(n_179), .C(n_219), .Y(n_218) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_28), .Y(n_512) );
INVx1_ASAP7_75t_L g566 ( .A(n_29), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_30), .A2(n_133), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_32), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_33), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_34), .A2(n_195), .B(n_481), .C(n_483), .Y(n_480) );
INVxp67_ASAP7_75t_L g567 ( .A(n_35), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_36), .B(n_221), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_37), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_38), .A2(n_143), .B(n_179), .C(n_489), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_40), .A2(n_197), .B(n_537), .C(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_41), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_42), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_43), .B(n_152), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_44), .B(n_133), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_45), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_46), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_47), .A2(n_141), .B(n_156), .C(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_48), .A2(n_86), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g194 ( .A(n_49), .Y(n_194) );
INVx1_ASAP7_75t_L g231 ( .A(n_50), .Y(n_231) );
INVx1_ASAP7_75t_L g502 ( .A(n_51), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_52), .B(n_133), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_53), .Y(n_183) );
CKINVDCx14_ASAP7_75t_R g535 ( .A(n_54), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_55), .Y(n_447) );
INVx1_ASAP7_75t_L g139 ( .A(n_56), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_57), .B(n_133), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_58), .B(n_187), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_59), .A2(n_178), .B(n_241), .C(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g161 ( .A(n_60), .Y(n_161) );
INVx1_ASAP7_75t_SL g482 ( .A(n_61), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_63), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_64), .B(n_187), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_65), .B(n_153), .Y(n_207) );
INVx1_ASAP7_75t_L g468 ( .A(n_66), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_67), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_68), .B(n_149), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_69), .A2(n_143), .B(n_156), .C(n_267), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_70), .Y(n_239) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_72), .A2(n_133), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_73), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_74), .A2(n_133), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_75), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_76), .A2(n_172), .B(n_562), .Y(n_561) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_77), .Y(n_487) );
INVx1_ASAP7_75t_L g522 ( .A(n_78), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_79), .B(n_148), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_80), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_81), .A2(n_133), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g525 ( .A(n_82), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_83), .Y(n_742) );
INVx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g515 ( .A(n_85), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_86), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_87), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_88), .B(n_196), .Y(n_208) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
OR2x2_ASAP7_75t_L g445 ( .A(n_89), .B(n_111), .Y(n_445) );
OR2x2_ASAP7_75t_L g452 ( .A(n_89), .B(n_112), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_90), .A2(n_143), .B(n_156), .C(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_91), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
INVxp67_ASAP7_75t_L g244 ( .A(n_93), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_94), .B(n_166), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_95), .A2(n_102), .B1(n_115), .B2(n_743), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g203 ( .A(n_97), .Y(n_203) );
INVx1_ASAP7_75t_L g268 ( .A(n_98), .Y(n_268) );
INVx2_ASAP7_75t_L g505 ( .A(n_99), .Y(n_505) );
AND2x2_ASAP7_75t_L g233 ( .A(n_100), .B(n_158), .Y(n_233) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g744 ( .A(n_105), .Y(n_744) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_108), .A2(n_450), .B1(n_732), .B2(n_735), .C1(n_741), .C2(n_742), .Y(n_449) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g455 ( .A(n_110), .B(n_112), .Y(n_455) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21x1_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_120), .B(n_448), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g448 ( .A1(n_116), .A2(n_446), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_443), .B(n_446), .Y(n_120) );
XOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx2_ASAP7_75t_L g453 ( .A(n_125), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_125), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_735) );
OR3x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_357), .C(n_400), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_284), .C(n_314), .D(n_331), .E(n_346), .Y(n_126) );
AOI221xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_199), .B1(n_246), .B2(n_252), .C(n_256), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_168), .Y(n_128) );
OR2x2_ASAP7_75t_L g261 ( .A(n_129), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g301 ( .A(n_129), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_129), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_129), .B(n_254), .Y(n_336) );
OR2x2_ASAP7_75t_L g348 ( .A(n_129), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_129), .B(n_307), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_129), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_129), .B(n_285), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_129), .B(n_293), .Y(n_399) );
AND2x2_ASAP7_75t_L g431 ( .A(n_129), .B(n_185), .Y(n_431) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_129), .Y(n_439) );
INVx5_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_130), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g258 ( .A(n_130), .B(n_234), .Y(n_258) );
BUFx2_ASAP7_75t_L g281 ( .A(n_130), .Y(n_281) );
AND2x2_ASAP7_75t_L g310 ( .A(n_130), .B(n_169), .Y(n_310) );
AND2x2_ASAP7_75t_L g365 ( .A(n_130), .B(n_262), .Y(n_365) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_158), .Y(n_131) );
BUFx2_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_134), .B(n_138), .Y(n_204) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_137), .Y(n_196) );
INVx1_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
INVx4_ASAP7_75t_SL g157 ( .A(n_138), .Y(n_157) );
BUFx3_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_142), .A2(n_157), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_142), .A2(n_157), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_142), .A2(n_157), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_142), .A2(n_157), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_142), .A2(n_157), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_142), .A2(n_157), .B(n_535), .C(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_SL g562 ( .A1(n_142), .A2(n_157), .B(n_563), .C(n_564), .Y(n_562) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_144), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_148), .A2(n_154), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_148), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
O2A1O1Ixp5_ASAP7_75t_L g514 ( .A1(n_148), .A2(n_470), .B(n_515), .C(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g242 ( .A(n_150), .Y(n_242) );
INVx2_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_152), .B(n_244), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_152), .A2(n_177), .B(n_490), .C(n_491), .Y(n_489) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_152), .A2(n_242), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_153), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
INVx1_ASAP7_75t_L g526 ( .A(n_155), .Y(n_526) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g181 ( .A(n_158), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_158), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_158), .A2(n_204), .B(n_487), .C(n_488), .Y(n_486) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_158), .A2(n_533), .B(n_540), .Y(n_532) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g167 ( .A(n_159), .B(n_160), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx3_ASAP7_75t_L g187 ( .A(n_165), .Y(n_187) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_202), .B(n_212), .Y(n_201) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_165), .A2(n_265), .B(n_273), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_165), .B(n_274), .Y(n_273) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_165), .A2(n_464), .B(n_471), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_165), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_165), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_166), .A2(n_217), .B(n_218), .Y(n_216) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_168), .B(n_319), .Y(n_328) );
OAI32xp33_ASAP7_75t_L g342 ( .A1(n_168), .A2(n_278), .A3(n_343), .B1(n_344), .B2(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_168), .B(n_344), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_168), .B(n_261), .Y(n_385) );
INVx1_ASAP7_75t_SL g414 ( .A(n_168), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g423 ( .A(n_168), .B(n_201), .C(n_365), .D(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_185), .Y(n_168) );
INVx5_ASAP7_75t_L g255 ( .A(n_169), .Y(n_255) );
AND2x2_ASAP7_75t_L g285 ( .A(n_169), .B(n_186), .Y(n_285) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_169), .Y(n_364) );
AND2x2_ASAP7_75t_L g434 ( .A(n_169), .B(n_381), .Y(n_434) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
AOI21xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_173), .B(n_180), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_178), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_181), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_184), .A2(n_511), .B(n_517), .Y(n_510) );
AND2x4_ASAP7_75t_L g307 ( .A(n_185), .B(n_255), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_185), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g341 ( .A(n_185), .B(n_262), .Y(n_341) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g254 ( .A(n_186), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g293 ( .A(n_186), .B(n_264), .Y(n_293) );
AND2x2_ASAP7_75t_L g302 ( .A(n_186), .B(n_263), .Y(n_302) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_198), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_195), .B(n_482), .Y(n_481) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g537 ( .A(n_196), .Y(n_537) );
INVx2_ASAP7_75t_L g470 ( .A(n_197), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_199), .A2(n_371), .B1(n_373), .B2(n_375), .C1(n_378), .C2(n_379), .Y(n_370) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_223), .Y(n_199) );
AND2x2_ASAP7_75t_L g303 ( .A(n_200), .B(n_304), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_200), .B(n_281), .C(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_215), .Y(n_200) );
INVx5_ASAP7_75t_SL g251 ( .A(n_201), .Y(n_251) );
OAI322xp33_ASAP7_75t_L g256 ( .A1(n_201), .A2(n_257), .A3(n_259), .B1(n_260), .B2(n_275), .C1(n_278), .C2(n_280), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_201), .B(n_249), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_201), .B(n_235), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_204), .A2(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_204), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_222), .Y(n_219) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx2_ASAP7_75t_L g560 ( .A(n_214), .Y(n_560) );
INVx2_ASAP7_75t_L g249 ( .A(n_215), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_215), .B(n_225), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_223), .B(n_288), .Y(n_343) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g322 ( .A(n_224), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
OR2x2_ASAP7_75t_L g250 ( .A(n_225), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_225), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g290 ( .A(n_225), .B(n_235), .Y(n_290) );
AND2x2_ASAP7_75t_L g313 ( .A(n_225), .B(n_249), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_225), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g329 ( .A(n_225), .B(n_288), .Y(n_329) );
AND2x2_ASAP7_75t_L g337 ( .A(n_225), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_225), .B(n_297), .Y(n_387) );
INVx5_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g277 ( .A(n_226), .B(n_251), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_226), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g304 ( .A(n_226), .B(n_235), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_226), .B(n_351), .Y(n_392) );
OR2x2_ASAP7_75t_L g408 ( .A(n_226), .B(n_352), .Y(n_408) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_226), .B(n_369), .Y(n_415) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_226), .Y(n_422) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
AND2x2_ASAP7_75t_L g276 ( .A(n_234), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g326 ( .A(n_234), .B(n_249), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_234), .B(n_251), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_234), .B(n_288), .Y(n_410) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_235), .B(n_251), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_235), .B(n_249), .Y(n_298) );
OR2x2_ASAP7_75t_L g352 ( .A(n_235), .B(n_249), .Y(n_352) );
AND2x2_ASAP7_75t_L g369 ( .A(n_235), .B(n_248), .Y(n_369) );
INVxp67_ASAP7_75t_L g391 ( .A(n_235), .Y(n_391) );
AND2x2_ASAP7_75t_L g418 ( .A(n_235), .B(n_288), .Y(n_418) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_235), .Y(n_425) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_236), .A2(n_477), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_236), .A2(n_500), .B(n_506), .Y(n_499) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_236), .A2(n_520), .B(n_527), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_241), .A2(n_268), .B(n_269), .C(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_242), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_242), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_248), .B(n_299), .Y(n_372) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g288 ( .A(n_249), .B(n_251), .Y(n_288) );
OR2x2_ASAP7_75t_L g355 ( .A(n_249), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
OR2x2_ASAP7_75t_L g360 ( .A(n_250), .B(n_352), .Y(n_360) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g259 ( .A(n_254), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_254), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g260 ( .A(n_255), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_255), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_255), .B(n_262), .Y(n_295) );
INVx2_ASAP7_75t_L g340 ( .A(n_255), .Y(n_340) );
AND2x2_ASAP7_75t_L g353 ( .A(n_255), .B(n_293), .Y(n_353) );
AND2x2_ASAP7_75t_L g378 ( .A(n_255), .B(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
INVx2_ASAP7_75t_SL g317 ( .A(n_261), .Y(n_317) );
INVx1_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx2_ASAP7_75t_L g381 ( .A(n_264), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_272), .Y(n_265) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g483 ( .A(n_271), .Y(n_483) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g350 ( .A(n_277), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g356 ( .A(n_277), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_277), .A2(n_359), .B1(n_361), .B2(n_366), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_277), .B(n_369), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_278), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g312 ( .A(n_279), .Y(n_312) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
OR2x2_ASAP7_75t_L g294 ( .A(n_281), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_281), .B(n_285), .Y(n_345) );
AND2x2_ASAP7_75t_L g368 ( .A(n_281), .B(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_291), .C(n_305), .Y(n_284) );
INVx1_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_285), .A2(n_417), .B1(n_419), .B2(n_420), .C(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g435 ( .A(n_288), .Y(n_435) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g384 ( .A(n_290), .B(n_323), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_296), .C(n_300), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OAI32xp33_ASAP7_75t_L g409 ( .A1(n_298), .A2(n_299), .A3(n_362), .B1(n_399), .B2(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_L g441 ( .A(n_301), .B(n_340), .Y(n_441) );
AND2x2_ASAP7_75t_L g388 ( .A(n_302), .B(n_340), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_302), .B(n_310), .Y(n_406) );
AOI31xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_308), .A3(n_309), .B(n_311), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_307), .B(n_319), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_307), .B(n_317), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_307), .A2(n_337), .B1(n_427), .B2(n_430), .C(n_432), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g332 ( .A(n_312), .B(n_333), .Y(n_332) );
AOI222xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_321), .B1(n_324), .B2(n_327), .C1(n_329), .C2(n_330), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g397 ( .A(n_316), .Y(n_397) );
INVx1_ASAP7_75t_L g419 ( .A(n_319), .Y(n_419) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_322), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g338 ( .A(n_323), .Y(n_338) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B1(n_337), .B2(n_339), .C(n_342), .Y(n_331) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g428 ( .A(n_334), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
INVx1_ASAP7_75t_L g349 ( .A(n_341), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_344), .B(n_431), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B1(n_353), .B2(n_354), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g440 ( .A(n_353), .Y(n_440) );
INVxp33_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_355), .B(n_399), .Y(n_398) );
OAI32xp33_ASAP7_75t_L g389 ( .A1(n_356), .A2(n_390), .A3(n_391), .B1(n_392), .B2(n_393), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_370), .C(n_382), .D(n_394), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NAND2xp33_ASAP7_75t_SL g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_365), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_379), .A2(n_395), .B1(n_412), .B2(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g430 ( .A(n_381), .B(n_431), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B1(n_386), .B2(n_388), .C(n_389), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_391), .B(n_422), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_411), .C(n_426), .D(n_437), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B(n_407), .C(n_409), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g442 ( .A(n_429), .Y(n_442) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B(n_442), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_445), .B(n_447), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_456), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g738 ( .A(n_452), .Y(n_738) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_L g739 ( .A(n_455), .Y(n_739) );
INVx3_ASAP7_75t_L g740 ( .A(n_456), .Y(n_740) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_687), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_624), .C(n_658), .D(n_674), .Y(n_457) );
NAND4xp25_ASAP7_75t_SL g458 ( .A(n_459), .B(n_553), .C(n_588), .D(n_604), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_494), .B1(n_528), .B2(n_541), .C1(n_546), .C2(n_552), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g720 ( .A1(n_461), .A2(n_721), .A3(n_722), .B(n_724), .Y(n_720) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
AND2x2_ASAP7_75t_L g695 ( .A(n_462), .B(n_475), .Y(n_695) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g545 ( .A(n_463), .Y(n_545) );
AND2x2_ASAP7_75t_L g552 ( .A(n_463), .B(n_485), .Y(n_552) );
AND2x2_ASAP7_75t_L g609 ( .A(n_463), .B(n_476), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_473), .B(n_639), .Y(n_638) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_474), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_474), .B(n_556), .Y(n_599) );
AND2x2_ASAP7_75t_L g692 ( .A(n_474), .B(n_632), .Y(n_692) );
OAI321xp33_ASAP7_75t_L g726 ( .A1(n_474), .A2(n_545), .A3(n_699), .B1(n_727), .B2(n_729), .C(n_730), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_474), .B(n_531), .C(n_639), .D(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
AND2x2_ASAP7_75t_L g594 ( .A(n_475), .B(n_543), .Y(n_594) );
AND2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_545), .Y(n_613) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g544 ( .A(n_476), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g569 ( .A(n_476), .B(n_485), .Y(n_569) );
AND2x2_ASAP7_75t_L g655 ( .A(n_476), .B(n_543), .Y(n_655) );
INVx3_ASAP7_75t_SL g543 ( .A(n_485), .Y(n_543) );
AND2x2_ASAP7_75t_L g587 ( .A(n_485), .B(n_574), .Y(n_587) );
OR2x2_ASAP7_75t_L g620 ( .A(n_485), .B(n_545), .Y(n_620) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_485), .Y(n_627) );
AND2x2_ASAP7_75t_L g656 ( .A(n_485), .B(n_544), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_485), .B(n_629), .Y(n_671) );
AND2x2_ASAP7_75t_L g703 ( .A(n_485), .B(n_695), .Y(n_703) );
AND2x2_ASAP7_75t_L g712 ( .A(n_485), .B(n_557), .Y(n_712) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
INVx1_ASAP7_75t_SL g680 ( .A(n_496), .Y(n_680) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g548 ( .A(n_497), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g530 ( .A(n_498), .B(n_509), .Y(n_530) );
AND2x2_ASAP7_75t_L g616 ( .A(n_498), .B(n_532), .Y(n_616) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g586 ( .A(n_499), .B(n_519), .Y(n_586) );
OR2x2_ASAP7_75t_L g597 ( .A(n_499), .B(n_532), .Y(n_597) );
AND2x2_ASAP7_75t_L g623 ( .A(n_499), .B(n_532), .Y(n_623) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_499), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_507), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_507), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g596 ( .A(n_508), .B(n_597), .Y(n_596) );
AOI322xp5_ASAP7_75t_L g682 ( .A1(n_508), .A2(n_586), .A3(n_592), .B1(n_623), .B2(n_673), .C1(n_683), .C2(n_685), .Y(n_682) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_519), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_509), .B(n_531), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_509), .B(n_532), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_509), .B(n_549), .Y(n_603) );
AND2x2_ASAP7_75t_L g657 ( .A(n_509), .B(n_623), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_509), .Y(n_661) );
AND2x2_ASAP7_75t_L g673 ( .A(n_509), .B(n_519), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_509), .B(n_548), .Y(n_705) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g570 ( .A(n_510), .B(n_519), .Y(n_570) );
BUFx3_ASAP7_75t_L g584 ( .A(n_510), .Y(n_584) );
AND3x2_ASAP7_75t_L g666 ( .A(n_510), .B(n_646), .C(n_667), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_519), .B(n_530), .C(n_531), .Y(n_529) );
INVx1_ASAP7_75t_SL g549 ( .A(n_519), .Y(n_549) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_519), .Y(n_651) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g645 ( .A(n_530), .B(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g652 ( .A(n_530), .Y(n_652) );
AND2x2_ASAP7_75t_L g690 ( .A(n_531), .B(n_668), .Y(n_690) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
AND2x2_ASAP7_75t_L g646 ( .A(n_532), .B(n_549), .Y(n_646) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
OR2x2_ASAP7_75t_L g590 ( .A(n_543), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g709 ( .A(n_543), .B(n_609), .Y(n_709) );
AND2x2_ASAP7_75t_L g723 ( .A(n_543), .B(n_545), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_544), .B(n_557), .Y(n_664) );
AND2x2_ASAP7_75t_L g711 ( .A(n_544), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g574 ( .A(n_545), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g591 ( .A(n_545), .B(n_557), .Y(n_591) );
INVx1_ASAP7_75t_L g601 ( .A(n_545), .Y(n_601) );
AND2x2_ASAP7_75t_L g632 ( .A(n_545), .B(n_557), .Y(n_632) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_547), .A2(n_675), .B1(n_679), .B2(n_681), .C(n_682), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g578 ( .A(n_548), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_551), .B(n_585), .Y(n_728) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_570), .A3(n_571), .B1(n_572), .B2(n_578), .C1(n_580), .C2(n_587), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_556), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_556), .B(n_619), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_556), .A2(n_569), .B(n_643), .C(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_556), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_556), .B(n_613), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_556), .B(n_695), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_556), .B(n_723), .Y(n_722) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_557), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_557), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g684 ( .A(n_557), .B(n_571), .Y(n_684) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_568), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_559), .A2(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g576 ( .A(n_561), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_568), .Y(n_577) );
INVx1_ASAP7_75t_L g659 ( .A(n_569), .Y(n_659) );
OAI31xp33_ASAP7_75t_L g669 ( .A1(n_569), .A2(n_594), .A3(n_670), .B(n_672), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_569), .B(n_575), .Y(n_721) );
INVx1_ASAP7_75t_SL g582 ( .A(n_570), .Y(n_582) );
AND2x2_ASAP7_75t_L g615 ( .A(n_570), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g696 ( .A(n_570), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g581 ( .A(n_571), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
AND2x2_ASAP7_75t_L g633 ( .A(n_571), .B(n_586), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_571), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g725 ( .A(n_571), .B(n_673), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_573), .B(n_643), .Y(n_716) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g612 ( .A(n_575), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g630 ( .A(n_575), .Y(n_630) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_581), .B(n_583), .Y(n_580) );
OAI211xp5_ASAP7_75t_SL g624 ( .A1(n_582), .A2(n_625), .B(n_631), .C(n_647), .Y(n_624) );
OR2x2_ASAP7_75t_L g699 ( .A(n_582), .B(n_680), .Y(n_699) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_584), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_584), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g605 ( .A(n_586), .B(n_606), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_595), .C(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g639 ( .A(n_591), .Y(n_639) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_594), .B(n_632), .Y(n_637) );
INVx1_ASAP7_75t_L g643 ( .A(n_594), .Y(n_643) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g602 ( .A(n_597), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g635 ( .A(n_597), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g697 ( .A(n_597), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B(n_602), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_600), .A2(n_611), .B(n_614), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B(n_610), .C(n_617), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_605), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_608), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g621 ( .A(n_609), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_611), .A2(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_616), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g641 ( .A(n_616), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_621), .B(n_622), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g672 ( .A(n_623), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_629), .B(n_655), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_629), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g708 ( .A(n_629), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g718 ( .A(n_629), .B(n_656), .Y(n_718) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_634), .C(n_642), .Y(n_631) );
INVx1_ASAP7_75t_L g678 ( .A(n_632), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_638), .B2(n_640), .Y(n_634) );
OR2x2_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_636), .B(n_697), .Y(n_719) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g713 ( .A(n_646), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_653), .B1(n_656), .B2(n_657), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g731 ( .A(n_651), .Y(n_731) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g677 ( .A(n_655), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B(n_662), .C(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_677), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NOR5xp2_ASAP7_75t_L g687 ( .A(n_688), .B(n_706), .C(n_714), .D(n_720), .E(n_726), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_691), .B(n_693), .C(n_700), .Y(n_688) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_698), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_703), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B(n_713), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g729 ( .A(n_709), .Y(n_729) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_732), .Y(n_741) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
endmodule