module fake_netlist_6_1826_n_655 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_655);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_655;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_625;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_229;
wire n_542;
wire n_644;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_624;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_612;
wire n_633;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_151;
wire n_412;
wire n_640;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_17),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_58),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_65),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_19),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_49),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_77),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_93),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_15),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_27),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_28),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_0),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_8),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_42),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_29),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_52),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_97),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_23),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_45),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_63),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_55),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_53),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_132),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_24),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_12),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_120),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_36),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_11),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_115),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_104),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_22),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_86),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_173),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

CKINVDCx6p67_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_1),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_2),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_2),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_3),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_140),
.B(n_3),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_4),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_135),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_143),
.B(n_144),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_4),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_13),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_5),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_5),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_6),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_7),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

BUFx8_ASAP7_75t_SL g245 ( 
.A(n_151),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_175),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_7),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_139),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_142),
.B(n_8),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_201),
.B1(n_199),
.B2(n_146),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_148),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_198),
.B1(n_179),
.B2(n_194),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_196),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_250),
.A2(n_190),
.B1(n_186),
.B2(n_185),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g257 ( 
.A1(n_205),
.A2(n_183),
.B1(n_182),
.B2(n_181),
.Y(n_257)
);

NOR2x1p5_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_149),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

OR2x6_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_9),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_150),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_212),
.A2(n_180),
.B1(n_178),
.B2(n_177),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_10),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_171),
.B1(n_170),
.B2(n_168),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_166),
.B1(n_164),
.B2(n_162),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_152),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_159),
.B1(n_157),
.B2(n_153),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_160),
.B1(n_18),
.B2(n_20),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_16),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_R g278 ( 
.A1(n_213),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_31),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_35),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_212),
.A2(n_216),
.B1(n_215),
.B2(n_242),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_40),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_41),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_43),
.Y(n_286)
);

OR2x6_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_216),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_233),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_233),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_228),
.B(n_61),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_62),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_219),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_242),
.A2(n_236),
.B1(n_237),
.B2(n_251),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_64),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_206),
.B(n_66),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_236),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_211),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_232),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_246),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_245),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_266),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_287),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_273),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_229),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_291),
.B(n_208),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_234),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_217),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_211),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_234),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_260),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_229),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

BUFx6f_ASAP7_75t_SL g334 ( 
.A(n_281),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g336 ( 
.A(n_289),
.B(n_217),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_253),
.B(n_208),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_279),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_234),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_208),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_275),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_262),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_252),
.B(n_78),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_231),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_231),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_269),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_256),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_265),
.B(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_278),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_266),
.B(n_221),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_304),
.B(n_231),
.Y(n_369)
);

XNOR2x2_ASAP7_75t_L g370 ( 
.A(n_262),
.B(n_80),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_272),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_372),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_221),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_81),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_223),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_223),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_350),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_309),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_221),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_220),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_305),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_339),
.B(n_223),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_325),
.B(n_310),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_320),
.B(n_220),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_358),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_366),
.B(n_82),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_366),
.B(n_84),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_306),
.B(n_87),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_222),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_356),
.B(n_222),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_363),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_222),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_344),
.B(n_209),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_209),
.Y(n_416)
);

BUFx8_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

AND2x4_ASAP7_75t_SL g418 ( 
.A(n_363),
.B(n_90),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_209),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_91),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_327),
.B(n_92),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_94),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_361),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_367),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_95),
.Y(n_427)
);

INVx3_ASAP7_75t_SL g428 ( 
.A(n_336),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_355),
.B(n_353),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_98),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_340),
.A2(n_99),
.B(n_100),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_331),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_336),
.B(n_101),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_393),
.B(n_322),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_365),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_391),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_373),
.B(n_362),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_349),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_322),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

OR2x6_ASAP7_75t_SL g452 ( 
.A(n_385),
.B(n_370),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_382),
.B(n_369),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_307),
.Y(n_455)
);

BUFx6f_ASAP7_75t_SL g456 ( 
.A(n_389),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_373),
.B(n_364),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_378),
.B(n_364),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_429),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_374),
.B(n_330),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_378),
.B(n_334),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_354),
.Y(n_467)
);

NAND2x1p5_ASAP7_75t_L g468 ( 
.A(n_414),
.B(n_338),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_428),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_374),
.B(n_330),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_368),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_316),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_436),
.B(n_338),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_434),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_417),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_368),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_378),
.B(n_316),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_449),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_428),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_440),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_461),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_449),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_397),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_460),
.A2(n_435),
.B1(n_405),
.B2(n_403),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_455),
.Y(n_496)
);

BUFx4_ASAP7_75t_SL g497 ( 
.A(n_482),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_442),
.B(n_414),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_472),
.B(n_435),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_453),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_448),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

BUFx8_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

CKINVDCx8_ASAP7_75t_R g508 ( 
.A(n_471),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_459),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_475),
.Y(n_511)
);

INVx3_ASAP7_75t_SL g512 ( 
.A(n_470),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_436),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

CKINVDCx11_ASAP7_75t_R g515 ( 
.A(n_512),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_505),
.Y(n_516)
);

NAND2x1p5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_442),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_450),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_452),
.B1(n_481),
.B2(n_465),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_450),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_503),
.A2(n_472),
.B1(n_467),
.B2(n_403),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

CKINVDCx6p67_ASAP7_75t_R g523 ( 
.A(n_489),
.Y(n_523)
);

CKINVDCx11_ASAP7_75t_R g524 ( 
.A(n_508),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_487),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_494),
.A2(n_405),
.B1(n_460),
.B2(n_396),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_460),
.B1(n_396),
.B2(n_459),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_510),
.A2(n_460),
.B1(n_427),
.B2(n_454),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_486),
.A2(n_481),
.B1(n_456),
.B2(n_418),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_487),
.B(n_511),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_490),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_510),
.A2(n_481),
.B1(n_476),
.B2(n_414),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_495),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_488),
.A2(n_427),
.B1(n_480),
.B2(n_432),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_L g538 ( 
.A1(n_488),
.A2(n_480),
.B1(n_441),
.B2(n_443),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_513),
.B(n_477),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_499),
.B(n_401),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_409),
.B1(n_418),
.B2(n_466),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_516),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_530),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_532),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_537),
.B(n_477),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_425),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_519),
.A2(n_501),
.B1(n_509),
.B2(n_407),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_478),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_526),
.A2(n_496),
.B1(n_478),
.B2(n_381),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_519),
.A2(n_466),
.B1(n_390),
.B2(n_493),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_535),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_523),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_526),
.A2(n_423),
.B(n_424),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_537),
.A2(n_409),
.B1(n_466),
.B2(n_408),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_532),
.Y(n_558)
);

BUFx4f_ASAP7_75t_SL g559 ( 
.A(n_522),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_520),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_534),
.A2(n_507),
.B1(n_466),
.B2(n_482),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_538),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_515),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_538),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_529),
.B(n_446),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

NOR2x1_ASAP7_75t_R g567 ( 
.A(n_525),
.B(n_497),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_517),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_527),
.A2(n_466),
.B1(n_408),
.B2(n_404),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_536),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_528),
.B(n_513),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_542),
.A2(n_527),
.B1(n_528),
.B2(n_439),
.Y(n_573)
);

AOI221xp5_ASAP7_75t_L g574 ( 
.A1(n_551),
.A2(n_410),
.B1(n_437),
.B2(n_419),
.C(n_539),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_548),
.A2(n_439),
.B1(n_539),
.B2(n_384),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_387),
.B1(n_384),
.B2(n_399),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_549),
.B(n_430),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_553),
.A2(n_468),
.B1(n_511),
.B2(n_536),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_565),
.A2(n_491),
.B1(n_430),
.B2(n_468),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_542),
.A2(n_493),
.B1(n_531),
.B2(n_434),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_562),
.A2(n_387),
.B1(n_402),
.B2(n_398),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_557),
.A2(n_506),
.B1(n_495),
.B2(n_517),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_564),
.A2(n_404),
.B1(n_399),
.B2(n_402),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_413),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_557),
.A2(n_398),
.B1(n_412),
.B2(n_406),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_546),
.A2(n_561),
.B1(n_547),
.B2(n_572),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_546),
.A2(n_412),
.B1(n_406),
.B2(n_433),
.Y(n_587)
);

AOI222xp33_ASAP7_75t_L g588 ( 
.A1(n_570),
.A2(n_377),
.B1(n_437),
.B2(n_413),
.C1(n_422),
.C2(n_433),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_558),
.A2(n_487),
.B1(n_420),
.B2(n_502),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_569),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_556),
.A2(n_416),
.B(n_415),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_570),
.A2(n_506),
.B1(n_502),
.B2(n_436),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_572),
.A2(n_421),
.B1(n_431),
.B2(n_400),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_550),
.A2(n_559),
.B1(n_545),
.B2(n_555),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_586),
.A2(n_563),
.B(n_552),
.Y(n_596)
);

AOI221xp5_ASAP7_75t_L g597 ( 
.A1(n_584),
.A2(n_554),
.B1(n_544),
.B2(n_543),
.C(n_377),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_594),
.B(n_568),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_571),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_595),
.A2(n_567),
.B(n_559),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_569),
.C(n_555),
.Y(n_601)
);

OAI221xp5_ASAP7_75t_L g602 ( 
.A1(n_579),
.A2(n_550),
.B1(n_431),
.B2(n_421),
.C(n_571),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_573),
.A2(n_566),
.B1(n_400),
.B2(n_569),
.Y(n_603)
);

NAND4xp25_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_379),
.C(n_400),
.D(n_444),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_569),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_492),
.C(n_483),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_492),
.C(n_483),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_457),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_578),
.B(n_457),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_588),
.B(n_463),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_580),
.C(n_589),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_598),
.B(n_591),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_605),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_591),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_609),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_608),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_596),
.B(n_582),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_588),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_613),
.B(n_600),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_603),
.C(n_602),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_616),
.B(n_606),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_613),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_616),
.B(n_607),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_614),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_615),
.B(n_610),
.Y(n_625)
);

XOR2x2_ASAP7_75t_L g626 ( 
.A(n_621),
.B(n_617),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_622),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_612),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_618),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_624),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_627),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_629),
.Y(n_632)
);

OA22x2_ASAP7_75t_L g633 ( 
.A1(n_630),
.A2(n_623),
.B1(n_624),
.B2(n_620),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_626),
.A2(n_624),
.B1(n_604),
.B2(n_587),
.Y(n_634)
);

XOR2x2_ASAP7_75t_L g635 ( 
.A(n_630),
.B(n_479),
.Y(n_635)
);

OA22x2_ASAP7_75t_L g636 ( 
.A1(n_634),
.A2(n_628),
.B1(n_497),
.B2(n_479),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_631),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_632),
.Y(n_638)
);

NAND4xp25_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_633),
.C(n_635),
.D(n_583),
.Y(n_639)
);

AOI221xp5_ASAP7_75t_L g640 ( 
.A1(n_637),
.A2(n_592),
.B1(n_585),
.B2(n_593),
.C(n_492),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_639),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_641),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_642),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_636),
.B1(n_640),
.B2(n_483),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

NAND4xp25_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_458),
.C(n_451),
.D(n_475),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

AO22x2_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_463),
.B1(n_380),
.B2(n_376),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_648),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_469),
.B1(n_458),
.B2(n_451),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_649),
.A2(n_380),
.B1(n_106),
.B2(n_108),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_650),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_651),
.Y(n_653)
);

AOI221xp5_ASAP7_75t_L g654 ( 
.A1(n_653),
.A2(n_652),
.B1(n_111),
.B2(n_112),
.C(n_116),
.Y(n_654)
);

AOI211xp5_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_655)
);


endmodule