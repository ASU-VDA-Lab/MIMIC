module fake_ibex_1041_n_2718 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_502, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2718);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_502;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2718;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_530;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_709;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_510;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_1894;
wire n_2110;
wire n_1349;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_1380;
wire n_647;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2698;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1946;
wire n_1726;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_786;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2714;
wire n_2669;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2303;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_2704;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx2_ASAP7_75t_L g503 ( 
.A(n_153),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_362),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_78),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_57),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_424),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_37),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_11),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_207),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_181),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_48),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_398),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_355),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_30),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_41),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_162),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_60),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_493),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_297),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_129),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_274),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_233),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_405),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_345),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_240),
.B(n_496),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_55),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_440),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_499),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_126),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_480),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_112),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_120),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_404),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_12),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_335),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_338),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_81),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_221),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_107),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_375),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_125),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_356),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_314),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_70),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_71),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_189),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_408),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_173),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_39),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_410),
.B(n_402),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_351),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_19),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_327),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_81),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_331),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_469),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_150),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_381),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_333),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_67),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_296),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_69),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_501),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_48),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_140),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_439),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_111),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_460),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_445),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_353),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_179),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_313),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_354),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_203),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_140),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_268),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_326),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_301),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_43),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_400),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_271),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_429),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_235),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_256),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_57),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_230),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_382),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_360),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_248),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_231),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_267),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_50),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_434),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_284),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_219),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_37),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_198),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_64),
.Y(n_602)
);

INVxp33_ASAP7_75t_R g603 ( 
.A(n_30),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_359),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_261),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_427),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_23),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_201),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_99),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_218),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_107),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_156),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_97),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_350),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_486),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_227),
.B(n_390),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_259),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_374),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_292),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_311),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_272),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_210),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_491),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_256),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_420),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_442),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_260),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_392),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_329),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_275),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_330),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_304),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_187),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_218),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_306),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_295),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_83),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_443),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_299),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_368),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_106),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_448),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_426),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_456),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_394),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_130),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_370),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_492),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_162),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_425),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_441),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_9),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_236),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_245),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_298),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_254),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_66),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_254),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_444),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_38),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_323),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_447),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_238),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_23),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_47),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_418),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_319),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_177),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_28),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_485),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_183),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_194),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_393),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_233),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_415),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_377),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_307),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_224),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_148),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_243),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_437),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_159),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_5),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_478),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_257),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_321),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_320),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_45),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_282),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_52),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_462),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_148),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_436),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_71),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_371),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_260),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_310),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_389),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_13),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_397),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_102),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_230),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_433),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_303),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_32),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_364),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_168),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_236),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_204),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_244),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_158),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_385),
.B(n_204),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_387),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_358),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_44),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_153),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_461),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_0),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_317),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_251),
.Y(n_721)
);

XOR2xp5_ASAP7_75t_R g722 ( 
.A(n_498),
.B(n_315),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_188),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_56),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_175),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_200),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_108),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_383),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_302),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_477),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_252),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_352),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_463),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_283),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_189),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_190),
.Y(n_736)
);

XOR2xp5_ASAP7_75t_L g737 ( 
.A(n_160),
.B(n_51),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_110),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_235),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_487),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_126),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_168),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_341),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_278),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_294),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_139),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_0),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_18),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_470),
.Y(n_749)
);

CKINVDCx11_ASAP7_75t_R g750 ( 
.A(n_73),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_157),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_399),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_118),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_231),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_15),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_395),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_13),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_269),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_472),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_305),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_278),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_40),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_401),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_340),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_104),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_386),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_367),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_243),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_471),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_170),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_50),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_164),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_452),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_293),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_59),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_154),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_43),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_24),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_110),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_134),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_450),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_421),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_407),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_438),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_141),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_89),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_379),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_123),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_312),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_432),
.Y(n_790)
);

BUFx5_ASAP7_75t_L g791 ( 
.A(n_357),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_44),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_114),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_67),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_222),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_363),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_220),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_98),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_114),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_102),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_476),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_135),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_199),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_10),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_451),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_122),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_26),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_483),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_267),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_490),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_344),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_376),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_184),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_328),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_489),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_40),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_34),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_64),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_198),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_203),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_179),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_121),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_227),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_125),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_369),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_134),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_8),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_116),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_46),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_342),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_273),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_271),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_361),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_184),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_193),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_422),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_300),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_403),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_115),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_282),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_34),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_414),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_378),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_39),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_409),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_259),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_166),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_86),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_208),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_89),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_417),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_481),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_121),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_488),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_459),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_449),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_568),
.B(n_1),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_791),
.Y(n_858)
);

BUFx8_ASAP7_75t_SL g859 ( 
.A(n_539),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_791),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_582),
.B(n_1),
.Y(n_861)
);

CKINVDCx6p67_ASAP7_75t_R g862 ( 
.A(n_542),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_564),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_835),
.B(n_2),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_791),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_670),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_547),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_670),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_683),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_546),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_546),
.Y(n_872)
);

INVx5_ASAP7_75t_L g873 ( 
.A(n_542),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_564),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_703),
.B(n_798),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_561),
.A2(n_286),
.B(n_285),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_564),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_568),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_520),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_638),
.Y(n_880)
);

BUFx8_ASAP7_75t_SL g881 ( 
.A(n_539),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_638),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_564),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_542),
.Y(n_884)
);

OAI22x1_ASAP7_75t_R g885 ( 
.A1(n_540),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_601),
.Y(n_886)
);

BUFx12f_ASAP7_75t_L g887 ( 
.A(n_750),
.Y(n_887)
);

OAI22x1_ASAP7_75t_L g888 ( 
.A1(n_737),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_586),
.B(n_7),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_624),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_533),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_791),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_624),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_653),
.B(n_9),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_749),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_624),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_624),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_673),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_555),
.Y(n_899)
);

NOR2x1_ASAP7_75t_L g900 ( 
.A(n_681),
.B(n_287),
.Y(n_900)
);

BUFx8_ASAP7_75t_L g901 ( 
.A(n_586),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_714),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_681),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_799),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_520),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_714),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_803),
.B(n_14),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_668),
.B(n_16),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_791),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_846),
.B(n_17),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_846),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_791),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_643),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_714),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_714),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_668),
.B(n_17),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_853),
.Y(n_917)
);

BUFx12f_ASAP7_75t_L g918 ( 
.A(n_533),
.Y(n_918)
);

OAI22x1_ASAP7_75t_SL g919 ( 
.A1(n_540),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_704),
.B(n_20),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_782),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_609),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_609),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_561),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_782),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_782),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_555),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_504),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_508),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_503),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_782),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_619),
.Y(n_934)
);

XNOR2x2_ASAP7_75t_L g935 ( 
.A(n_603),
.B(n_21),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_605),
.B(n_21),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_704),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_563),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_534),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_534),
.Y(n_940)
);

CKINVDCx16_ASAP7_75t_R g941 ( 
.A(n_625),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_519),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_563),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_519),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_529),
.B(n_502),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_672),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_619),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_585),
.A2(n_289),
.B(n_288),
.Y(n_948)
);

OAI22x1_ASAP7_75t_R g949 ( 
.A1(n_625),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_672),
.B(n_25),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_509),
.B(n_27),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_585),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_566),
.B(n_27),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_663),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_634),
.Y(n_955)
);

BUFx8_ASAP7_75t_SL g956 ( 
.A(n_634),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_519),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_663),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_742),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_724),
.B(n_28),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_742),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_742),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_510),
.B(n_29),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_742),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_758),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_758),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_761),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_761),
.B(n_29),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_543),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_650),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_592),
.Y(n_971)
);

OA21x2_ASAP7_75t_L g972 ( 
.A1(n_606),
.A2(n_291),
.B(n_290),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_758),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_813),
.B(n_31),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_643),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_922),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_913),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_913),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_857),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_975),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_922),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_940),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_975),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_867),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_955),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_873),
.B(n_884),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_868),
.B(n_543),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_859),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_859),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_887),
.B(n_571),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_867),
.B(n_571),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_881),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_955),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_923),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_941),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_881),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_939),
.Y(n_997)
);

NAND2x1_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_527),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_956),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_956),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_894),
.B(n_678),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_858),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_891),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_918),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_857),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_866),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_869),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_939),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_862),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_969),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_969),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_858),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_875),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_929),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_929),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_936),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_931),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_860),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_868),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_871),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_950),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_931),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_870),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_901),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_870),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_871),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_950),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_872),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_873),
.B(n_813),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_880),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_860),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_882),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_885),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_865),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_960),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_873),
.B(n_575),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_873),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_884),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_865),
.A2(n_607),
.B(n_606),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_960),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_884),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_968),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_974),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_884),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_911),
.B(n_550),
.Y(n_1045)
);

BUFx10_ASAP7_75t_L g1046 ( 
.A(n_907),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_974),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_911),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_861),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_935),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_907),
.Y(n_1051)
);

AND2x6_ASAP7_75t_L g1052 ( 
.A(n_910),
.B(n_678),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_919),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_864),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_910),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_917),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_892),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_872),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_917),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_949),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_878),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_930),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_930),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_879),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_879),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_905),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_905),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_888),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_953),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_953),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_909),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_886),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_903),
.B(n_550),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_970),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_904),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_899),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_899),
.Y(n_1077)
);

BUFx8_ASAP7_75t_SL g1078 ( 
.A(n_903),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_928),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_928),
.Y(n_1080)
);

CKINVDCx6p67_ASAP7_75t_R g1081 ( 
.A(n_889),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_876),
.A2(n_713),
.B(n_617),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_909),
.Y(n_1083)
);

NOR2x1p5_ASAP7_75t_L g1084 ( 
.A(n_946),
.B(n_551),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_934),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_934),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_898),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_947),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_947),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_954),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_954),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_895),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_889),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_937),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_937),
.B(n_607),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_908),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_908),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_863),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_946),
.B(n_551),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_916),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_920),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_920),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_951),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_951),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_937),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_937),
.B(n_817),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_963),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_963),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_932),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_925),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_912),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_938),
.Y(n_1112)
);

XNOR2xp5_ASAP7_75t_L g1113 ( 
.A(n_900),
.B(n_650),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_938),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_967),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_943),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_958),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_952),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_912),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_948),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_958),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_924),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_971),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_971),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_924),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_944),
.Y(n_1126)
);

NOR2xp67_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_505),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_945),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_962),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_945),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_863),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_893),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_893),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_893),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_893),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_863),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_942),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_915),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_915),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_942),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_874),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_957),
.B(n_575),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_972),
.A2(n_552),
.B(n_535),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_957),
.B(n_636),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_933),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_933),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_957),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_933),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_959),
.B(n_636),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_933),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_959),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_961),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_961),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_961),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_964),
.B(n_729),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_964),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_964),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_972),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_965),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_874),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_965),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_965),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_966),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_966),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_973),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_1096),
.B(n_553),
.C(n_521),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1102),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1093),
.B(n_530),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_L g1169 ( 
.A(n_1006),
.B(n_530),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1085),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1025),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1120),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1101),
.B(n_532),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1056),
.B(n_532),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1062),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1063),
.B(n_1076),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1029),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_984),
.B(n_537),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_1039),
.A2(n_648),
.B(n_640),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1059),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1085),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1029),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1058),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_984),
.B(n_537),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1049),
.B(n_664),
.C(n_590),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1046),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1014),
.B(n_538),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_1120),
.B(n_572),
.C(n_557),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1108),
.B(n_538),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1061),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_1005),
.B(n_979),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1046),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1050),
.B(n_693),
.C(n_524),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1112),
.B(n_544),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1072),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1001),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1028),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1128),
.B(n_729),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1015),
.B(n_544),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1020),
.B(n_545),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1045),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1026),
.B(n_545),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1075),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1019),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1048),
.B(n_1116),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1123),
.B(n_549),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1086),
.B(n_549),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_1007),
.B(n_558),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1106),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1073),
.B(n_558),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1106),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1080),
.B(n_701),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1099),
.B(n_701),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1079),
.B(n_1077),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1110),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1088),
.B(n_814),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1089),
.B(n_814),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1009),
.B(n_1003),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1017),
.B(n_815),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1114),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1022),
.B(n_833),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1090),
.B(n_833),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1001),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1109),
.B(n_514),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1091),
.B(n_515),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_987),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1163),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1001),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_982),
.B(n_700),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1008),
.B(n_1075),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1004),
.B(n_554),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_L g1233 ( 
.A(n_1068),
.B(n_754),
.C(n_747),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1069),
.A2(n_783),
.B1(n_810),
.B2(n_781),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1118),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1070),
.A2(n_783),
.B1(n_810),
.B2(n_781),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1158),
.B(n_583),
.C(n_576),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1081),
.B(n_676),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1030),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1115),
.B(n_1125),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1051),
.B(n_525),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1055),
.B(n_694),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1040),
.B(n_526),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1016),
.B(n_560),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1087),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_997),
.B(n_556),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1130),
.B(n_1012),
.C(n_1002),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1124),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_SL g1249 ( 
.A(n_1001),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1023),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1002),
.A2(n_648),
.B(n_640),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1032),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1036),
.Y(n_1253)
);

AOI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_1066),
.A2(n_816),
.B1(n_818),
.B2(n_700),
.C(n_559),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1084),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1021),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1027),
.B(n_845),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1010),
.B(n_816),
.Y(n_1258)
);

INVxp33_ASAP7_75t_L g1259 ( 
.A(n_990),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1011),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1035),
.B(n_569),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1042),
.B(n_573),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1024),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1043),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1047),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_986),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1018),
.B(n_620),
.C(n_604),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1117),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1018),
.Y(n_1269)
);

INVxp33_ASAP7_75t_L g1270 ( 
.A(n_990),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1054),
.B(n_580),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1097),
.B(n_581),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1082),
.A2(n_630),
.B(n_627),
.Y(n_1273)
);

CKINVDCx11_ASAP7_75t_R g1274 ( 
.A(n_999),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1142),
.Y(n_1275)
);

NOR3xp33_ASAP7_75t_L g1276 ( 
.A(n_1067),
.B(n_802),
.C(n_776),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1037),
.B(n_591),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1038),
.B(n_597),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1052),
.B(n_1041),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1044),
.B(n_615),
.Y(n_1280)
);

BUFx2_ASAP7_75t_R g1281 ( 
.A(n_988),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1036),
.B(n_991),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1031),
.B(n_649),
.C(n_639),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1100),
.B(n_616),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_SL g1285 ( 
.A(n_1052),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1105),
.B(n_621),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1142),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1095),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1092),
.A2(n_823),
.B1(n_824),
.B2(n_819),
.C(n_818),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1034),
.B(n_626),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1034),
.B(n_629),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1121),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1095),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1127),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_991),
.B(n_722),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_989),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1057),
.B(n_632),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1071),
.B(n_633),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_977),
.B(n_819),
.Y(n_1299)
);

AO221x1_ASAP7_75t_L g1300 ( 
.A1(n_1103),
.A2(n_738),
.B1(n_797),
.B2(n_725),
.C(n_654),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1071),
.B(n_637),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1083),
.B(n_641),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1111),
.B(n_644),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1144),
.B(n_645),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1119),
.B(n_646),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1122),
.B(n_1082),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1104),
.B(n_652),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1122),
.B(n_656),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1107),
.B(n_660),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1143),
.B(n_667),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1144),
.B(n_685),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_992),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1094),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1132),
.Y(n_1314)
);

NOR2xp67_ASAP7_75t_L g1315 ( 
.A(n_978),
.B(n_823),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1139),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1126),
.Y(n_1317)
);

NAND2xp33_ASAP7_75t_L g1318 ( 
.A(n_1149),
.B(n_687),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1129),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_976),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1152),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1143),
.B(n_511),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1154),
.Y(n_1323)
);

AO221x1_ASAP7_75t_L g1324 ( 
.A1(n_1149),
.A2(n_738),
.B1(n_797),
.B2(n_725),
.C(n_654),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1065),
.A2(n_517),
.B(n_523),
.C(n_513),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1155),
.B(n_692),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1133),
.B(n_696),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1134),
.B(n_699),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1098),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1156),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1157),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1155),
.B(n_707),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1013),
.B(n_828),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_980),
.B(n_730),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_983),
.B(n_829),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1135),
.B(n_733),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_994),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1159),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_SL g1340 ( 
.A(n_996),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1138),
.B(n_756),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1078),
.B(n_759),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1145),
.B(n_760),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1146),
.B(n_763),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1113),
.B(n_766),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1148),
.B(n_662),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1150),
.B(n_671),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_995),
.B(n_831),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1162),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1164),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1000),
.B(n_774),
.Y(n_1351)
);

AND2x6_ASAP7_75t_SL g1352 ( 
.A(n_981),
.B(n_528),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1074),
.B(n_789),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1053),
.B(n_796),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_L g1355 ( 
.A(n_1098),
.B(n_805),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1098),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1033),
.B(n_808),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1137),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1060),
.B(n_811),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1140),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1147),
.B(n_674),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1151),
.B(n_812),
.Y(n_1362)
);

XOR2xp5_ASAP7_75t_L g1363 ( 
.A(n_985),
.B(n_804),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_993),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1153),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1161),
.B(n_677),
.Y(n_1366)
);

NOR3xp33_ASAP7_75t_L g1367 ( 
.A(n_1165),
.B(n_848),
.C(n_826),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1098),
.B(n_836),
.Y(n_1368)
);

AO221x1_ASAP7_75t_L g1369 ( 
.A1(n_1141),
.A2(n_804),
.B1(n_822),
.B2(n_809),
.C(n_807),
.Y(n_1369)
);

OR2x2_ASAP7_75t_SL g1370 ( 
.A(n_1131),
.B(n_807),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1131),
.B(n_682),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1141),
.B(n_842),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1136),
.B(n_688),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1141),
.B(n_851),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1141),
.B(n_852),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1136),
.B(n_824),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1096),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1096),
.B(n_705),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1096),
.B(n_715),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1096),
.B(n_718),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1025),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1096),
.B(n_732),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_998),
.B(n_817),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1096),
.B(n_855),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1096),
.B(n_856),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1096),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1096),
.B(n_740),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1096),
.B(n_743),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_998),
.B(n_841),
.Y(n_1389)
);

BUFx5_ASAP7_75t_L g1390 ( 
.A(n_1120),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1096),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1096),
.B(n_745),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1096),
.B(n_752),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1096),
.B(n_767),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1096),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1096),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1096),
.B(n_769),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1096),
.B(n_773),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1096),
.B(n_787),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1096),
.B(n_790),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_L g1401 ( 
.A(n_1001),
.B(n_651),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1096),
.B(n_801),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1096),
.B(n_825),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1096),
.B(n_830),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1096),
.B(n_837),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1096),
.B(n_827),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1096),
.B(n_838),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1096),
.B(n_854),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1167),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1377),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1386),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1391),
.B(n_829),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1395),
.Y(n_1413)
);

NOR3xp33_ASAP7_75t_SL g1414 ( 
.A(n_1296),
.B(n_831),
.C(n_507),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1205),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1396),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1172),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1228),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1204),
.B(n_531),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1258),
.B(n_809),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1237),
.A2(n_822),
.B1(n_541),
.B2(n_548),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1406),
.B(n_506),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1196),
.B(n_512),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1216),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1378),
.B(n_516),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1190),
.Y(n_1426)
);

AND2x2_ASAP7_75t_SL g1427 ( 
.A(n_1199),
.B(n_841),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_518),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1312),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1379),
.B(n_1380),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1379),
.B(n_522),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1180),
.B(n_562),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1198),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1198),
.B(n_565),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1380),
.B(n_567),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1249),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1382),
.B(n_570),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1237),
.A2(n_578),
.B1(n_579),
.B2(n_536),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1224),
.B(n_847),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1224),
.B(n_574),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1221),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1250),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1397),
.A2(n_589),
.B(n_594),
.C(n_588),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1195),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1383),
.B(n_595),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1199),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_SL g1447 ( 
.A(n_1357),
.B(n_584),
.C(n_577),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1227),
.A2(n_1202),
.B1(n_1206),
.B2(n_1230),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1245),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1383),
.B(n_600),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1400),
.A2(n_613),
.B(n_618),
.C(n_602),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1338),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_SL g1453 ( 
.A(n_1171),
.B(n_593),
.C(n_587),
.Y(n_1453)
);

OR2x4_ASAP7_75t_L g1454 ( 
.A(n_1345),
.B(n_622),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1210),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1212),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1189),
.B(n_596),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1274),
.Y(n_1458)
);

BUFx4f_ASAP7_75t_L g1459 ( 
.A(n_1295),
.Y(n_1459)
);

NOR2x2_ASAP7_75t_L g1460 ( 
.A(n_1295),
.B(n_1363),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1383),
.B(n_631),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1312),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1229),
.B(n_598),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1381),
.B(n_599),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1229),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1229),
.B(n_608),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1177),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1172),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1387),
.B(n_610),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1402),
.A2(n_658),
.B(n_659),
.C(n_647),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1235),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1333),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1387),
.A2(n_675),
.B1(n_690),
.B2(n_661),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1260),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1231),
.A2(n_612),
.B1(n_614),
.B2(n_611),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1325),
.A2(n_697),
.B(n_709),
.C(n_691),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1197),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1268),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1352),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1191),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1388),
.B(n_623),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1388),
.B(n_628),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1240),
.B(n_635),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1392),
.B(n_642),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1175),
.B(n_655),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1183),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1186),
.B(n_657),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1234),
.B(n_665),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1182),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1256),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1264),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1239),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1265),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1376),
.Y(n_1494)
);

AND2x6_ASAP7_75t_SL g1495 ( 
.A(n_1295),
.B(n_710),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1191),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1252),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1392),
.B(n_666),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1192),
.B(n_669),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1292),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1248),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1393),
.B(n_679),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1364),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1246),
.B(n_680),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1306),
.A2(n_1310),
.B(n_1322),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1249),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1317),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1322),
.A2(n_720),
.B(n_698),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1215),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1188),
.A2(n_720),
.B(n_698),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1394),
.B(n_684),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1348),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1336),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1390),
.B(n_686),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1394),
.B(n_689),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1319),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1389),
.B(n_711),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1336),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1398),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1269),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1263),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1285),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1253),
.B(n_847),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1389),
.B(n_716),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1389),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1255),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1398),
.B(n_695),
.Y(n_1527)
);

INVx5_ASAP7_75t_L g1528 ( 
.A(n_1191),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1399),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1390),
.B(n_702),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1340),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1320),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1399),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1335),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1285),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1390),
.B(n_706),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1403),
.B(n_708),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1314),
.B(n_719),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1236),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1403),
.B(n_712),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1340),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1170),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1316),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1323),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1408),
.B(n_717),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1384),
.A2(n_723),
.B1(n_727),
.B2(n_721),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1385),
.A2(n_731),
.B1(n_744),
.B2(n_739),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1288),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1293),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1407),
.B(n_748),
.Y(n_1550)
);

AND2x6_ASAP7_75t_L g1551 ( 
.A(n_1266),
.B(n_728),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1405),
.B(n_753),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1404),
.B(n_757),
.Y(n_1553)
);

OR2x6_ASAP7_75t_SL g1554 ( 
.A(n_1281),
.B(n_762),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1287),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1361),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1275),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1251),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1185),
.A2(n_772),
.B1(n_777),
.B2(n_765),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1166),
.B(n_779),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1181),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1254),
.A2(n_734),
.B1(n_735),
.B2(n_726),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1276),
.A2(n_741),
.B(n_746),
.C(n_736),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1356),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1194),
.B(n_785),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1289),
.A2(n_793),
.B1(n_795),
.B2(n_786),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1330),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1211),
.B(n_849),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1370),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1219),
.B(n_751),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1214),
.B(n_850),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1361),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1282),
.B(n_755),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1331),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1207),
.B(n_768),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1339),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1201),
.B(n_770),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1213),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1193),
.A2(n_775),
.B(n_780),
.C(n_771),
.Y(n_1579)
);

NOR2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1300),
.B(n_1324),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1366),
.Y(n_1581)
);

AOI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1233),
.A2(n_792),
.B(n_794),
.C(n_788),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1371),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1203),
.B(n_800),
.Y(n_1584)
);

NAND2x2_ASAP7_75t_L g1585 ( 
.A(n_1369),
.B(n_33),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1371),
.Y(n_1586)
);

AND3x1_ASAP7_75t_L g1587 ( 
.A(n_1359),
.B(n_1353),
.C(n_1354),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1367),
.A2(n_820),
.B1(n_821),
.B2(n_806),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1188),
.A2(n_784),
.B(n_764),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1313),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1373),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1168),
.B(n_1173),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1299),
.B(n_832),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1349),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_L g1595 ( 
.A(n_1342),
.B(n_35),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1242),
.A2(n_839),
.B1(n_844),
.B2(n_834),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1307),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1309),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1272),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1178),
.B(n_843),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1373),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1267),
.A2(n_1283),
.B1(n_1247),
.B2(n_1346),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_SL g1603 ( 
.A(n_1321),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1184),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_SL g1605 ( 
.A(n_1259),
.B(n_1270),
.C(n_1284),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1257),
.B(n_1273),
.Y(n_1606)
);

AND2x6_ASAP7_75t_SL g1607 ( 
.A(n_1351),
.B(n_35),
.Y(n_1607)
);

AND2x6_ASAP7_75t_SL g1608 ( 
.A(n_1271),
.B(n_36),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1244),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_R g1610 ( 
.A(n_1318),
.B(n_36),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1179),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1283),
.A2(n_840),
.B1(n_778),
.B2(n_973),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1176),
.B(n_1232),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1179),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1273),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1262),
.A2(n_840),
.B1(n_778),
.B2(n_877),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1390),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1315),
.Y(n_1618)
);

AND2x6_ASAP7_75t_SL g1619 ( 
.A(n_1238),
.B(n_38),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1169),
.B(n_41),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1401),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1174),
.B(n_42),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1261),
.B(n_45),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1294),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1187),
.A2(n_883),
.B1(n_890),
.B2(n_877),
.Y(n_1625)
);

INVx5_ASAP7_75t_L g1626 ( 
.A(n_1329),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1200),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1225),
.B(n_51),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1220),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1350),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1209),
.B(n_883),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1277),
.B(n_52),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1243),
.Y(n_1633)
);

AND3x1_ASAP7_75t_L g1634 ( 
.A(n_1222),
.B(n_53),
.C(n_54),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1346),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1208),
.B(n_53),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1241),
.A2(n_897),
.B1(n_902),
.B2(n_896),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1217),
.B(n_1218),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1347),
.A2(n_897),
.B1(n_902),
.B2(n_896),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1290),
.A2(n_902),
.B(n_897),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1223),
.A2(n_1304),
.B1(n_1326),
.B2(n_1311),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1334),
.B(n_56),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1347),
.B(n_58),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1329),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1226),
.B(n_58),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1343),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1291),
.B(n_59),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1329),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1301),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1302),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_SL g1652 ( 
.A(n_1358),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1332),
.A2(n_914),
.B1(n_921),
.B2(n_906),
.Y(n_1653)
);

NOR2x2_ASAP7_75t_L g1654 ( 
.A(n_1278),
.B(n_60),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1303),
.A2(n_914),
.B1(n_921),
.B2(n_906),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1305),
.B(n_61),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1308),
.B(n_61),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1280),
.B(n_62),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1327),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1279),
.B(n_62),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1368),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1344),
.A2(n_1362),
.B1(n_1374),
.B2(n_1372),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1375),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1329),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1328),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1286),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1337),
.Y(n_1667)
);

NOR2x2_ASAP7_75t_L g1668 ( 
.A(n_1360),
.B(n_63),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1341),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1355),
.A2(n_1365),
.B1(n_926),
.B2(n_927),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1356),
.B(n_921),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1167),
.A2(n_927),
.B1(n_926),
.B2(n_70),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1338),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1167),
.B(n_68),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1205),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1564),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1452),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1539),
.B(n_68),
.Y(n_1678)
);

INVx6_ASAP7_75t_L g1679 ( 
.A(n_1531),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1443),
.A2(n_73),
.B(n_69),
.C(n_72),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1505),
.A2(n_927),
.B(n_926),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1626),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1582),
.B(n_72),
.C(n_74),
.Y(n_1683)
);

OA22x2_ASAP7_75t_L g1684 ( 
.A1(n_1509),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1430),
.B(n_1519),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1626),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1648),
.A2(n_1533),
.B(n_1529),
.Y(n_1687)
);

OAI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1425),
.A2(n_75),
.B(n_76),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1415),
.B(n_1509),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1626),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1429),
.B(n_77),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1635),
.B(n_77),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1451),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1675),
.Y(n_1694)
);

AOI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1432),
.A2(n_79),
.B(n_80),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1410),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1411),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1413),
.Y(n_1698)
);

BUFx4f_ASAP7_75t_L g1699 ( 
.A(n_1479),
.Y(n_1699)
);

AO22x1_ASAP7_75t_L g1700 ( 
.A1(n_1531),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1454),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1556),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1462),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1420),
.B(n_87),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1409),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1416),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1472),
.B(n_1488),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1611),
.A2(n_309),
.B(n_308),
.Y(n_1708)
);

OR2x6_ASAP7_75t_L g1709 ( 
.A(n_1436),
.B(n_88),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1474),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1651),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1425),
.B(n_91),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1512),
.B(n_92),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1428),
.B(n_93),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1614),
.A2(n_318),
.B(n_316),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1446),
.B(n_94),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1492),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_94),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1458),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1428),
.B(n_95),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1543),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1431),
.B(n_95),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1673),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1418),
.B(n_96),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1572),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1465),
.Y(n_1727)
);

AOI22x1_ASAP7_75t_L g1728 ( 
.A1(n_1640),
.A2(n_324),
.B1(n_325),
.B2(n_322),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1435),
.B(n_1437),
.Y(n_1729)
);

NOR2x1p5_ASAP7_75t_SL g1730 ( 
.A(n_1558),
.B(n_1583),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1628),
.A2(n_103),
.B(n_100),
.C(n_101),
.Y(n_1731)
);

NOR3xp33_ASAP7_75t_L g1732 ( 
.A(n_1453),
.B(n_101),
.C(n_103),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1541),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1534),
.B(n_104),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1532),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1448),
.B(n_1599),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1581),
.A2(n_108),
.B(n_105),
.C(n_106),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1426),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_R g1739 ( 
.A(n_1459),
.B(n_109),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1586),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1442),
.B(n_113),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1497),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1508),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1470),
.A2(n_122),
.B(n_119),
.C(n_120),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1674),
.A2(n_124),
.B1(n_119),
.B2(n_123),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1610),
.B(n_127),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1481),
.B(n_128),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1504),
.B(n_128),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1419),
.B(n_129),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1569),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1563),
.A2(n_135),
.B(n_131),
.C(n_133),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1459),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1521),
.B(n_133),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1444),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1482),
.A2(n_334),
.B(n_332),
.Y(n_1755)
);

O2A1O1Ixp5_ASAP7_75t_SL g1756 ( 
.A1(n_1655),
.A2(n_337),
.B(n_339),
.C(n_336),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1591),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1449),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1609),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1507),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1484),
.B(n_139),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1484),
.B(n_1498),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1503),
.B(n_141),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1498),
.B(n_142),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_SL g1765 ( 
.A1(n_1647),
.A2(n_346),
.B(n_347),
.C(n_343),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1601),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1602),
.A2(n_349),
.B(n_348),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_SL g1768 ( 
.A(n_1629),
.B(n_143),
.C(n_144),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1478),
.B(n_1500),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1516),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1419),
.B(n_145),
.Y(n_1771)
);

OAI22x1_ASAP7_75t_L g1772 ( 
.A1(n_1580),
.A2(n_1668),
.B1(n_1632),
.B2(n_1620),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1585),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1480),
.B(n_146),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1579),
.A2(n_151),
.B(n_147),
.C(n_149),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1454),
.B(n_149),
.Y(n_1776)
);

OAI21xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1643),
.A2(n_151),
.B(n_152),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1502),
.B(n_1511),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1526),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1511),
.A2(n_155),
.B1(n_152),
.B2(n_154),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1476),
.A2(n_1473),
.B(n_1643),
.C(n_1537),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1418),
.B(n_156),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1578),
.B(n_159),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1465),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1548),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_R g1786 ( 
.A(n_1495),
.B(n_161),
.Y(n_1786)
);

OAI22x1_ASAP7_75t_L g1787 ( 
.A1(n_1632),
.A2(n_1620),
.B1(n_1554),
.B2(n_1460),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1570),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_1570),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1570),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1515),
.B(n_163),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1602),
.A2(n_366),
.B(n_365),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1667),
.B(n_163),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1537),
.B(n_164),
.Y(n_1794)
);

OAI22x1_ASAP7_75t_L g1795 ( 
.A1(n_1523),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1652),
.B(n_165),
.Y(n_1796)
);

NOR3xp33_ASAP7_75t_L g1797 ( 
.A(n_1605),
.B(n_167),
.C(n_169),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1540),
.B(n_169),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1540),
.B(n_170),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1555),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1496),
.B(n_171),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1549),
.B(n_172),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1490),
.Y(n_1803)
);

OAI21xp33_ASAP7_75t_L g1804 ( 
.A1(n_1438),
.A2(n_1596),
.B(n_1421),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_SL g1805 ( 
.A(n_1496),
.B(n_172),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1491),
.B(n_173),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1493),
.B(n_174),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1582),
.B(n_174),
.C(n_175),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1469),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_1809)
);

OR2x6_ASAP7_75t_L g1810 ( 
.A(n_1525),
.B(n_176),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1633),
.A2(n_373),
.B(n_372),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1445),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1501),
.Y(n_1813)
);

NOR2xp67_ASAP7_75t_L g1814 ( 
.A(n_1496),
.B(n_380),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1464),
.B(n_180),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_SL g1816 ( 
.A(n_1613),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1551),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_1817)
);

OA22x2_ASAP7_75t_L g1818 ( 
.A1(n_1613),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1644),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1527),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1485),
.B(n_191),
.C(n_192),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1494),
.B(n_191),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1551),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1562),
.B(n_1669),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_R g1825 ( 
.A(n_1506),
.B(n_192),
.Y(n_1825)
);

AO32x2_ASAP7_75t_L g1826 ( 
.A1(n_1655),
.A2(n_195),
.A3(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1575),
.B(n_196),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1424),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1545),
.A2(n_197),
.B(n_200),
.C(n_202),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1441),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1604),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1659),
.B(n_205),
.Y(n_1832)
);

OR2x6_ASAP7_75t_L g1833 ( 
.A(n_1613),
.B(n_206),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1523),
.B(n_209),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1551),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_SL g1836 ( 
.A(n_1447),
.B(n_1666),
.C(n_1414),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1551),
.A2(n_1634),
.B1(n_1538),
.B2(n_1587),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1665),
.B(n_211),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1514),
.A2(n_388),
.B(n_384),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1608),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1657),
.A2(n_211),
.B(n_212),
.C(n_213),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1575),
.B(n_212),
.Y(n_1842)
);

OR2x6_ASAP7_75t_SL g1843 ( 
.A(n_1654),
.B(n_213),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1412),
.B(n_214),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1577),
.B(n_214),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1584),
.B(n_215),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1550),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1592),
.B(n_220),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1487),
.B(n_221),
.C(n_222),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1607),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1455),
.B(n_223),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1564),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1623),
.A2(n_1589),
.B(n_1510),
.C(n_1656),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1536),
.A2(n_416),
.B(n_497),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1634),
.A2(n_1538),
.B1(n_1587),
.B2(n_1622),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1471),
.Y(n_1856)
);

BUFx2_ASAP7_75t_SL g1857 ( 
.A(n_1652),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1552),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1456),
.B(n_225),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1619),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1650),
.B(n_226),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1552),
.A2(n_226),
.B(n_228),
.C(n_229),
.Y(n_1862)
);

OAI21xp33_ASAP7_75t_L g1863 ( 
.A1(n_1553),
.A2(n_228),
.B(n_229),
.Y(n_1863)
);

O2A1O1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1553),
.A2(n_232),
.B(n_234),
.C(n_237),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1467),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1450),
.Y(n_1866)
);

OAI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1623),
.A2(n_1589),
.B(n_1510),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1461),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1600),
.A2(n_419),
.B(n_495),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1565),
.A2(n_413),
.B(n_494),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1461),
.B(n_234),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1664),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1520),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1489),
.B(n_237),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1565),
.A2(n_1568),
.B(n_1422),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1621),
.A2(n_1568),
.B1(n_1528),
.B2(n_1457),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1636),
.A2(n_239),
.B(n_241),
.C(n_242),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1638),
.B(n_241),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1517),
.B(n_242),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1645),
.A2(n_244),
.B(n_245),
.C(n_246),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1528),
.B(n_246),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1517),
.B(n_247),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1588),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.C(n_250),
.Y(n_1883)
);

OR2x6_ASAP7_75t_L g1884 ( 
.A(n_1646),
.B(n_249),
.Y(n_1884)
);

AO32x2_ASAP7_75t_L g1885 ( 
.A1(n_1544),
.A2(n_251),
.A3(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1576),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1524),
.B(n_258),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1621),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_1888)
);

BUFx12f_ASAP7_75t_L g1889 ( 
.A(n_1593),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1524),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1528),
.B(n_263),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1477),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1630),
.B(n_264),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1594),
.Y(n_1894)
);

AND2x4_ASAP7_75t_SL g1895 ( 
.A(n_1644),
.B(n_265),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1571),
.B(n_265),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1560),
.B(n_266),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1465),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1660),
.A2(n_431),
.B(n_484),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1593),
.Y(n_1900)
);

O2A1O1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1618),
.A2(n_270),
.B(n_272),
.C(n_273),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1660),
.A2(n_270),
.B1(n_274),
.B2(n_275),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1557),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_SL g1904 ( 
.A(n_1499),
.B(n_276),
.C(n_277),
.Y(n_1904)
);

A2O1A1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1658),
.A2(n_277),
.B(n_279),
.C(n_280),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1506),
.B(n_279),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1641),
.A2(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1483),
.B(n_284),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1624),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1433),
.Y(n_1910)
);

AO21x1_ASAP7_75t_L g1911 ( 
.A1(n_1617),
.A2(n_391),
.B(n_396),
.Y(n_1911)
);

CKINVDCx6p67_ASAP7_75t_R g1912 ( 
.A(n_1603),
.Y(n_1912)
);

BUFx12f_ASAP7_75t_L g1913 ( 
.A(n_1567),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1417),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1468),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1590),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_R g1917 ( 
.A(n_1522),
.B(n_406),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1627),
.A2(n_411),
.B(n_412),
.C(n_423),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1475),
.B(n_428),
.Y(n_1919)
);

AND2x6_ASAP7_75t_L g1920 ( 
.A(n_1522),
.B(n_435),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1603),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1642),
.B(n_446),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1574),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1535),
.B(n_500),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1649),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1535),
.B(n_482),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1566),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1439),
.A2(n_464),
.B1(n_465),
.B2(n_466),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1546),
.B(n_468),
.Y(n_1929)
);

O2A1O1Ixp33_ASAP7_75t_SL g1930 ( 
.A1(n_1671),
.A2(n_473),
.B(n_474),
.C(n_475),
.Y(n_1930)
);

BUFx12f_ASAP7_75t_L g1931 ( 
.A(n_1631),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1547),
.B(n_479),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1661),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1513),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1595),
.A2(n_1559),
.B1(n_1663),
.B2(n_1573),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1486),
.B(n_1662),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1423),
.A2(n_1434),
.B(n_1440),
.C(n_1463),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1542),
.A2(n_1561),
.B1(n_1672),
.B2(n_1466),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_SL g1939 ( 
.A(n_1616),
.B(n_1653),
.C(n_1639),
.Y(n_1939)
);

INVx4_ASAP7_75t_L g1940 ( 
.A(n_1433),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1631),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_SL g1942 ( 
.A(n_1631),
.B(n_1649),
.C(n_1637),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1518),
.A2(n_1612),
.B(n_1670),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1625),
.A2(n_1430),
.B1(n_1065),
.B2(n_1427),
.Y(n_1944)
);

O2A1O1Ixp5_ASAP7_75t_L g1945 ( 
.A1(n_1606),
.A2(n_1615),
.B(n_1602),
.C(n_1530),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1539),
.B(n_1103),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_R g1947 ( 
.A(n_1452),
.B(n_1673),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1409),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1564),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1505),
.A2(n_1430),
.B(n_1306),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1539),
.A2(n_1065),
.B1(n_1066),
.B2(n_1064),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1430),
.B(n_1519),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1430),
.B(n_1519),
.Y(n_1953)
);

BUFx2_ASAP7_75t_SL g1954 ( 
.A(n_1788),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1867),
.A2(n_1687),
.B(n_1945),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1719),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1867),
.A2(n_1853),
.B(n_1778),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1685),
.B(n_1952),
.Y(n_1958)
);

NAND2x1p5_ASAP7_75t_L g1959 ( 
.A(n_1682),
.B(n_1686),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_SL g1960 ( 
.A1(n_1837),
.A2(n_1792),
.B(n_1767),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1947),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1736),
.B(n_1724),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1676),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1943),
.A2(n_1715),
.B(n_1756),
.Y(n_1964)
);

AO21x2_ASAP7_75t_L g1965 ( 
.A1(n_1688),
.A2(n_1863),
.B(n_1875),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1789),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1707),
.B(n_1689),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_SL g1968 ( 
.A1(n_1837),
.A2(n_1953),
.B(n_1745),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1729),
.A2(n_1781),
.B(n_1762),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1703),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1876),
.A2(n_1714),
.B(n_1712),
.Y(n_1971)
);

OAI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1897),
.A2(n_1722),
.B(n_1720),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_L g1973 ( 
.A1(n_1728),
.A2(n_1899),
.B(n_1869),
.Y(n_1973)
);

BUFx2_ASAP7_75t_R g1974 ( 
.A(n_1677),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1735),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1886),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1793),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1721),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1779),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1785),
.B(n_1824),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_SL g1981 ( 
.A(n_1718),
.B(n_1774),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1699),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1686),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1718),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1717),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1690),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1705),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1946),
.B(n_1951),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1718),
.B(n_1834),
.Y(n_1989)
);

BUFx4f_ASAP7_75t_SL g1990 ( 
.A(n_1912),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1738),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1804),
.B(n_1706),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1694),
.B(n_1710),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1727),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1866),
.B(n_1832),
.Y(n_1995)
);

INVxp67_ASAP7_75t_SL g1996 ( 
.A(n_1793),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1699),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1742),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1758),
.Y(n_1999)
);

OAI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1747),
.A2(n_1764),
.B(n_1761),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1834),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1760),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1894),
.Y(n_2003)
);

AO21x2_ASAP7_75t_L g2004 ( 
.A1(n_1688),
.A2(n_1863),
.B(n_1911),
.Y(n_2004)
);

BUFx2_ASAP7_75t_SL g2005 ( 
.A(n_1816),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1769),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_SL g2007 ( 
.A1(n_1745),
.A2(n_1780),
.B(n_1858),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1794),
.A2(n_1799),
.B(n_1798),
.Y(n_2008)
);

OAI21x1_ASAP7_75t_SL g2009 ( 
.A1(n_1780),
.A2(n_1858),
.B(n_1784),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1679),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1769),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1834),
.Y(n_2012)
);

INVx6_ASAP7_75t_L g2013 ( 
.A(n_1769),
.Y(n_2013)
);

BUFx2_ASAP7_75t_SL g2014 ( 
.A(n_1816),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_1913),
.Y(n_2015)
);

BUFx12f_ASAP7_75t_L g2016 ( 
.A(n_1679),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1727),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1770),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1893),
.Y(n_2019)
);

AO21x2_ASAP7_75t_L g2020 ( 
.A1(n_1765),
.A2(n_1814),
.B(n_1855),
.Y(n_2020)
);

AOI22x1_ASAP7_75t_L g2021 ( 
.A1(n_1772),
.A2(n_1839),
.B1(n_1854),
.B2(n_1811),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1827),
.A2(n_1842),
.B(n_1692),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1777),
.A2(n_1804),
.B(n_1802),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1790),
.B(n_1813),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1696),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1872),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1697),
.Y(n_2027)
);

OAI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1777),
.A2(n_1846),
.B(n_1845),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1723),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1784),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1739),
.Y(n_2031)
);

CKINVDCx11_ASAP7_75t_R g2032 ( 
.A(n_1843),
.Y(n_2032)
);

AOI22x1_ASAP7_75t_L g2033 ( 
.A1(n_1787),
.A2(n_1795),
.B1(n_1791),
.B2(n_1817),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1931),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1754),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1822),
.A2(n_1807),
.B(n_1806),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_1893),
.Y(n_2037)
);

AO21x2_ASAP7_75t_L g2038 ( 
.A1(n_1814),
.A2(n_1855),
.B(n_1801),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1895),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_1868),
.Y(n_2040)
);

INVxp67_ASAP7_75t_SL g2041 ( 
.A(n_1852),
.Y(n_2041)
);

BUFx10_ASAP7_75t_L g2042 ( 
.A(n_1763),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1890),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1800),
.B(n_1903),
.Y(n_2044)
);

CKINVDCx20_ASAP7_75t_R g2045 ( 
.A(n_1733),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_1852),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_1797),
.B(n_1732),
.C(n_1768),
.Y(n_2047)
);

BUFx12f_ASAP7_75t_L g2048 ( 
.A(n_1921),
.Y(n_2048)
);

OAI21xp33_ASAP7_75t_L g2049 ( 
.A1(n_1678),
.A2(n_1704),
.B(n_1848),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1803),
.B(n_1948),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1819),
.B(n_1730),
.Y(n_2051)
);

INVx3_ASAP7_75t_SL g2052 ( 
.A(n_1763),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1805),
.B(n_1823),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1910),
.A2(n_1941),
.B(n_1928),
.Y(n_2054)
);

NAND2x1p5_ASAP7_75t_L g2055 ( 
.A(n_1940),
.B(n_1835),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1698),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1889),
.Y(n_2057)
);

AO21x2_ASAP7_75t_L g2058 ( 
.A1(n_1881),
.A2(n_1891),
.B(n_1939),
.Y(n_2058)
);

AO21x2_ASAP7_75t_L g2059 ( 
.A1(n_1918),
.A2(n_1936),
.B(n_1743),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1763),
.Y(n_2060)
);

OAI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1896),
.A2(n_1844),
.B(n_1851),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1819),
.A2(n_1937),
.B(n_1938),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1713),
.B(n_1871),
.Y(n_2063)
);

INVx6_ASAP7_75t_L g2064 ( 
.A(n_1940),
.Y(n_2064)
);

BUFx2_ASAP7_75t_SL g2065 ( 
.A(n_1920),
.Y(n_2065)
);

CKINVDCx14_ASAP7_75t_R g2066 ( 
.A(n_1786),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1753),
.B(n_1833),
.Y(n_2067)
);

BUFx3_ASAP7_75t_L g2068 ( 
.A(n_1753),
.Y(n_2068)
);

INVx5_ASAP7_75t_L g2069 ( 
.A(n_1914),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1753),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_1938),
.A2(n_1922),
.B(n_1873),
.Y(n_2071)
);

INVx3_ASAP7_75t_SL g2072 ( 
.A(n_1752),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1810),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1865),
.B(n_1828),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1925),
.Y(n_2075)
);

CKINVDCx16_ASAP7_75t_R g2076 ( 
.A(n_1709),
.Y(n_2076)
);

INVx8_ASAP7_75t_L g2077 ( 
.A(n_1709),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1830),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1833),
.B(n_1909),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1914),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1914),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1810),
.Y(n_2082)
);

INVx5_ASAP7_75t_L g2083 ( 
.A(n_1915),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1856),
.Y(n_2084)
);

INVx5_ASAP7_75t_L g2085 ( 
.A(n_1915),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_1709),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1892),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1810),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_1852),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1833),
.B(n_1933),
.Y(n_2090)
);

INVx3_ASAP7_75t_SL g2091 ( 
.A(n_1884),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1859),
.A2(n_1874),
.B(n_1878),
.Y(n_2092)
);

CKINVDCx16_ASAP7_75t_R g2093 ( 
.A(n_1825),
.Y(n_2093)
);

BUFx2_ASAP7_75t_SL g2094 ( 
.A(n_1920),
.Y(n_2094)
);

CKINVDCx20_ASAP7_75t_R g2095 ( 
.A(n_1857),
.Y(n_2095)
);

AO21x2_ASAP7_75t_L g2096 ( 
.A1(n_1841),
.A2(n_1737),
.B(n_1942),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1701),
.A2(n_1683),
.B1(n_1808),
.B2(n_1836),
.Y(n_2097)
);

AO21x2_ASAP7_75t_L g2098 ( 
.A1(n_1711),
.A2(n_1731),
.B(n_1759),
.Y(n_2098)
);

BUFx2_ASAP7_75t_R g2099 ( 
.A(n_1840),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_1906),
.Y(n_2100)
);

INVx8_ASAP7_75t_L g2101 ( 
.A(n_1884),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1861),
.B(n_1783),
.Y(n_2102)
);

OAI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_1932),
.A2(n_1680),
.B(n_1744),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_1906),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1884),
.Y(n_2105)
);

OA21x2_ASAP7_75t_L g2106 ( 
.A1(n_1683),
.A2(n_1808),
.B(n_1927),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1693),
.A2(n_1944),
.B(n_1929),
.Y(n_2107)
);

BUFx12f_ASAP7_75t_L g2108 ( 
.A(n_1850),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1916),
.Y(n_2109)
);

CKINVDCx16_ASAP7_75t_R g2110 ( 
.A(n_1796),
.Y(n_2110)
);

NAND2x1p5_ASAP7_75t_L g2111 ( 
.A(n_1949),
.B(n_1934),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1944),
.B(n_1935),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1684),
.Y(n_2113)
);

OAI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1919),
.A2(n_1877),
.B(n_1880),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1924),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1701),
.A2(n_1776),
.B1(n_1748),
.B2(n_1818),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1838),
.B(n_1815),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1725),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1900),
.B(n_1924),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1782),
.Y(n_2120)
);

INVx4_ASAP7_75t_L g2121 ( 
.A(n_1920),
.Y(n_2121)
);

AO21x2_ASAP7_75t_L g2122 ( 
.A1(n_1716),
.A2(n_1905),
.B(n_1864),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_1879),
.B(n_1887),
.Y(n_2123)
);

NAND3xp33_ASAP7_75t_L g2124 ( 
.A(n_1773),
.B(n_1829),
.C(n_1862),
.Y(n_2124)
);

BUFx2_ASAP7_75t_SL g2125 ( 
.A(n_1920),
.Y(n_2125)
);

HB1xp67_ASAP7_75t_L g2126 ( 
.A(n_1898),
.Y(n_2126)
);

BUFx8_ASAP7_75t_L g2127 ( 
.A(n_1885),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_1902),
.A2(n_1847),
.B(n_1901),
.Y(n_2128)
);

INVx5_ASAP7_75t_L g2129 ( 
.A(n_1949),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_1935),
.A2(n_1809),
.B(n_1820),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1860),
.Y(n_2131)
);

BUFx2_ASAP7_75t_R g2132 ( 
.A(n_1746),
.Y(n_2132)
);

INVx8_ASAP7_75t_L g2133 ( 
.A(n_1926),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1923),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1751),
.A2(n_1775),
.B(n_1882),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1849),
.Y(n_2136)
);

INVx5_ASAP7_75t_L g2137 ( 
.A(n_1926),
.Y(n_2137)
);

NAND2x1p5_ASAP7_75t_L g2138 ( 
.A(n_1749),
.B(n_1771),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1917),
.Y(n_2139)
);

AOI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_1930),
.A2(n_1695),
.B(n_1907),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1734),
.Y(n_2141)
);

NAND2x1p5_ASAP7_75t_L g2142 ( 
.A(n_1691),
.B(n_1741),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_1700),
.Y(n_2143)
);

INVx4_ASAP7_75t_L g2144 ( 
.A(n_1904),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_1740),
.A2(n_1766),
.B(n_1757),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1702),
.A2(n_1726),
.B(n_1888),
.Y(n_2146)
);

AO21x2_ASAP7_75t_L g2147 ( 
.A1(n_1831),
.A2(n_1821),
.B(n_1908),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1883),
.B(n_1812),
.Y(n_2148)
);

OAI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1750),
.A2(n_1885),
.B(n_1826),
.Y(n_2149)
);

INVx6_ASAP7_75t_SL g2150 ( 
.A(n_1826),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_1679),
.Y(n_2151)
);

BUFx12f_ASAP7_75t_L g2152 ( 
.A(n_1679),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_1788),
.Y(n_2153)
);

HB1xp67_ASAP7_75t_L g2154 ( 
.A(n_1718),
.Y(n_2154)
);

INVx4_ASAP7_75t_L g2155 ( 
.A(n_1679),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1703),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1946),
.B(n_1539),
.Y(n_2157)
);

NAND2x1_ASAP7_75t_L g2158 ( 
.A(n_1682),
.B(n_1686),
.Y(n_2158)
);

AO21x2_ASAP7_75t_L g2159 ( 
.A1(n_1767),
.A2(n_1792),
.B(n_1606),
.Y(n_2159)
);

INVx3_ASAP7_75t_SL g2160 ( 
.A(n_1679),
.Y(n_2160)
);

AOI22x1_ASAP7_75t_L g2161 ( 
.A1(n_1875),
.A2(n_1870),
.B1(n_1580),
.B2(n_1755),
.Y(n_2161)
);

OA21x2_ASAP7_75t_L g2162 ( 
.A1(n_1945),
.A2(n_1615),
.B(n_1767),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1685),
.B(n_1952),
.Y(n_2163)
);

INVx4_ASAP7_75t_L g2164 ( 
.A(n_1679),
.Y(n_2164)
);

NAND2x1p5_ASAP7_75t_L g2165 ( 
.A(n_1682),
.B(n_1686),
.Y(n_2165)
);

OR2x6_ASAP7_75t_L g2166 ( 
.A(n_1718),
.B(n_1834),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_L g2167 ( 
.A1(n_1681),
.A2(n_1950),
.B(n_1708),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1685),
.B(n_1952),
.Y(n_2168)
);

BUFx10_ASAP7_75t_L g2169 ( 
.A(n_1679),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_1703),
.Y(n_2170)
);

AOI22x1_ASAP7_75t_L g2171 ( 
.A1(n_1875),
.A2(n_1870),
.B1(n_1580),
.B2(n_1755),
.Y(n_2171)
);

BUFx2_ASAP7_75t_SL g2172 ( 
.A(n_1788),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1685),
.Y(n_2173)
);

AO21x2_ASAP7_75t_L g2174 ( 
.A1(n_1767),
.A2(n_1792),
.B(n_1606),
.Y(n_2174)
);

CKINVDCx20_ASAP7_75t_R g2175 ( 
.A(n_1719),
.Y(n_2175)
);

OR2x6_ASAP7_75t_SL g2176 ( 
.A(n_1677),
.B(n_1452),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_1681),
.A2(n_1950),
.B(n_1708),
.Y(n_2177)
);

OAI21x1_ASAP7_75t_L g2178 ( 
.A1(n_1681),
.A2(n_1950),
.B(n_1708),
.Y(n_2178)
);

CKINVDCx8_ASAP7_75t_R g2179 ( 
.A(n_1857),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1685),
.B(n_1952),
.Y(n_2180)
);

AO21x2_ASAP7_75t_L g2181 ( 
.A1(n_1767),
.A2(n_1792),
.B(n_1606),
.Y(n_2181)
);

OAI21x1_ASAP7_75t_L g2182 ( 
.A1(n_1681),
.A2(n_1950),
.B(n_1708),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1685),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_1685),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1867),
.A2(n_1950),
.B(n_1687),
.Y(n_2185)
);

AOI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_1950),
.A2(n_1505),
.B(n_1430),
.Y(n_2186)
);

INVxp67_ASAP7_75t_SL g2187 ( 
.A(n_1685),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1958),
.Y(n_2188)
);

OA21x2_ASAP7_75t_L g2189 ( 
.A1(n_1955),
.A2(n_2185),
.B(n_1964),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2050),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1979),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1958),
.Y(n_2192)
);

BUFx2_ASAP7_75t_L g2193 ( 
.A(n_1989),
.Y(n_2193)
);

CKINVDCx20_ASAP7_75t_R g2194 ( 
.A(n_1956),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_1989),
.A2(n_2166),
.B1(n_2187),
.B2(n_1977),
.Y(n_2195)
);

CKINVDCx11_ASAP7_75t_R g2196 ( 
.A(n_2176),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2180),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2050),
.Y(n_2198)
);

BUFx3_ASAP7_75t_L g2199 ( 
.A(n_1956),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2187),
.B(n_2163),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1967),
.B(n_1962),
.Y(n_2201)
);

OAI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_2166),
.A2(n_1981),
.B1(n_2076),
.B2(n_2133),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2157),
.A2(n_1988),
.B1(n_2166),
.B2(n_2007),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1977),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_2175),
.Y(n_2205)
);

BUFx2_ASAP7_75t_L g2206 ( 
.A(n_1975),
.Y(n_2206)
);

INVx1_ASAP7_75t_SL g2207 ( 
.A(n_2184),
.Y(n_2207)
);

CKINVDCx11_ASAP7_75t_R g2208 ( 
.A(n_2175),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2033),
.A2(n_1968),
.B1(n_2049),
.B2(n_2116),
.Y(n_2209)
);

AOI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_2116),
.A2(n_2112),
.B1(n_2047),
.B2(n_2012),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_1975),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1978),
.Y(n_2212)
);

INVx4_ASAP7_75t_L g2213 ( 
.A(n_2012),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2035),
.Y(n_2214)
);

INVx6_ASAP7_75t_L g2215 ( 
.A(n_2169),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2163),
.B(n_2168),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2186),
.A2(n_2185),
.B(n_1996),
.Y(n_2217)
);

HB1xp67_ASAP7_75t_L g2218 ( 
.A(n_2184),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_1981),
.A2(n_1996),
.B1(n_2112),
.B2(n_2168),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_2121),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_2144),
.B(n_2001),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2173),
.B(n_2183),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1991),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1999),
.Y(n_2224)
);

OAI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2133),
.A2(n_2012),
.B1(n_2052),
.B2(n_2093),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2002),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2018),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2109),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_SL g2229 ( 
.A1(n_2077),
.A2(n_2133),
.B1(n_2101),
.B2(n_2001),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1987),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2074),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_1982),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_SL g2233 ( 
.A1(n_2031),
.A2(n_2094),
.B1(n_2125),
.B2(n_2065),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_2095),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2169),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_2051),
.Y(n_2236)
);

BUFx2_ASAP7_75t_L g2237 ( 
.A(n_1966),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_2019),
.Y(n_2238)
);

BUFx12f_ASAP7_75t_SL g2239 ( 
.A(n_2060),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2078),
.Y(n_2240)
);

BUFx2_ASAP7_75t_R g2241 ( 
.A(n_1997),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2084),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2047),
.A2(n_2012),
.B1(n_2077),
.B2(n_2144),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2137),
.A2(n_2052),
.B1(n_2121),
.B2(n_1984),
.Y(n_2244)
);

OAI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_2091),
.A2(n_2077),
.B1(n_2110),
.B2(n_2137),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2087),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_2060),
.A2(n_2101),
.B1(n_2102),
.B2(n_2009),
.Y(n_2247)
);

OA21x2_ASAP7_75t_L g2248 ( 
.A1(n_1955),
.A2(n_2177),
.B(n_2167),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_SL g2249 ( 
.A1(n_2101),
.A2(n_2154),
.B1(n_2067),
.B2(n_2105),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_1959),
.Y(n_2250)
);

OA21x2_ASAP7_75t_L g2251 ( 
.A1(n_2178),
.A2(n_2182),
.B(n_1971),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2025),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2027),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2056),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_1990),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1969),
.B(n_1980),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1969),
.B(n_1980),
.Y(n_2257)
);

INVx6_ASAP7_75t_L g2258 ( 
.A(n_2016),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_1990),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2137),
.A2(n_2091),
.B1(n_2097),
.B2(n_2115),
.Y(n_2260)
);

HB1xp67_ASAP7_75t_L g2261 ( 
.A(n_2051),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2107),
.A2(n_2147),
.B1(n_2097),
.B2(n_2113),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1992),
.B(n_1957),
.Y(n_2263)
);

OAI22xp33_ASAP7_75t_SL g2264 ( 
.A1(n_2082),
.A2(n_2073),
.B1(n_2143),
.B2(n_2053),
.Y(n_2264)
);

BUFx3_ASAP7_75t_L g2265 ( 
.A(n_2095),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2136),
.A2(n_2031),
.B1(n_2148),
.B2(n_2107),
.Y(n_2266)
);

AOI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2147),
.A2(n_2139),
.B1(n_2032),
.B2(n_2136),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_2152),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2069),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2063),
.B(n_1995),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2070),
.A2(n_2082),
.B1(n_2068),
.B2(n_2127),
.Y(n_2271)
);

OAI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2139),
.A2(n_2053),
.B1(n_2143),
.B2(n_2086),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_1985),
.B(n_1998),
.Y(n_2273)
);

BUFx6f_ASAP7_75t_L g2274 ( 
.A(n_2069),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2090),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2090),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2024),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_2069),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2126),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_2069),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_1970),
.Y(n_2281)
);

OAI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2023),
.A2(n_2186),
.B(n_1957),
.Y(n_2282)
);

BUFx8_ASAP7_75t_L g2283 ( 
.A(n_2015),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2024),
.Y(n_2284)
);

INVx6_ASAP7_75t_L g2285 ( 
.A(n_2155),
.Y(n_2285)
);

OA21x2_ASAP7_75t_L g2286 ( 
.A1(n_2023),
.A2(n_1960),
.B(n_1973),
.Y(n_2286)
);

BUFx2_ASAP7_75t_SL g2287 ( 
.A(n_2179),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2044),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2079),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1985),
.B(n_1998),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_2083),
.Y(n_2291)
);

BUFx4f_ASAP7_75t_L g2292 ( 
.A(n_2160),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_1993),
.B(n_2003),
.Y(n_2293)
);

BUFx2_ASAP7_75t_R g2294 ( 
.A(n_1961),
.Y(n_2294)
);

AO21x2_ASAP7_75t_L g2295 ( 
.A1(n_2004),
.A2(n_2149),
.B(n_1965),
.Y(n_2295)
);

INVx4_ASAP7_75t_L g2296 ( 
.A(n_2160),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_2083),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1992),
.B(n_2028),
.Y(n_2298)
);

AO21x2_ASAP7_75t_L g2299 ( 
.A1(n_2004),
.A2(n_2149),
.B(n_1965),
.Y(n_2299)
);

AO21x2_ASAP7_75t_L g2300 ( 
.A1(n_2159),
.A2(n_2181),
.B(n_2174),
.Y(n_2300)
);

BUFx12f_ASAP7_75t_L g2301 ( 
.A(n_2032),
.Y(n_2301)
);

OR2x6_ASAP7_75t_L g2302 ( 
.A(n_2005),
.B(n_2014),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1959),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2079),
.B(n_2100),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2134),
.Y(n_2305)
);

CKINVDCx6p67_ASAP7_75t_R g2306 ( 
.A(n_2072),
.Y(n_2306)
);

BUFx12f_ASAP7_75t_L g2307 ( 
.A(n_2155),
.Y(n_2307)
);

OA21x2_ASAP7_75t_L g2308 ( 
.A1(n_2028),
.A2(n_2071),
.B(n_2062),
.Y(n_2308)
);

OAI21xp33_ASAP7_75t_SL g2309 ( 
.A1(n_2130),
.A2(n_2145),
.B(n_2146),
.Y(n_2309)
);

CKINVDCx11_ASAP7_75t_R g2310 ( 
.A(n_2045),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2150),
.A2(n_2143),
.B1(n_2104),
.B2(n_2037),
.Y(n_2311)
);

AOI22x1_ASAP7_75t_SL g2312 ( 
.A1(n_1966),
.A2(n_2045),
.B1(n_2164),
.B2(n_2131),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_2135),
.A2(n_2141),
.B1(n_2143),
.B2(n_2148),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_SL g2314 ( 
.A1(n_2066),
.A2(n_1954),
.B1(n_2172),
.B2(n_2088),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2118),
.Y(n_2315)
);

AOI21x1_ASAP7_75t_L g2316 ( 
.A1(n_2140),
.A2(n_2162),
.B(n_2106),
.Y(n_2316)
);

BUFx8_ASAP7_75t_L g2317 ( 
.A(n_2048),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2120),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_2156),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_SL g2320 ( 
.A1(n_2127),
.A2(n_2042),
.B1(n_2066),
.B2(n_2013),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2064),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2064),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2022),
.B(n_2000),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_2064),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2132),
.B(n_2153),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_2170),
.Y(n_2326)
);

CKINVDCx11_ASAP7_75t_R g2327 ( 
.A(n_2108),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2040),
.B(n_2043),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2165),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2022),
.B(n_2000),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2083),
.Y(n_2331)
);

CKINVDCx6p67_ASAP7_75t_R g2332 ( 
.A(n_2072),
.Y(n_2332)
);

AOI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2124),
.A2(n_2158),
.B(n_2054),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2042),
.Y(n_2334)
);

OAI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2117),
.A2(n_2039),
.B1(n_2003),
.B2(n_2138),
.Y(n_2335)
);

NAND2x1p5_ASAP7_75t_L g2336 ( 
.A(n_2085),
.B(n_2129),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2142),
.Y(n_2337)
);

OA21x2_ASAP7_75t_L g2338 ( 
.A1(n_2161),
.A2(n_2171),
.B(n_1972),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2310),
.Y(n_2339)
);

OR2x6_ASAP7_75t_L g2340 ( 
.A(n_2195),
.B(n_2055),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2212),
.Y(n_2341)
);

INVx1_ASAP7_75t_SL g2342 ( 
.A(n_2279),
.Y(n_2342)
);

NOR3xp33_ASAP7_75t_SL g2343 ( 
.A(n_2202),
.B(n_2114),
.C(n_2135),
.Y(n_2343)
);

INVx4_ASAP7_75t_SL g2344 ( 
.A(n_2258),
.Y(n_2344)
);

OAI21xp33_ASAP7_75t_L g2345 ( 
.A1(n_2209),
.A2(n_2142),
.B(n_2114),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2214),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2201),
.B(n_2006),
.Y(n_2347)
);

CKINVDCx16_ASAP7_75t_R g2348 ( 
.A(n_2194),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2207),
.B(n_2026),
.Y(n_2349)
);

NAND2xp33_ASAP7_75t_R g2350 ( 
.A(n_2312),
.B(n_1983),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2207),
.B(n_2011),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2292),
.Y(n_2352)
);

CKINVDCx16_ASAP7_75t_R g2353 ( 
.A(n_2259),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_SL g2354 ( 
.A(n_2225),
.B(n_2061),
.C(n_2008),
.Y(n_2354)
);

AND2x4_ASAP7_75t_SL g2355 ( 
.A(n_2259),
.B(n_2164),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_2196),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2230),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2264),
.B(n_2085),
.Y(n_2358)
);

NOR2x1_ASAP7_75t_SL g2359 ( 
.A(n_2302),
.B(n_2085),
.Y(n_2359)
);

CKINVDCx16_ASAP7_75t_R g2360 ( 
.A(n_2287),
.Y(n_2360)
);

CKINVDCx16_ASAP7_75t_R g2361 ( 
.A(n_2301),
.Y(n_2361)
);

AOI22xp33_ASAP7_75t_SL g2362 ( 
.A1(n_2195),
.A2(n_2013),
.B1(n_2119),
.B2(n_2021),
.Y(n_2362)
);

A2O1A1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2266),
.A2(n_2128),
.B(n_2008),
.C(n_1972),
.Y(n_2363)
);

AOI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2203),
.A2(n_2150),
.B1(n_2096),
.B2(n_2138),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_SL g2365 ( 
.A(n_2245),
.B(n_2061),
.C(n_1974),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2292),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2216),
.B(n_2119),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2216),
.B(n_2123),
.Y(n_2368)
);

NAND2xp33_ASAP7_75t_R g2369 ( 
.A(n_2302),
.B(n_2030),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_2208),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2222),
.B(n_2013),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_2279),
.Y(n_2372)
);

NOR2x1p5_ASAP7_75t_L g2373 ( 
.A(n_2306),
.B(n_2057),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2270),
.B(n_2075),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2283),
.Y(n_2375)
);

CKINVDCx20_ASAP7_75t_R g2376 ( 
.A(n_2317),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2228),
.Y(n_2377)
);

NAND2xp33_ASAP7_75t_R g2378 ( 
.A(n_2302),
.B(n_2017),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2328),
.B(n_2165),
.Y(n_2379)
);

NAND3xp33_ASAP7_75t_SL g2380 ( 
.A(n_2267),
.B(n_2055),
.C(n_2092),
.Y(n_2380)
);

INVx1_ASAP7_75t_SL g2381 ( 
.A(n_2236),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2218),
.B(n_2030),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2240),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2273),
.Y(n_2384)
);

NOR3xp33_ASAP7_75t_SL g2385 ( 
.A(n_2232),
.B(n_1974),
.C(n_2099),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2290),
.B(n_1994),
.Y(n_2386)
);

INVxp67_ASAP7_75t_L g2387 ( 
.A(n_2191),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2242),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2258),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2288),
.B(n_1994),
.Y(n_2390)
);

OAI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2323),
.A2(n_2103),
.B(n_2092),
.Y(n_2391)
);

INVx8_ASAP7_75t_L g2392 ( 
.A(n_2307),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_R g2393 ( 
.A(n_2283),
.B(n_2029),
.Y(n_2393)
);

HB1xp67_ASAP7_75t_L g2394 ( 
.A(n_2204),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2246),
.Y(n_2395)
);

OR2x6_ASAP7_75t_L g2396 ( 
.A(n_2244),
.B(n_2017),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2204),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2188),
.B(n_1976),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2200),
.B(n_1986),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2223),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2200),
.B(n_1986),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2192),
.B(n_2034),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2293),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2190),
.B(n_2198),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_2239),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2224),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2256),
.B(n_2096),
.Y(n_2407)
);

OR2x2_ASAP7_75t_SL g2408 ( 
.A(n_2285),
.B(n_2099),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_SL g2409 ( 
.A1(n_2320),
.A2(n_2010),
.B(n_2151),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2197),
.B(n_2132),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2226),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2227),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_SL g2413 ( 
.A(n_2243),
.B(n_2036),
.C(n_2103),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2233),
.B(n_2085),
.Y(n_2414)
);

OR2x4_ASAP7_75t_L g2415 ( 
.A(n_2325),
.B(n_2221),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_SL g2416 ( 
.A(n_2255),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2336),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2231),
.B(n_2036),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_SL g2419 ( 
.A1(n_2193),
.A2(n_2038),
.B1(n_2020),
.B2(n_2122),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_R g2420 ( 
.A(n_2317),
.B(n_2129),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_R g2421 ( 
.A(n_2332),
.B(n_2129),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_R g2422 ( 
.A(n_2268),
.B(n_2129),
.Y(n_2422)
);

INVx2_ASAP7_75t_SL g2423 ( 
.A(n_2215),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2329),
.B(n_2098),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2252),
.Y(n_2425)
);

OAI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_2219),
.A2(n_2046),
.B1(n_2041),
.B2(n_2089),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2266),
.B(n_2059),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2327),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2336),
.Y(n_2429)
);

NAND2xp33_ASAP7_75t_SL g2430 ( 
.A(n_2213),
.B(n_2038),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2281),
.Y(n_2431)
);

AOI22xp33_ASAP7_75t_SL g2432 ( 
.A1(n_2314),
.A2(n_2020),
.B1(n_2058),
.B2(n_2059),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2294),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2330),
.B(n_2058),
.Y(n_2434)
);

NAND2xp33_ASAP7_75t_SL g2435 ( 
.A(n_2213),
.B(n_1963),
.Y(n_2435)
);

OR2x6_ASAP7_75t_L g2436 ( 
.A(n_2244),
.B(n_2111),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2253),
.Y(n_2437)
);

NAND2x1p5_ASAP7_75t_L g2438 ( 
.A(n_2296),
.B(n_1963),
.Y(n_2438)
);

BUFx12f_ASAP7_75t_L g2439 ( 
.A(n_2296),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2236),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2330),
.B(n_2080),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2305),
.B(n_2080),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2254),
.Y(n_2443)
);

INVx5_ASAP7_75t_L g2444 ( 
.A(n_2269),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_R g2445 ( 
.A(n_2250),
.B(n_2081),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2256),
.B(n_2181),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_L g2447 ( 
.A(n_2372),
.Y(n_2447)
);

CKINVDCx20_ASAP7_75t_R g2448 ( 
.A(n_2376),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2394),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2397),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2441),
.Y(n_2451)
);

AOI33xp33_ASAP7_75t_L g2452 ( 
.A1(n_2341),
.A2(n_2262),
.A3(n_2210),
.B1(n_2320),
.B2(n_2271),
.B3(n_2249),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2424),
.B(n_2282),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2407),
.B(n_2282),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2357),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2346),
.Y(n_2456)
);

BUFx2_ASAP7_75t_L g2457 ( 
.A(n_2340),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2403),
.B(n_2257),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2422),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2342),
.B(n_2298),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2407),
.B(n_2189),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2434),
.B(n_2427),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2342),
.B(n_2298),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2414),
.B(n_2365),
.Y(n_2464)
);

NOR2x1_ASAP7_75t_L g2465 ( 
.A(n_2409),
.B(n_2272),
.Y(n_2465)
);

AOI221xp5_ASAP7_75t_L g2466 ( 
.A1(n_2409),
.A2(n_2335),
.B1(n_2284),
.B2(n_2277),
.C(n_2309),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2340),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2345),
.A2(n_2313),
.B1(n_2260),
.B2(n_2271),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2377),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2383),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2388),
.B(n_2263),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2395),
.B(n_2263),
.Y(n_2472)
);

NOR2x1_ASAP7_75t_L g2473 ( 
.A(n_2405),
.B(n_2220),
.Y(n_2473)
);

AOI22x1_ASAP7_75t_L g2474 ( 
.A1(n_2353),
.A2(n_2314),
.B1(n_2220),
.B2(n_2250),
.Y(n_2474)
);

HB1xp67_ASAP7_75t_L g2475 ( 
.A(n_2440),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2384),
.B(n_2295),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2446),
.B(n_2299),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2400),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2340),
.B(n_2261),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2406),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2446),
.B(n_2299),
.Y(n_2481)
);

AND2x2_ASAP7_75t_SL g2482 ( 
.A(n_2414),
.B(n_2261),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2381),
.B(n_2257),
.Y(n_2483)
);

OR2x6_ASAP7_75t_L g2484 ( 
.A(n_2396),
.B(n_2217),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2411),
.B(n_2286),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2412),
.B(n_2286),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2381),
.B(n_2217),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2425),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_L g2489 ( 
.A1(n_2345),
.A2(n_2260),
.B1(n_2247),
.B2(n_2276),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2391),
.B(n_2300),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2391),
.B(n_2300),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2437),
.Y(n_2492)
);

INVxp67_ASAP7_75t_SL g2493 ( 
.A(n_2399),
.Y(n_2493)
);

INVxp67_ASAP7_75t_SL g2494 ( 
.A(n_2401),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2443),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2404),
.B(n_2275),
.Y(n_2496)
);

HB1xp67_ASAP7_75t_L g2497 ( 
.A(n_2382),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2349),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2386),
.B(n_2308),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2444),
.Y(n_2500)
);

OR2x2_ASAP7_75t_L g2501 ( 
.A(n_2418),
.B(n_2238),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2396),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2426),
.Y(n_2503)
);

HB1xp67_ASAP7_75t_L g2504 ( 
.A(n_2379),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2436),
.B(n_2333),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2456),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2485),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2485),
.Y(n_2508)
);

INVxp67_ASAP7_75t_SL g2509 ( 
.A(n_2450),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2453),
.B(n_2343),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2471),
.B(n_2472),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2471),
.B(n_2472),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2456),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2453),
.B(n_2419),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2486),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2451),
.B(n_2363),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2449),
.Y(n_2517)
);

OAI21xp33_ASAP7_75t_L g2518 ( 
.A1(n_2465),
.A2(n_2362),
.B(n_2354),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2460),
.B(n_2351),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2499),
.B(n_2248),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2502),
.B(n_2396),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2499),
.B(n_2248),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2460),
.B(n_2367),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2454),
.B(n_2432),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2454),
.B(n_2316),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2451),
.B(n_2390),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2463),
.B(n_2483),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2486),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2448),
.B(n_2389),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2458),
.B(n_2368),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2461),
.B(n_2251),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2463),
.B(n_2483),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2447),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2455),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2449),
.B(n_2371),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2493),
.B(n_2364),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_2501),
.B(n_2426),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2494),
.B(n_2442),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2501),
.B(n_2413),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2520),
.B(n_2462),
.Y(n_2540)
);

BUFx2_ASAP7_75t_SL g2541 ( 
.A(n_2517),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2517),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2520),
.B(n_2462),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2522),
.B(n_2487),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2534),
.Y(n_2545)
);

INVx3_ASAP7_75t_L g2546 ( 
.A(n_2521),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2527),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_2539),
.B(n_2473),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2510),
.B(n_2490),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2521),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_2527),
.B(n_2476),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2522),
.B(n_2487),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2507),
.B(n_2508),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2507),
.B(n_2508),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2515),
.B(n_2528),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2510),
.B(n_2490),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2515),
.B(n_2477),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2506),
.Y(n_2558)
);

NAND2x1_ASAP7_75t_SL g2559 ( 
.A(n_2521),
.B(n_2505),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2506),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2532),
.B(n_2476),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2528),
.B(n_2477),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2525),
.B(n_2481),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2513),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2532),
.B(n_2498),
.Y(n_2565)
);

INVx1_ASAP7_75t_SL g2566 ( 
.A(n_2519),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2525),
.B(n_2481),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2533),
.B(n_2361),
.Y(n_2568)
);

OAI322xp33_ASAP7_75t_L g2569 ( 
.A1(n_2549),
.A2(n_2539),
.A3(n_2519),
.B1(n_2535),
.B2(n_2537),
.C1(n_2530),
.C2(n_2512),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2547),
.Y(n_2570)
);

BUFx2_ASAP7_75t_L g2571 ( 
.A(n_2542),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_SL g2572 ( 
.A1(n_2541),
.A2(n_2482),
.B1(n_2459),
.B2(n_2467),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_SL g2573 ( 
.A(n_2548),
.B(n_2474),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2547),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2565),
.Y(n_2575)
);

AOI32xp33_ASAP7_75t_L g2576 ( 
.A1(n_2548),
.A2(n_2518),
.A3(n_2459),
.B1(n_2509),
.B2(n_2467),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2545),
.Y(n_2577)
);

AOI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2549),
.A2(n_2524),
.B1(n_2514),
.B2(n_2464),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2565),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2568),
.B(n_2356),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2542),
.B(n_2474),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2558),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2558),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2566),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2546),
.B(n_2502),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2540),
.B(n_2497),
.Y(n_2586)
);

NAND3xp33_ASAP7_75t_L g2587 ( 
.A(n_2556),
.B(n_2452),
.C(n_2387),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2545),
.Y(n_2588)
);

OR2x6_ASAP7_75t_L g2589 ( 
.A(n_2541),
.B(n_2457),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2551),
.B(n_2511),
.Y(n_2590)
);

INVxp67_ASAP7_75t_SL g2591 ( 
.A(n_2545),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2566),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2560),
.Y(n_2593)
);

NAND4xp25_ASAP7_75t_L g2594 ( 
.A(n_2556),
.B(n_2350),
.C(n_2206),
.D(n_2468),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2563),
.A2(n_2524),
.B1(n_2514),
.B2(n_2516),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2560),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2546),
.B(n_2457),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2540),
.B(n_2531),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2564),
.Y(n_2599)
);

OA222x2_ASAP7_75t_L g2600 ( 
.A1(n_2546),
.A2(n_2484),
.B1(n_2535),
.B2(n_2538),
.C1(n_2366),
.C2(n_2352),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_2551),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2582),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2576),
.B(n_2466),
.C(n_2529),
.Y(n_2603)
);

OAI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2587),
.A2(n_2380),
.B(n_2229),
.Y(n_2604)
);

O2A1O1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_2594),
.A2(n_2237),
.B(n_2211),
.C(n_2205),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2595),
.B(n_2563),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2570),
.B(n_2567),
.Y(n_2607)
);

OAI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2594),
.A2(n_2546),
.B1(n_2550),
.B2(n_2484),
.Y(n_2608)
);

OAI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2589),
.A2(n_2550),
.B1(n_2484),
.B2(n_2561),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2601),
.B(n_2561),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2581),
.A2(n_2482),
.B(n_2359),
.Y(n_2611)
);

OAI21xp33_ASAP7_75t_SL g2612 ( 
.A1(n_2589),
.A2(n_2559),
.B(n_2543),
.Y(n_2612)
);

NOR2x1_ASAP7_75t_L g2613 ( 
.A(n_2589),
.B(n_2373),
.Y(n_2613)
);

OAI21xp33_ASAP7_75t_L g2614 ( 
.A1(n_2578),
.A2(n_2559),
.B(n_2552),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2583),
.Y(n_2615)
);

AOI21xp33_ASAP7_75t_SL g2616 ( 
.A1(n_2587),
.A2(n_2392),
.B(n_2360),
.Y(n_2616)
);

OAI221xp5_ASAP7_75t_L g2617 ( 
.A1(n_2572),
.A2(n_2550),
.B1(n_2536),
.B2(n_2489),
.C(n_2385),
.Y(n_2617)
);

OAI21xp33_ASAP7_75t_L g2618 ( 
.A1(n_2601),
.A2(n_2552),
.B(n_2544),
.Y(n_2618)
);

AOI211xp5_ASAP7_75t_L g2619 ( 
.A1(n_2569),
.A2(n_2393),
.B(n_2420),
.C(n_2433),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2593),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2596),
.Y(n_2621)
);

OAI322xp33_ASAP7_75t_L g2622 ( 
.A1(n_2608),
.A2(n_2573),
.A3(n_2574),
.B1(n_2579),
.B2(n_2575),
.C1(n_2584),
.C2(n_2592),
.Y(n_2622)
);

AOI221xp5_ASAP7_75t_L g2623 ( 
.A1(n_2616),
.A2(n_2571),
.B1(n_2591),
.B2(n_2599),
.C(n_2580),
.Y(n_2623)
);

NAND2x1p5_ASAP7_75t_L g2624 ( 
.A(n_2613),
.B(n_2431),
.Y(n_2624)
);

OAI211xp5_ASAP7_75t_L g2625 ( 
.A1(n_2619),
.A2(n_2421),
.B(n_2392),
.C(n_2370),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2610),
.Y(n_2626)
);

OR2x2_ASAP7_75t_L g2627 ( 
.A(n_2607),
.B(n_2590),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2612),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2603),
.A2(n_2573),
.B1(n_2439),
.B2(n_2374),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2618),
.B(n_2600),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2614),
.B(n_2598),
.Y(n_2631)
);

AOI222xp33_ASAP7_75t_L g2632 ( 
.A1(n_2617),
.A2(n_2597),
.B1(n_2544),
.B2(n_2586),
.C1(n_2567),
.C2(n_2344),
.Y(n_2632)
);

OR2x2_ASAP7_75t_L g2633 ( 
.A(n_2606),
.B(n_2543),
.Y(n_2633)
);

OAI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2611),
.A2(n_2597),
.B1(n_2408),
.B2(n_2550),
.Y(n_2634)
);

INVx1_ASAP7_75t_SL g2635 ( 
.A(n_2602),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2615),
.Y(n_2636)
);

OAI21xp33_ASAP7_75t_L g2637 ( 
.A1(n_2604),
.A2(n_2588),
.B(n_2577),
.Y(n_2637)
);

OR2x2_ASAP7_75t_L g2638 ( 
.A(n_2620),
.B(n_2557),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2621),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2609),
.B(n_2557),
.Y(n_2640)
);

OAI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2604),
.A2(n_2415),
.B1(n_2585),
.B2(n_2504),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2605),
.A2(n_2585),
.B1(n_2553),
.B2(n_2348),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2610),
.Y(n_2643)
);

XOR2xp5_ASAP7_75t_L g2644 ( 
.A(n_2629),
.B(n_2428),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2624),
.B(n_2625),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2635),
.B(n_2475),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2626),
.B(n_2562),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2628),
.B(n_2554),
.Y(n_2648)
);

AOI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2634),
.A2(n_2392),
.B(n_2375),
.Y(n_2649)
);

OAI21xp5_ASAP7_75t_SL g2650 ( 
.A1(n_2629),
.A2(n_2355),
.B(n_2229),
.Y(n_2650)
);

A2O1A1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2628),
.A2(n_2339),
.B(n_2265),
.C(n_2234),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2643),
.Y(n_2652)
);

O2A1O1Ixp33_ASAP7_75t_L g2653 ( 
.A1(n_2637),
.A2(n_2199),
.B(n_2423),
.C(n_2235),
.Y(n_2653)
);

NAND3xp33_ASAP7_75t_SL g2654 ( 
.A(n_2632),
.B(n_2438),
.C(n_2445),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2630),
.A2(n_2537),
.B1(n_2484),
.B2(n_2523),
.Y(n_2655)
);

OAI21xp33_ASAP7_75t_L g2656 ( 
.A1(n_2637),
.A2(n_2526),
.B(n_2491),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2642),
.A2(n_2358),
.B(n_2435),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2633),
.B(n_2562),
.Y(n_2658)
);

AOI221xp5_ASAP7_75t_L g2659 ( 
.A1(n_2622),
.A2(n_2553),
.B1(n_2478),
.B2(n_2470),
.C(n_2469),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2636),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2652),
.Y(n_2661)
);

NOR3xp33_ASAP7_75t_L g2662 ( 
.A(n_2650),
.B(n_2622),
.C(n_2641),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_SL g2663 ( 
.A1(n_2645),
.A2(n_2631),
.B1(n_2500),
.B2(n_2319),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2644),
.B(n_2623),
.Y(n_2664)
);

OAI21xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2659),
.A2(n_2640),
.B(n_2627),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2646),
.Y(n_2666)
);

NOR2x1_ASAP7_75t_L g2667 ( 
.A(n_2649),
.B(n_2326),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2660),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2651),
.A2(n_2639),
.B(n_2638),
.Y(n_2669)
);

NAND3xp33_ASAP7_75t_L g2670 ( 
.A(n_2655),
.B(n_2334),
.C(n_2318),
.Y(n_2670)
);

NOR3xp33_ASAP7_75t_L g2671 ( 
.A(n_2654),
.B(n_2324),
.C(n_2315),
.Y(n_2671)
);

AOI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2653),
.A2(n_2264),
.B(n_2311),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_SL g2673 ( 
.A1(n_2657),
.A2(n_2344),
.B(n_2311),
.Y(n_2673)
);

OAI211xp5_ASAP7_75t_SL g2674 ( 
.A1(n_2656),
.A2(n_2249),
.B(n_2337),
.C(n_2321),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2648),
.Y(n_2675)
);

AOI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2658),
.A2(n_2416),
.B1(n_2378),
.B2(n_2369),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_R g2677 ( 
.A(n_2664),
.B(n_2416),
.Y(n_2677)
);

AOI221xp5_ASAP7_75t_L g2678 ( 
.A1(n_2662),
.A2(n_2647),
.B1(n_2347),
.B2(n_2470),
.C(n_2478),
.Y(n_2678)
);

O2A1O1Ixp5_ASAP7_75t_SL g2679 ( 
.A1(n_2668),
.A2(n_2322),
.B(n_2215),
.C(n_2303),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2675),
.A2(n_2491),
.B1(n_2505),
.B2(n_2479),
.Y(n_2680)
);

INVx1_ASAP7_75t_SL g2681 ( 
.A(n_2667),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2661),
.A2(n_2402),
.B(n_2294),
.C(n_2304),
.Y(n_2682)
);

NAND4xp25_ASAP7_75t_L g2683 ( 
.A(n_2663),
.B(n_2410),
.C(n_2500),
.D(n_2241),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2666),
.Y(n_2684)
);

OAI221xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2665),
.A2(n_2241),
.B1(n_2523),
.B2(n_2436),
.C(n_2503),
.Y(n_2685)
);

AOI322xp5_ASAP7_75t_L g2686 ( 
.A1(n_2676),
.A2(n_2671),
.A3(n_2673),
.B1(n_2674),
.B2(n_2553),
.C1(n_2554),
.C2(n_2555),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2669),
.B(n_2555),
.Y(n_2687)
);

NAND4xp75_ASAP7_75t_L g2688 ( 
.A(n_2672),
.B(n_2398),
.C(n_2289),
.D(n_2338),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2684),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2687),
.B(n_2670),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2681),
.Y(n_2691)
);

NOR2x1_ASAP7_75t_L g2692 ( 
.A(n_2683),
.B(n_2417),
.Y(n_2692)
);

NAND2x1p5_ASAP7_75t_L g2693 ( 
.A(n_2677),
.B(n_2444),
.Y(n_2693)
);

AO22x2_ASAP7_75t_SL g2694 ( 
.A1(n_2685),
.A2(n_2417),
.B1(n_2429),
.B2(n_2303),
.Y(n_2694)
);

AO22x2_ASAP7_75t_L g2695 ( 
.A1(n_2688),
.A2(n_2331),
.B1(n_2480),
.B2(n_2429),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_2682),
.B(n_2678),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2686),
.B(n_2553),
.Y(n_2697)
);

NOR2x1_ASAP7_75t_L g2698 ( 
.A(n_2679),
.B(n_2480),
.Y(n_2698)
);

NOR2x1_ASAP7_75t_L g2699 ( 
.A(n_2680),
.B(n_2269),
.Y(n_2699)
);

NAND4xp75_ASAP7_75t_L g2700 ( 
.A(n_2691),
.B(n_2338),
.C(n_2503),
.D(n_2496),
.Y(n_2700)
);

OAI221xp5_ASAP7_75t_L g2701 ( 
.A1(n_2693),
.A2(n_2444),
.B1(n_2430),
.B2(n_2492),
.C(n_2488),
.Y(n_2701)
);

NAND4xp75_ASAP7_75t_L g2702 ( 
.A(n_2692),
.B(n_2488),
.C(n_2492),
.D(n_2495),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2689),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2690),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2698),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2696),
.B(n_2495),
.Y(n_2706)
);

NOR2x1_ASAP7_75t_L g2707 ( 
.A(n_2697),
.B(n_2274),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2704),
.B(n_2699),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_2703),
.Y(n_2709)
);

CKINVDCx20_ASAP7_75t_R g2710 ( 
.A(n_2706),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2708),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_L g2712 ( 
.A1(n_2711),
.A2(n_2707),
.B1(n_2694),
.B2(n_2710),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_2712),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2713),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2714),
.A2(n_2709),
.B1(n_2705),
.B2(n_2700),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2715),
.A2(n_2695),
.B1(n_2701),
.B2(n_2702),
.Y(n_2716)
);

AOI221xp5_ASAP7_75t_L g2717 ( 
.A1(n_2716),
.A2(n_2695),
.B1(n_2280),
.B2(n_2278),
.C(n_2297),
.Y(n_2717)
);

AOI211xp5_ASAP7_75t_L g2718 ( 
.A1(n_2717),
.A2(n_2291),
.B(n_2297),
.C(n_2274),
.Y(n_2718)
);


endmodule