module fake_jpeg_29980_n_65 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_65);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_5),
.B(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_18),
.C(n_16),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_13),
.C(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_13),
.B(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_24),
.B1(n_10),
.B2(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_43),
.B1(n_34),
.B2(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_42),
.A3(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_34),
.B2(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_19),
.B1(n_34),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_45),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_3),
.C(n_7),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_52),
.B1(n_46),
.B2(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_0),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_2),
.Y(n_64)
);

NAND2x1_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_2),
.Y(n_65)
);


endmodule