module fake_jpeg_21893_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_47),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_47),
.B1(n_45),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_36),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_61),
.B1(n_19),
.B2(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_19),
.B1(n_36),
.B2(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_77),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_71),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_74),
.B1(n_97),
.B2(n_48),
.Y(n_105)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_39),
.B1(n_47),
.B2(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_78),
.B1(n_93),
.B2(n_42),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_31),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_47),
.B1(n_25),
.B2(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_81),
.Y(n_106)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_84),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_24),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_18),
.B1(n_17),
.B2(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_48),
.B1(n_46),
.B2(n_42),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_70),
.B1(n_98),
.B2(n_68),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_104),
.B1(n_108),
.B2(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_81),
.B1(n_66),
.B2(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_112),
.B1(n_126),
.B2(n_86),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_40),
.B1(n_37),
.B2(n_44),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_71),
.B1(n_69),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_124),
.B1(n_30),
.B2(n_28),
.Y(n_149)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_41),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_17),
.B1(n_40),
.B2(n_37),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_131),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_137),
.B1(n_144),
.B2(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_139),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_40),
.B(n_67),
.C(n_37),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_138),
.B(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_96),
.B1(n_72),
.B2(n_90),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_44),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_95),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_91),
.B1(n_89),
.B2(n_23),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_114),
.B1(n_128),
.B2(n_129),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_44),
.B1(n_85),
.B2(n_43),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_44),
.B1(n_85),
.B2(n_43),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_43),
.C(n_41),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_126),
.C(n_123),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_103),
.B1(n_28),
.B2(n_30),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_41),
.B1(n_23),
.B2(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_151),
.B1(n_157),
.B2(n_101),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_124),
.B1(n_108),
.B2(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_26),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_41),
.B1(n_23),
.B2(n_20),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_121),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_179),
.B(n_27),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_165),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_175),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_168),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_155),
.B1(n_134),
.B2(n_138),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_171),
.B1(n_174),
.B2(n_157),
.Y(n_192)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_107),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_110),
.B(n_123),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_182),
.B(n_35),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_103),
.C(n_94),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_184),
.B1(n_137),
.B2(n_141),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_101),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_151),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_119),
.B(n_109),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_111),
.B1(n_99),
.B2(n_30),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_99),
.C(n_111),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_186),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_99),
.C(n_107),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_107),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_150),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_164),
.C(n_160),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_135),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_198),
.B(n_201),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_192),
.A2(n_199),
.B1(n_203),
.B2(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_149),
.B1(n_141),
.B2(n_131),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_207),
.B1(n_214),
.B2(n_9),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_143),
.B1(n_26),
.B2(n_34),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_20),
.B1(n_28),
.B2(n_33),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_35),
.B1(n_27),
.B2(n_21),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_208),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_33),
.B1(n_136),
.B2(n_32),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_33),
.B1(n_136),
.B2(n_32),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_131),
.B1(n_29),
.B2(n_35),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_219),
.B(n_181),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_161),
.CI(n_172),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_217),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_213),
.B(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_29),
.B1(n_35),
.B2(n_27),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_158),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_27),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_160),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_21),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_189),
.Y(n_235)
);

NAND2x1_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_0),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_166),
.B1(n_187),
.B2(n_178),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_222),
.B(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_233),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_231),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_201),
.B(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_164),
.B(n_181),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_209),
.B(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_205),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_159),
.C(n_169),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_0),
.C(n_1),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_0),
.C(n_1),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_1),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_201),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_207),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_221),
.B1(n_194),
.B2(n_198),
.Y(n_255)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_235),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_258),
.B(n_263),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_266),
.B1(n_245),
.B2(n_228),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_256),
.B1(n_10),
.B2(n_14),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_211),
.B1(n_215),
.B2(n_205),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_223),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_220),
.B(n_215),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_214),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_9),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_243),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_229),
.B1(n_227),
.B2(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_236),
.C(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_274),
.C(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_263),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_261),
.C(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_224),
.C(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_246),
.B1(n_242),
.B2(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_230),
.C(n_242),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_283),
.C(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_237),
.B1(n_225),
.B2(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_237),
.C(n_247),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_10),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_266),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_285),
.B1(n_283),
.B2(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_249),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_16),
.B(n_13),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_248),
.B1(n_265),
.B2(n_262),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_300),
.B1(n_270),
.B2(n_282),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_272),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_16),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_264),
.B1(n_253),
.B2(n_5),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_274),
.B(n_271),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_302),
.A2(n_297),
.B(n_4),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_273),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_275),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_3),
.C(n_4),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_291),
.C(n_296),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_290),
.C(n_301),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_294),
.B(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_317),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_298),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_12),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_12),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_310),
.Y(n_322)
);

AOI221xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_308),
.B1(n_303),
.B2(n_307),
.C(n_11),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_303),
.B1(n_312),
.B2(n_309),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_324),
.A2(n_316),
.B(n_314),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_328),
.B(n_315),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_16),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_318),
.B(n_4),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_329),
.B(n_333),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_323),
.B(n_332),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_330),
.B(n_6),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_3),
.B(n_6),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B(n_7),
.Y(n_341)
);


endmodule