module fake_jpeg_811_n_508 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_50),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_52),
.Y(n_141)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_75),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_87),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_89),
.Y(n_122)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_95),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_100),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_35),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_30),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_46),
.B1(n_18),
.B2(n_25),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_70),
.B1(n_77),
.B2(n_73),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_18),
.B1(n_40),
.B2(n_35),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_124),
.B1(n_138),
.B2(n_144),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_51),
.A2(n_18),
.B1(n_40),
.B2(n_35),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_40),
.B1(n_46),
.B2(n_29),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_137),
.B1(n_142),
.B2(n_66),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_68),
.A2(n_40),
.B1(n_47),
.B2(n_38),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_136),
.A2(n_0),
.B(n_2),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_39),
.B1(n_34),
.B2(n_15),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_39),
.B1(n_34),
.B2(n_38),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_15),
.B1(n_19),
.B2(n_44),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_62),
.A2(n_47),
.B1(n_26),
.B2(n_21),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_20),
.B1(n_96),
.B2(n_80),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_158),
.B1(n_57),
.B2(n_86),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_63),
.B(n_19),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_161),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_74),
.A2(n_49),
.B1(n_50),
.B2(n_88),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_78),
.B(n_44),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_98),
.C(n_97),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_189),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_168),
.A2(n_185),
.B1(n_197),
.B2(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_20),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_178),
.B1(n_184),
.B2(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_54),
.B1(n_76),
.B2(n_60),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_181),
.Y(n_220)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_0),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_83),
.B1(n_71),
.B2(n_69),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_190),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_65),
.B1(n_45),
.B2(n_3),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_141),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_121),
.A2(n_139),
.B1(n_156),
.B2(n_112),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_204),
.B1(n_155),
.B2(n_112),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_196),
.Y(n_237)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_142),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_110),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_201),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_45),
.B(n_9),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_110),
.B(n_145),
.C(n_105),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_0),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_103),
.B(n_14),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_207),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_136),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_3),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_223),
.B1(n_232),
.B2(n_145),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_152),
.B1(n_129),
.B2(n_135),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_171),
.B(n_148),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_160),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_199),
.B(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_174),
.B(n_135),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_146),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_185),
.A2(n_108),
.B1(n_113),
.B2(n_107),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_166),
.B1(n_199),
.B2(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_194),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_230),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_166),
.B1(n_175),
.B2(n_168),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_264),
.B1(n_265),
.B2(n_268),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_200),
.B(n_205),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_240),
.B(n_244),
.Y(n_298)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_255),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_204),
.B1(n_187),
.B2(n_176),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_252),
.A2(n_269),
.B(n_273),
.Y(n_282)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_233),
.C(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_226),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_262),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_217),
.B1(n_240),
.B2(n_239),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_163),
.C(n_202),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_261),
.B(n_215),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_274),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_202),
.B1(n_201),
.B2(n_197),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_183),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_272),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_209),
.A2(n_173),
.B1(n_133),
.B2(n_104),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_228),
.A2(n_236),
.B1(n_223),
.B2(n_233),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_271),
.B1(n_275),
.B2(n_210),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_170),
.B1(n_162),
.B2(n_179),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_214),
.B(n_173),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_224),
.A2(n_207),
.B(n_169),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_194),
.B1(n_182),
.B2(n_181),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_214),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_286),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_267),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_281),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_258),
.B(n_241),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_252),
.A2(n_238),
.B1(n_212),
.B2(n_236),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_289),
.B1(n_292),
.B2(n_264),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_265),
.A2(n_212),
.B1(n_211),
.B2(n_225),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_235),
.B1(n_243),
.B2(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_302),
.B1(n_271),
.B2(n_275),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_301),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_303),
.B(n_304),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_270),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_300),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_244),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_301),
.B(n_280),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_248),
.A2(n_221),
.B1(n_177),
.B2(n_216),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_261),
.A2(n_216),
.B(n_215),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_246),
.A2(n_210),
.A3(n_220),
.B1(n_227),
.B2(n_180),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_269),
.Y(n_311)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_300),
.B1(n_269),
.B2(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_309),
.A2(n_285),
.B1(n_282),
.B2(n_306),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_310),
.A2(n_321),
.B1(n_322),
.B2(n_328),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_311),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_260),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_325),
.C(n_286),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_314),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_315),
.B(n_316),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_260),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_256),
.B(n_251),
.C(n_245),
.D(n_266),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_318),
.B(n_330),
.CI(n_303),
.CON(n_360),
.SN(n_360)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_277),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_329),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_248),
.B1(n_268),
.B2(n_259),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_256),
.C(n_246),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_249),
.B1(n_257),
.B2(n_254),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_270),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_249),
.C(n_165),
.Y(n_330)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_227),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_333),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_278),
.B(n_189),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_213),
.Y(n_334)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_287),
.A2(n_271),
.B1(n_250),
.B2(n_253),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_335),
.A2(n_338),
.B1(n_296),
.B2(n_302),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_298),
.A2(n_250),
.B(n_188),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_304),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_292),
.A2(n_221),
.B1(n_177),
.B2(n_210),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_340),
.A2(n_313),
.B(n_309),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_284),
.Y(n_343)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_346),
.B(n_362),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_288),
.Y(n_348)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_289),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_368),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_353),
.C(n_363),
.Y(n_371)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_281),
.C(n_299),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_321),
.B1(n_336),
.B2(n_317),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_305),
.B1(n_220),
.B2(n_229),
.Y(n_390)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_305),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_326),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_282),
.C(n_206),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_322),
.B1(n_318),
.B2(n_308),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_107),
.C(n_118),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_369),
.C(n_337),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_306),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_118),
.C(n_128),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_305),
.Y(n_370)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_343),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_372),
.B(n_392),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_328),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_382),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_340),
.A2(n_313),
.B(n_311),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_381),
.A2(n_395),
.B(n_370),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_330),
.Y(n_382)
);

XOR2x2_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_317),
.C(n_335),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_394),
.C(n_341),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_390),
.B1(n_344),
.B2(n_357),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_391),
.B(n_397),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_358),
.B(n_291),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_128),
.C(n_213),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_229),
.B(n_213),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_350),
.B(n_229),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_342),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_143),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_220),
.Y(n_398)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_398),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_410),
.Y(n_427)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_401),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_393),
.A2(n_361),
.B1(n_365),
.B2(n_359),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_402),
.A2(n_411),
.B1(n_384),
.B2(n_385),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_363),
.C(n_368),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_404),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_369),
.C(n_367),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_345),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_348),
.C(n_347),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_418),
.C(n_421),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_379),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_383),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_417),
.Y(n_426)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_360),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_416),
.B(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_356),
.C(n_357),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_352),
.B1(n_360),
.B2(n_344),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_420),
.A2(n_395),
.B1(n_384),
.B2(n_379),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_147),
.C(n_111),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_386),
.A2(n_111),
.B(n_106),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_422),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_424),
.A2(n_431),
.B1(n_106),
.B2(n_133),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_391),
.C(n_394),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_430),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_427),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_435),
.B1(n_400),
.B2(n_413),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_397),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_375),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_438),
.Y(n_452)
);

BUFx24_ASAP7_75t_SL g434 ( 
.A(n_406),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_436),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_376),
.B1(n_377),
.B2(n_389),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_373),
.C(n_376),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_9),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_147),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_445),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_440),
.B(n_418),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_427),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_456),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_442),
.A2(n_404),
.B(n_408),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_448),
.A2(n_449),
.B(n_423),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_441),
.A2(n_410),
.B(n_422),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_426),
.A2(n_416),
.B1(n_407),
.B2(n_421),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_453),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_409),
.C(n_407),
.Y(n_453)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_104),
.C(n_5),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_457),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_11),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_4),
.C(n_5),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_5),
.C(n_7),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_460),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_439),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_446),
.B(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_461),
.B(n_475),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_467),
.B(n_472),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_423),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_464),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_443),
.A2(n_9),
.B(n_12),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_460),
.A2(n_12),
.B(n_13),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_13),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_457),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_444),
.B(n_13),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_478),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_445),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_452),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_479),
.A2(n_484),
.B(n_485),
.Y(n_491)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_482),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_453),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_468),
.A2(n_455),
.B(n_459),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_469),
.A2(n_468),
.B(n_470),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_454),
.C(n_456),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_486),
.B(n_487),
.Y(n_488)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_465),
.B(n_467),
.Y(n_490)
);

AOI21x1_ASAP7_75t_SL g498 ( 
.A1(n_490),
.A2(n_492),
.B(n_494),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_466),
.B(n_14),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_14),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_486),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_497),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_493),
.A2(n_491),
.B(n_495),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_483),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_488),
.B(n_480),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_498),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_7),
.B(n_501),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_505),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_7),
.B(n_503),
.Y(n_508)
);


endmodule