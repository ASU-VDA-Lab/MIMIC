module fake_jpeg_15807_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_34),
.B1(n_26),
.B2(n_25),
.Y(n_102)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_20),
.B1(n_35),
.B2(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_1),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_3),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_3),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_28),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_86),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_36),
.B1(n_6),
.B2(n_7),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_71),
.A2(n_72),
.B1(n_80),
.B2(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_40),
.B1(n_23),
.B2(n_25),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_81),
.B(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_79),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_20),
.B1(n_39),
.B2(n_35),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_32),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_18),
.B1(n_17),
.B2(n_40),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_17),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_52),
.B(n_39),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_96),
.B1(n_71),
.B2(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_84),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_109),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_114),
.B1(n_120),
.B2(n_122),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_13),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_121),
.Y(n_141)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_125),
.Y(n_149)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_15),
.B1(n_104),
.B2(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_71),
.B1(n_101),
.B2(n_74),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_139),
.B1(n_134),
.B2(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_135),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_89),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_101),
.B1(n_74),
.B2(n_78),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_147),
.B1(n_161),
.B2(n_165),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_131),
.B(n_107),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_148),
.B(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_150),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_90),
.B(n_93),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_103),
.C(n_84),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_122),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_166),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_110),
.A2(n_118),
.B(n_119),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_110),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_113),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_162),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_134),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_164),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_127),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_152),
.C(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_133),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_112),
.B(n_123),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_161),
.B1(n_166),
.B2(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_167),
.Y(n_188)
);

AO221x1_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_189),
.B1(n_145),
.B2(n_156),
.C(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_143),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_199),
.C(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_185),
.B1(n_171),
.B2(n_172),
.Y(n_209)
);

CKINVDCx6p67_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_159),
.B(n_163),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_203),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_154),
.C(n_151),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_151),
.C(n_157),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_144),
.B(n_164),
.C(n_179),
.D(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_213),
.B1(n_217),
.B2(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_186),
.C(n_175),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_218),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_185),
.B1(n_178),
.B2(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_204),
.B(n_198),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_190),
.B1(n_201),
.B2(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_207),
.C(n_210),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_222),
.B1(n_223),
.B2(n_215),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_233),
.A2(n_222),
.B(n_215),
.C(n_226),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_231),
.B(n_194),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_234),
.B(n_235),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_237),
.Y(n_238)
);


endmodule