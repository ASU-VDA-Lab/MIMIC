module fake_jpeg_8081_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_51),
.B1(n_16),
.B2(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_32),
.B(n_18),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_61),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_34),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_80),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_62),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_65),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_69),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_25),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_71),
.Y(n_99)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_37),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_73),
.B(n_29),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_37),
.C(n_33),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_33),
.C(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_40),
.B1(n_15),
.B2(n_33),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_34),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_46),
.B1(n_52),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_84),
.B1(n_87),
.B2(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_52),
.B1(n_42),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_42),
.B1(n_40),
.B2(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_11),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_42),
.B1(n_43),
.B2(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_101),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_77),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_40),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_104),
.B1(n_63),
.B2(n_75),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_72),
.B1(n_74),
.B2(n_60),
.Y(n_104)
);

OAI22x1_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_30),
.B1(n_15),
.B2(n_17),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_110),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_117),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_67),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_76),
.B1(n_71),
.B2(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_89),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_78),
.B(n_66),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_15),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_100),
.C(n_91),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_125),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_30),
.B(n_25),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_11),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NOR4xp25_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_14),
.C(n_3),
.D(n_4),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_88),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_131),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_101),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_146),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_112),
.C(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_162),
.C(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_106),
.B(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_133),
.B1(n_102),
.B2(n_90),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_109),
.B1(n_107),
.B2(n_105),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_161),
.B1(n_129),
.B2(n_90),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_122),
.A3(n_109),
.B1(n_116),
.B2(n_110),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_30),
.B1(n_25),
.B2(n_17),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_143),
.B1(n_138),
.B2(n_145),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_140),
.B1(n_134),
.B2(n_116),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_55),
.B(n_3),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_173),
.C(n_175),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_160),
.B1(n_149),
.B2(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_151),
.C(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_17),
.B(n_55),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_136),
.C(n_94),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_151),
.C(n_150),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_180),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_150),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_181),
.B(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_174),
.B1(n_4),
.B2(n_6),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_172),
.B(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_14),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_R g187 ( 
.A(n_178),
.B(n_170),
.Y(n_187)
);

OAI221xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_7),
.B1(n_9),
.B2(n_186),
.C(n_188),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_190),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_7),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_2),
.C(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_7),
.C(n_9),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_190),
.B(n_9),
.CI(n_6),
.CON(n_194),
.SN(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_196),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_6),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_199),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_192),
.B(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_195),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_194),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_200),
.B1(n_198),
.B2(n_194),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);


endmodule