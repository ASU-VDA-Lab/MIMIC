module fake_netlist_5_1901_n_4303 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_441, n_450, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4303);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_441;
input n_450;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4303;

wire n_924;
wire n_1263;
wire n_3304;
wire n_1378;
wire n_2417;
wire n_2253;
wire n_977;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_3241;
wire n_4129;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_3906;
wire n_4127;
wire n_880;
wire n_4138;
wire n_3297;
wire n_3086;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_4109;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3039;
wire n_3019;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_556;
wire n_2076;
wire n_2482;
wire n_3036;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1705;
wire n_659;
wire n_1294;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3834;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_2091;
wire n_1517;
wire n_2652;
wire n_2635;
wire n_2466;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3868;
wire n_3437;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_4187;
wire n_3089;
wire n_475;
wire n_1070;
wire n_1547;
wire n_777;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_521;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_1587;
wire n_680;
wire n_1473;
wire n_2682;
wire n_901;
wire n_553;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3542;
wire n_1167;
wire n_1626;
wire n_3436;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_3191;
wire n_571;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_3837;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_3593;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_3096;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_1002;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_593;
wire n_3487;
wire n_2258;
wire n_4069;
wire n_748;
wire n_1058;
wire n_1667;
wire n_586;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_647;
wire n_3433;
wire n_4024;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_561;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_4151;
wire n_4148;
wire n_1906;
wire n_1883;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3649;
wire n_3528;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4160;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_558;
wire n_3655;
wire n_2808;
wire n_702;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_809;
wire n_3923;
wire n_931;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_870;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_1888;
wire n_2009;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_843;
wire n_2491;
wire n_3747;
wire n_523;
wire n_1537;
wire n_913;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_776;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_498;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3113;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_568;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_3426;
wire n_3820;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3454;
wire n_636;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_2029;
wire n_742;
wire n_995;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_4232;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_974;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_761;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_512;
wire n_1591;
wire n_2033;
wire n_4071;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3077;
wire n_3929;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_860;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_495;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3824;
wire n_2662;
wire n_2740;
wire n_3751;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_4102;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_950;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_3033;
wire n_2824;
wire n_2650;
wire n_3298;
wire n_912;
wire n_968;
wire n_3548;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_483;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_762;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3632;
wire n_1966;
wire n_3231;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3482;
wire n_3417;
wire n_3866;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_918;
wire n_3854;
wire n_3529;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_4043;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2793;
wire n_2751;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_3869;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_4004;
wire n_4118;
wire n_2962;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3460;
wire n_3409;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_3697;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_487;
wire n_1726;
wire n_1584;
wire n_1835;
wire n_665;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_500;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_766;
wire n_1457;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3661;
wire n_3536;
wire n_3635;
wire n_4150;
wire n_827;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_3934;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_703;
wire n_698;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_737;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2774;
wire n_570;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_622;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_1567;
wire n_682;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3265;
wire n_3050;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_479;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_598;
wire n_685;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_499;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_722;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_1028;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_502;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_4061;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_3250;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3921;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_3772;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_4032;
wire n_2892;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_4212;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_491;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4245;
wire n_4288;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4222;
wire n_4216;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_3225;
wire n_1558;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_927;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_7),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_133),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_158),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_303),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_259),
.Y(n_480)
);

BUFx5_ASAP7_75t_L g481 ( 
.A(n_474),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_81),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_412),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_150),
.Y(n_484)
);

BUFx8_ASAP7_75t_SL g485 ( 
.A(n_106),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_340),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_234),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_261),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_271),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_228),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_366),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_63),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_360),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_271),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_239),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_84),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_135),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_144),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_186),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_280),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_24),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_20),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_276),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_329),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_263),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_228),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_387),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_130),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_40),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_378),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_303),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_467),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_32),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_344),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_11),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_190),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_198),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_40),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_1),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_135),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_339),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_218),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_440),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_379),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_151),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_222),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_184),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_112),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_26),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_306),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_162),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_173),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_232),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_98),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_279),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_417),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_416),
.Y(n_541)
);

CKINVDCx12_ASAP7_75t_R g542 ( 
.A(n_328),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_210),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_425),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_410),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_341),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_308),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_30),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_103),
.Y(n_549)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_1),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_435),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_5),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_294),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_151),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_459),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_403),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_134),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_222),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_372),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_344),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_199),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_347),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_269),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_83),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_144),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_468),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_57),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_114),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_49),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_422),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_145),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_101),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_22),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_117),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_466),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_206),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_212),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_111),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_207),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_330),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_108),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_71),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_373),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_460),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_400),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_170),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_322),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_227),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_99),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_266),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_206),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_332),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_112),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_223),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_274),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_145),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_378),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_186),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_436),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_82),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_201),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_333),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_184),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_193),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_28),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_9),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_193),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_183),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_366),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_148),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_295),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_95),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_204),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_103),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_411),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_259),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_2),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_92),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_249),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_67),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_354),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_20),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_245),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_53),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_394),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_94),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_443),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_446),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_24),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_310),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_224),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_248),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_342),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_125),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_63),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_230),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_153),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_83),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_181),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_207),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_202),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_118),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_62),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_0),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_354),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_242),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_35),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_239),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_377),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_176),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_247),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_143),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_462),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_313),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_95),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_11),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_53),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_295),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_342),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_152),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_210),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_290),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_57),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_240),
.Y(n_666)
);

BUFx8_ASAP7_75t_SL g667 ( 
.A(n_211),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_79),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_37),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_310),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_216),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_234),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_278),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_305),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_126),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_281),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_55),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_196),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_292),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_415),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_166),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_15),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_187),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_50),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_257),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_395),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_264),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_331),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_427),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_441),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_275),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_31),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_219),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_284),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_64),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_360),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_44),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_242),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_153),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_163),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_389),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_398),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_25),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_117),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_369),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_413),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_219),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_326),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_138),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_330),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_407),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_329),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_13),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_283),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_376),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_224),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_26),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_162),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_7),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_266),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_197),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_461),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_190),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_88),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_301),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_358),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_35),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_156),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_317),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_116),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_64),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_213),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_262),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_213),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_47),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_308),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_178),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_167),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_215),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_50),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_165),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_60),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_159),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_231),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_274),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_328),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_164),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_108),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_75),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_155),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_183),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_91),
.Y(n_752)
);

BUFx10_ASAP7_75t_L g753 ( 
.A(n_257),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_275),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_173),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_229),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_270),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_180),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_414),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_58),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_469),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_169),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_455),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_288),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_42),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_134),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_390),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_110),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_38),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_37),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_452),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_306),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_420),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_88),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_30),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_233),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_171),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_152),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_505),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_498),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_498),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_498),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_498),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_485),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_505),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_498),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_516),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_498),
.Y(n_788)
);

INVxp33_ASAP7_75t_L g789 ( 
.A(n_605),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_498),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_498),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_498),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_498),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_493),
.Y(n_794)
);

INVxp33_ASAP7_75t_SL g795 ( 
.A(n_605),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_493),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_493),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_653),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_493),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_493),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_493),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_485),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_493),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_543),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_543),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_543),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_543),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_761),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_653),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_761),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_543),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_543),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_543),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_542),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_521),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_773),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_521),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_492),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_475),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_521),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_583),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_667),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_583),
.Y(n_823)
);

BUFx2_ASAP7_75t_SL g824 ( 
.A(n_617),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_516),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_583),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_591),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_591),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_591),
.Y(n_829)
);

INVxp33_ASAP7_75t_SL g830 ( 
.A(n_492),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_592),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_592),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_592),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_667),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_560),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_642),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_642),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_642),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_541),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_663),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_663),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_560),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_663),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_694),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_694),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_694),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_718),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_718),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_544),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_718),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_730),
.Y(n_851)
);

INVxp33_ASAP7_75t_L g852 ( 
.A(n_687),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_730),
.Y(n_853)
);

INVxp33_ASAP7_75t_SL g854 ( 
.A(n_687),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_617),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_617),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_479),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_545),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_730),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_756),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_513),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_513),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_525),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_525),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_533),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_533),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_479),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_475),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_756),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_756),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_774),
.Y(n_871)
);

INVxp33_ASAP7_75t_L g872 ( 
.A(n_487),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_774),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_774),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_550),
.Y(n_875)
);

INVx4_ASAP7_75t_R g876 ( 
.A(n_483),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_479),
.Y(n_877)
);

INVxp33_ASAP7_75t_SL g878 ( 
.A(n_476),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_490),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_551),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_550),
.B(n_0),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_490),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_490),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_510),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_510),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_555),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_510),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_538),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_538),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_538),
.Y(n_890)
);

INVxp33_ASAP7_75t_SL g891 ( 
.A(n_477),
.Y(n_891)
);

CKINVDCx14_ASAP7_75t_R g892 ( 
.A(n_691),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_558),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_558),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_478),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_556),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_558),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_561),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_508),
.B(n_540),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_542),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_566),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_561),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_561),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_594),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_594),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_594),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_595),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_595),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_595),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_716),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_508),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_584),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_716),
.Y(n_913)
);

INVxp33_ASAP7_75t_SL g914 ( 
.A(n_482),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_716),
.Y(n_915)
);

CKINVDCx14_ASAP7_75t_R g916 ( 
.A(n_691),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_731),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_508),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_534),
.B(n_2),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_517),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_517),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_731),
.Y(n_922)
);

INVxp33_ASAP7_75t_SL g923 ( 
.A(n_484),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_731),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_764),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_764),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_779),
.A2(n_559),
.B1(n_613),
.B2(n_520),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_899),
.A2(n_759),
.B(n_540),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_794),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_920),
.B(n_856),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_808),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_855),
.B(n_480),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_784),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_780),
.A2(n_759),
.B(n_540),
.Y(n_935)
);

OAI22x1_ASAP7_75t_L g936 ( 
.A1(n_787),
.A2(n_825),
.B1(n_798),
.B2(n_733),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_877),
.B(n_480),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_808),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_808),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_809),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_861),
.B(n_759),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_877),
.B(n_480),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_794),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_796),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_814),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_808),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_875),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

OA21x2_ASAP7_75t_L g950 ( 
.A1(n_911),
.A2(n_570),
.B(n_534),
.Y(n_950)
);

BUFx12f_ASAP7_75t_L g951 ( 
.A(n_802),
.Y(n_951)
);

XNOR2xp5_ASAP7_75t_L g952 ( 
.A(n_830),
.B(n_661),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_796),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_810),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_810),
.Y(n_955)
);

INVx6_ASAP7_75t_L g956 ( 
.A(n_810),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_780),
.A2(n_575),
.B(n_570),
.Y(n_957)
);

BUFx8_ASAP7_75t_L g958 ( 
.A(n_895),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_862),
.B(n_575),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_881),
.B(n_690),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_797),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_895),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_797),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_799),
.Y(n_964)
);

OA21x2_ASAP7_75t_L g965 ( 
.A1(n_911),
.A2(n_589),
.B(n_585),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_799),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_800),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_800),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_819),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_868),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_856),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_801),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_879),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_839),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_918),
.A2(n_803),
.B(n_801),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_918),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_810),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_803),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_781),
.A2(n_589),
.B(n_585),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_559),
.B1(n_613),
.B2(n_520),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_921),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_804),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_863),
.B(n_600),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_879),
.B(n_766),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_804),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_805),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_864),
.B(n_600),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_892),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_805),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_806),
.Y(n_990)
);

INVx5_ASAP7_75t_L g991 ( 
.A(n_821),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_816),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_900),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_916),
.Y(n_994)
);

CKINVDCx6p67_ASAP7_75t_R g995 ( 
.A(n_901),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_781),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_806),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_821),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_835),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_782),
.A2(n_771),
.B(n_627),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_807),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_807),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_811),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_811),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_824),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_849),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_812),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_858),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_812),
.Y(n_1009)
);

AOI22x1_ASAP7_75t_SL g1010 ( 
.A1(n_822),
.A2(n_661),
.B1(n_664),
.B2(n_569),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_865),
.B(n_616),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_813),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_L g1013 ( 
.A(n_834),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_842),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_866),
.B(n_616),
.Y(n_1015)
);

INVxp33_ASAP7_75t_SL g1016 ( 
.A(n_880),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_813),
.B(n_627),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_823),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_789),
.A2(n_664),
.B1(n_713),
.B2(n_569),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_886),
.Y(n_1020)
);

BUFx12f_ASAP7_75t_L g1021 ( 
.A(n_896),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_823),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_782),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_831),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_783),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_882),
.B(n_511),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_831),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_840),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_912),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_840),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_882),
.B(n_511),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_869),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_878),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_869),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_857),
.B(n_867),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_883),
.Y(n_1036)
);

AOI22x1_ASAP7_75t_SL g1037 ( 
.A1(n_887),
.A2(n_713),
.B1(n_650),
.B2(n_671),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_783),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_786),
.Y(n_1039)
);

BUFx8_ASAP7_75t_SL g1040 ( 
.A(n_854),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_786),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_924),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_788),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_883),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_884),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_788),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_790),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_790),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_884),
.B(n_511),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_791),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_791),
.Y(n_1051)
);

CKINVDCx6p67_ASAP7_75t_R g1052 ( 
.A(n_824),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1035),
.B(n_885),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_999),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_974),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_939),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_975),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_1006),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_1008),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1035),
.B(n_885),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_1038),
.B(n_792),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1024),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_975),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_1016),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_975),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_939),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_975),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_932),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_976),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_932),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1005),
.B(n_960),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_976),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_992),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_995),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1039),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_969),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_969),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_1020),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1039),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_932),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_960),
.B(n_891),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1024),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1035),
.B(n_914),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1045),
.B(n_888),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_1020),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_970),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_1020),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1041),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1041),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1051),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1024),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1051),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1023),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_970),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_996),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_939),
.Y(n_1097)
);

OA21x2_ASAP7_75t_L g1098 ( 
.A1(n_935),
.A2(n_793),
.B(n_792),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1005),
.B(n_923),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1038),
.B(n_793),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_981),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_962),
.B(n_795),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1038),
.B(n_483),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1023),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_959),
.B(n_629),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1024),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1045),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_R g1108 ( 
.A(n_981),
.B(n_876),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_948),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1023),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_939),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1025),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_999),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1025),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1021),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1025),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_939),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_931),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1045),
.B(n_973),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1024),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1024),
.Y(n_1121)
);

AND2x6_ASAP7_75t_L g1122 ( 
.A(n_1017),
.B(n_761),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_931),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1038),
.B(n_690),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1034),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_996),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1034),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_959),
.B(n_629),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_L g1129 ( 
.A(n_1047),
.B(n_630),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1021),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1043),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_973),
.B(n_888),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1021),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1034),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_932),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1029),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1042),
.B(n_818),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_950),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_950),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_1014),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_950),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_995),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_950),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1034),
.Y(n_1145)
);

AND3x1_ASAP7_75t_L g1146 ( 
.A(n_1014),
.B(n_919),
.C(n_489),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1029),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_950),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1029),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1033),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_965),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_935),
.A2(n_817),
.B(n_815),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_965),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1040),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_988),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_941),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_988),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_965),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1034),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_965),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1047),
.B(n_889),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_988),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_988),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_994),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_965),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1043),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_994),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_994),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_932),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_994),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_932),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1043),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1034),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_935),
.A2(n_979),
.B(n_957),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1047),
.B(n_889),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1043),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_938),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_993),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_934),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1052),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_934),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_938),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_944),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_934),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_951),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_951),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_951),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1050),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_938),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1013),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_944),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1052),
.B(n_1013),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_944),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_939),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1050),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1013),
.Y(n_1196)
);

AND3x2_ASAP7_75t_L g1197 ( 
.A(n_962),
.B(n_757),
.C(n_733),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1047),
.B(n_890),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_945),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1050),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_939),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1050),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_973),
.B(n_893),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_958),
.B(n_852),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1017),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_959),
.B(n_701),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_938),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_930),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_993),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_958),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_996),
.B(n_893),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_930),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_953),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_953),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_963),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1036),
.B(n_894),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_R g1217 ( 
.A(n_958),
.B(n_655),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_941),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_963),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_959),
.B(n_701),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_945),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_938),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_996),
.B(n_894),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_958),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_967),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_948),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_936),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_971),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_967),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1036),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_972),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_945),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_961),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_961),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_961),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_971),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_964),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_971),
.Y(n_1238)
);

BUFx8_ASAP7_75t_L g1239 ( 
.A(n_983),
.Y(n_1239)
);

XNOR2xp5_ASAP7_75t_L g1240 ( 
.A(n_1019),
.B(n_571),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_971),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_952),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_952),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_946),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_996),
.B(n_897),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_938),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_955),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1019),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_972),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1010),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1010),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_946),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_955),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_978),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_936),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_978),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_936),
.Y(n_1257)
);

XOR2xp5_ASAP7_75t_L g1258 ( 
.A(n_1037),
.B(n_674),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_980),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_989),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_989),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_980),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1037),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_996),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_996),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1046),
.Y(n_1266)
);

NAND2xp33_ASAP7_75t_SL g1267 ( 
.A(n_928),
.B(n_519),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_964),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_933),
.B(n_872),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_955),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_928),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1046),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_983),
.B(n_771),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_933),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1044),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1082),
.B(n_680),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1269),
.B(n_983),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1076),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1192),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1205),
.Y(n_1280)
);

BUFx8_ASAP7_75t_SL g1281 ( 
.A(n_1154),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1275),
.B(n_1026),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1076),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1080),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1080),
.Y(n_1285)
);

NOR3xp33_ASAP7_75t_L g1286 ( 
.A(n_1072),
.B(n_598),
.C(n_757),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1152),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1119),
.B(n_1046),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1085),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1077),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1057),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1084),
.B(n_1026),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1152),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1152),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1205),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1085),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1053),
.B(n_983),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1108),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1089),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1089),
.Y(n_1300)
);

BUFx10_ASAP7_75t_L g1301 ( 
.A(n_1099),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1057),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1090),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1058),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1062),
.A2(n_929),
.B(n_957),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1152),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1098),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1259),
.A2(n_1011),
.B1(n_1015),
.B2(n_987),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1118),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1156),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1107),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1053),
.A2(n_1061),
.B(n_1216),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1138),
.B(n_580),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1058),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1064),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1105),
.A2(n_929),
.B1(n_1017),
.B2(n_1011),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1090),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1091),
.Y(n_1318)
);

INVx8_ASAP7_75t_L g1319 ( 
.A(n_1122),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1064),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1091),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1065),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1055),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1096),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1066),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1066),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1118),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1123),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1123),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1093),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1227),
.A2(n_669),
.B1(n_672),
.B2(n_580),
.Y(n_1331)
);

INVx4_ASAP7_75t_SL g1332 ( 
.A(n_1122),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1068),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1093),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1068),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1208),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1098),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1208),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1212),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1139),
.A2(n_979),
.B(n_957),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_SL g1341 ( 
.A(n_1131),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1107),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1212),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1119),
.B(n_1046),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1262),
.A2(n_1011),
.B1(n_1015),
.B2(n_987),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1070),
.B(n_1046),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1213),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1131),
.B(n_686),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1098),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1213),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1214),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1180),
.B(n_689),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1214),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1215),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1275),
.B(n_937),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1109),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1215),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_1218),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1219),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1219),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1105),
.A2(n_929),
.B1(n_1017),
.B2(n_1011),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_1209),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1225),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1105),
.A2(n_929),
.B1(n_1015),
.B2(n_987),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1225),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1229),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1098),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1229),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1069),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1070),
.B(n_1046),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1054),
.B(n_1113),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1231),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1249),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1141),
.B(n_669),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1249),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1254),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1180),
.B(n_1061),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1105),
.B(n_987),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1087),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1139),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1103),
.B(n_929),
.C(n_1015),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1178),
.B(n_672),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1254),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1218),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1133),
.B(n_937),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1256),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1073),
.B(n_1046),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1073),
.B(n_1132),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1124),
.B(n_998),
.Y(n_1390)
);

INVx8_ASAP7_75t_L g1391 ( 
.A(n_1122),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1256),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1062),
.A2(n_1000),
.B(n_979),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1140),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1069),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1244),
.B(n_678),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1260),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1128),
.B(n_942),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1140),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1261),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1261),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1133),
.B(n_943),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1161),
.B(n_1198),
.C(n_1175),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1244),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1142),
.B(n_998),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1166),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1166),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1274),
.B(n_678),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1255),
.B(n_702),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1102),
.B(n_684),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1142),
.B(n_998),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1144),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1239),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1069),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1172),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1144),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1148),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1203),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1148),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1151),
.B(n_998),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1151),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1153),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1153),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1257),
.B(n_706),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1059),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1158),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1217),
.B(n_711),
.Y(n_1428)
);

AND2x6_ASAP7_75t_L g1429 ( 
.A(n_1158),
.B(n_761),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1239),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1172),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1216),
.B(n_722),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1160),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1230),
.B(n_684),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1160),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1203),
.B(n_984),
.C(n_943),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1176),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1165),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1165),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1176),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1183),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1188),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1128),
.B(n_942),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1188),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1100),
.B(n_942),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1195),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1183),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1191),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1191),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1195),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_SL g1451 ( 
.A(n_1128),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1078),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1069),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1200),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1239),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1193),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1128),
.B(n_984),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1056),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1096),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1227),
.A2(n_700),
.B1(n_598),
.B2(n_523),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1206),
.B(n_1220),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1200),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1193),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1202),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1199),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1096),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1146),
.A2(n_1267),
.B1(n_1220),
.B2(n_1206),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1206),
.A2(n_1000),
.B1(n_942),
.B2(n_761),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1096),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1199),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_SL g1471 ( 
.A(n_1206),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1221),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1221),
.Y(n_1473)
);

BUFx10_ASAP7_75t_L g1474 ( 
.A(n_1150),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1232),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1202),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1220),
.A2(n_1000),
.B1(n_761),
.B2(n_523),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1220),
.B(n_763),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1060),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1211),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1223),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1273),
.B(n_1048),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1095),
.B(n_700),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1069),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1273),
.A2(n_750),
.B1(n_755),
.B2(n_732),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1101),
.B(n_486),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1232),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1245),
.Y(n_1488)
);

INVx5_ASAP7_75t_L g1489 ( 
.A(n_1122),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1094),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1197),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1273),
.B(n_1031),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_1240),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1094),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1233),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1233),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1252),
.B(n_488),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1074),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1273),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_SL g1500 ( 
.A(n_1170),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1056),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1063),
.B(n_898),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1271),
.B(n_491),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1204),
.B(n_1031),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1248),
.B(n_1049),
.C(n_496),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1056),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1234),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1104),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1079),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1075),
.Y(n_1510)
);

NAND2xp33_ASAP7_75t_R g1511 ( 
.A(n_1242),
.B(n_767),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1226),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1126),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1109),
.B(n_495),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1174),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1240),
.Y(n_1516)
);

AND2x6_ASAP7_75t_L g1517 ( 
.A(n_1264),
.B(n_761),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1104),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1234),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1235),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1380),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1302),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1302),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1302),
.Y(n_1524)
);

AO221x1_ASAP7_75t_L g1525 ( 
.A1(n_1331),
.A2(n_489),
.B1(n_497),
.B2(n_494),
.C(n_487),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1313),
.B(n_1210),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1407),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1292),
.B(n_1224),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1407),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1295),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1342),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1277),
.B(n_1129),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1302),
.B(n_1239),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1358),
.B(n_1228),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1386),
.B(n_1264),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1358),
.B(n_1236),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1302),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1397),
.B(n_1238),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1408),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_L g1540 ( 
.A(n_1461),
.B(n_1241),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1408),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1372),
.B(n_1385),
.Y(n_1542)
);

AND2x6_ASAP7_75t_L g1543 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1323),
.B(n_1086),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1304),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_SL g1546 ( 
.A(n_1474),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1414),
.B(n_519),
.Y(n_1547)
);

BUFx8_ASAP7_75t_L g1548 ( 
.A(n_1500),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1419),
.B(n_1088),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1416),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1411),
.B(n_1130),
.C(n_1115),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1416),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1405),
.B(n_1134),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1386),
.B(n_1265),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1419),
.B(n_1137),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1312),
.B(n_1149),
.Y(n_1556)
);

NOR2xp67_ASAP7_75t_L g1557 ( 
.A(n_1279),
.B(n_1147),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1503),
.B(n_1265),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1290),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1304),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1403),
.B(n_1266),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1304),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1355),
.B(n_1266),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1431),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1312),
.B(n_1157),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1304),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1375),
.B(n_1179),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1310),
.B(n_1181),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1304),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1325),
.B(n_1272),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1355),
.B(n_1155),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1309),
.B(n_1162),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1309),
.B(n_1163),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1457),
.B(n_1110),
.Y(n_1574)
);

INVxp33_ASAP7_75t_L g1575 ( 
.A(n_1409),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1325),
.B(n_1126),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1325),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1325),
.B(n_1126),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1457),
.A2(n_1122),
.B1(n_1112),
.B2(n_1114),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1437),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1308),
.A2(n_1112),
.B(n_1114),
.C(n_1110),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1289),
.B(n_1116),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1289),
.B(n_1296),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1325),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1437),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1296),
.B(n_1116),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1297),
.B(n_1056),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1295),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_L g1589 ( 
.A(n_1461),
.B(n_1164),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1369),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1338),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1295),
.B(n_1167),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1297),
.B(n_1067),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1327),
.B(n_1168),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1327),
.B(n_1184),
.Y(n_1595)
);

INVxp33_ASAP7_75t_SL g1596 ( 
.A(n_1323),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1328),
.B(n_1185),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1291),
.B(n_1067),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1280),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1278),
.B(n_1067),
.Y(n_1600)
);

NOR3xp33_ASAP7_75t_L g1601 ( 
.A(n_1497),
.B(n_1263),
.C(n_1187),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1278),
.B(n_1067),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1383),
.B(n_1186),
.Y(n_1603)
);

BUFx8_ASAP7_75t_L g1604 ( 
.A(n_1500),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1283),
.B(n_1097),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1369),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1440),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1338),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1329),
.B(n_1190),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1283),
.B(n_1097),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1284),
.B(n_1097),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_L g1612 ( 
.A(n_1279),
.B(n_1196),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1440),
.Y(n_1613)
);

BUFx5_ASAP7_75t_L g1614 ( 
.A(n_1461),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1434),
.B(n_898),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1284),
.B(n_1097),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1285),
.B(n_1111),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1329),
.B(n_1126),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1282),
.B(n_1111),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1442),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1489),
.B(n_1063),
.Y(n_1621)
);

NOR3xp33_ASAP7_75t_L g1622 ( 
.A(n_1514),
.B(n_1251),
.C(n_1250),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1282),
.B(n_1111),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1285),
.B(n_1111),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1299),
.B(n_1117),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1442),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1280),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1299),
.B(n_1117),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_L g1629 ( 
.A(n_1356),
.B(n_903),
.C(n_902),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1399),
.A2(n_1122),
.B1(n_1174),
.B2(n_1092),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1339),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1300),
.B(n_1117),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1505),
.B(n_1117),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1489),
.B(n_1083),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1300),
.B(n_1194),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1426),
.B(n_902),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1303),
.B(n_1194),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1489),
.B(n_1083),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1303),
.B(n_1194),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1311),
.B(n_1092),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1444),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1317),
.B(n_1194),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1339),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1489),
.B(n_1106),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1369),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1343),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1317),
.B(n_1201),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1318),
.B(n_1201),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1467),
.B(n_1071),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_L g1650 ( 
.A(n_1461),
.B(n_1122),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1318),
.B(n_1321),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1378),
.B(n_1201),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1414),
.B(n_519),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1483),
.Y(n_1654)
);

BUFx5_ASAP7_75t_L g1655 ( 
.A(n_1461),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1321),
.B(n_1201),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1330),
.B(n_1270),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1452),
.B(n_1207),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1343),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1362),
.B(n_1207),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1350),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_SL g1662 ( 
.A(n_1474),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1356),
.B(n_904),
.C(n_903),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1350),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1444),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1446),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1489),
.B(n_1106),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1467),
.B(n_1280),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_SL g1670 ( 
.A(n_1474),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1354),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1446),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1334),
.B(n_1270),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1450),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1308),
.B(n_1345),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1354),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1336),
.B(n_1347),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1345),
.B(n_1207),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1486),
.B(n_503),
.C(n_501),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1450),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1516),
.B(n_905),
.C(n_904),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1281),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1286),
.B(n_507),
.C(n_504),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_L g1684 ( 
.A(n_1461),
.B(n_481),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1454),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1336),
.B(n_1270),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1347),
.B(n_1270),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1512),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1351),
.B(n_1120),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1351),
.B(n_1120),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1454),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1512),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1462),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1462),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1489),
.B(n_1121),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1511),
.B(n_515),
.C(n_514),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1491),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_L g1698 ( 
.A(n_1461),
.B(n_481),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1499),
.B(n_1121),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1342),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1499),
.B(n_1125),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_L g1702 ( 
.A(n_1342),
.B(n_481),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1301),
.B(n_905),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1353),
.B(n_1125),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1464),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1464),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1379),
.B(n_1127),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1491),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1365),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1353),
.B(n_1127),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1379),
.B(n_1413),
.Y(n_1711)
);

XNOR2x2_ASAP7_75t_L g1712 ( 
.A(n_1485),
.B(n_1258),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1357),
.B(n_1135),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1365),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1342),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_L g1716 ( 
.A(n_1342),
.B(n_481),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1357),
.B(n_1135),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1436),
.B(n_1485),
.Y(n_1718)
);

BUFx8_ASAP7_75t_L g1719 ( 
.A(n_1500),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1379),
.B(n_1071),
.Y(n_1720)
);

AND2x6_ASAP7_75t_SL g1721 ( 
.A(n_1504),
.B(n_494),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1314),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1410),
.B(n_907),
.C(n_906),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1311),
.B(n_1379),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1413),
.B(n_1145),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1359),
.B(n_1145),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1436),
.B(n_522),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1276),
.B(n_524),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1366),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1399),
.B(n_1071),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1359),
.B(n_1159),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1366),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1399),
.B(n_1071),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1301),
.B(n_906),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1371),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1476),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_L g1737 ( 
.A(n_1319),
.B(n_481),
.Y(n_1737)
);

INVxp33_ASAP7_75t_L g1738 ( 
.A(n_1425),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1476),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1301),
.B(n_907),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1371),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1504),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1369),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1360),
.B(n_1159),
.Y(n_1744)
);

AO221x1_ASAP7_75t_L g1745 ( 
.A1(n_1460),
.A2(n_499),
.B1(n_502),
.B2(n_500),
.C(n_497),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1373),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1479),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1373),
.Y(n_1748)
);

BUFx5_ASAP7_75t_L g1749 ( 
.A(n_1429),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1360),
.B(n_1173),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1417),
.B(n_1173),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1363),
.B(n_1235),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1363),
.B(n_1237),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1368),
.B(n_1237),
.Y(n_1754)
);

AO221x1_ASAP7_75t_L g1755 ( 
.A1(n_1368),
.A2(n_500),
.B1(n_506),
.B2(n_502),
.C(n_499),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1374),
.B(n_530),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1376),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1376),
.Y(n_1758)
);

AND2x2_ASAP7_75t_SL g1759 ( 
.A(n_1477),
.B(n_1174),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1417),
.B(n_1071),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1591),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1559),
.Y(n_1762)
);

AO22x2_ASAP7_75t_L g1763 ( 
.A1(n_1712),
.A2(n_1258),
.B1(n_681),
.B2(n_564),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1591),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1718),
.A2(n_1493),
.B1(n_1432),
.B2(n_1504),
.C(n_1298),
.Y(n_1765)
);

AO22x2_ASAP7_75t_L g1766 ( 
.A1(n_1669),
.A2(n_681),
.B1(n_564),
.B2(n_532),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1608),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1608),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1631),
.Y(n_1769)
);

AO22x2_ASAP7_75t_L g1770 ( 
.A1(n_1675),
.A2(n_681),
.B1(n_564),
.B2(n_532),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1631),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1558),
.B(n_1389),
.Y(n_1772)
);

BUFx8_ASAP7_75t_L g1773 ( 
.A(n_1546),
.Y(n_1773)
);

AO22x2_ASAP7_75t_L g1774 ( 
.A1(n_1675),
.A2(n_766),
.B1(n_532),
.B2(n_603),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1643),
.Y(n_1775)
);

AO22x2_ASAP7_75t_L g1776 ( 
.A1(n_1654),
.A2(n_603),
.B1(n_693),
.B2(n_523),
.Y(n_1776)
);

AO22x2_ASAP7_75t_L g1777 ( 
.A1(n_1533),
.A2(n_693),
.B1(n_714),
.B2(n_603),
.Y(n_1777)
);

AO22x2_ASAP7_75t_L g1778 ( 
.A1(n_1533),
.A2(n_714),
.B1(n_738),
.B2(n_693),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1521),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1643),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1575),
.B(n_1479),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1558),
.B(n_1374),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1724),
.B(n_1455),
.Y(n_1783)
);

NOR2xp67_ASAP7_75t_L g1784 ( 
.A(n_1747),
.B(n_1498),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1566),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1563),
.B(n_1377),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1724),
.B(n_1455),
.Y(n_1787)
);

AO22x2_ASAP7_75t_L g1788 ( 
.A1(n_1649),
.A2(n_738),
.B1(n_766),
.B2(n_714),
.Y(n_1788)
);

OAI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1526),
.A2(n_1504),
.B1(n_1352),
.B2(n_1348),
.C(n_1498),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1528),
.A2(n_1471),
.B1(n_1451),
.B2(n_1492),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1527),
.Y(n_1791)
);

AO22x2_ASAP7_75t_L g1792 ( 
.A1(n_1721),
.A2(n_1703),
.B1(n_1740),
.B2(n_1734),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1724),
.B(n_1430),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1542),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1530),
.B(n_1430),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1615),
.B(n_1301),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1567),
.B(n_1474),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1563),
.B(n_1377),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1603),
.B(n_1322),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1529),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1646),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1539),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1619),
.B(n_1384),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1541),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1646),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1659),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1550),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1552),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1659),
.Y(n_1809)
);

AO22x2_ASAP7_75t_L g1810 ( 
.A1(n_1565),
.A2(n_1692),
.B1(n_1564),
.B2(n_1580),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1585),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1661),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1661),
.Y(n_1813)
);

AO22x2_ASAP7_75t_L g1814 ( 
.A1(n_1607),
.A2(n_738),
.B1(n_1387),
.B2(n_1384),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1613),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1620),
.Y(n_1816)
);

AO22x2_ASAP7_75t_L g1817 ( 
.A1(n_1626),
.A2(n_1392),
.B1(n_1393),
.B2(n_1387),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1528),
.A2(n_1471),
.B1(n_1451),
.B2(n_1492),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1688),
.B(n_1542),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1641),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1664),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1619),
.B(n_1392),
.Y(n_1822)
);

AO22x2_ASAP7_75t_L g1823 ( 
.A1(n_1666),
.A2(n_1398),
.B1(n_1393),
.B2(n_509),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1697),
.B(n_1399),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1568),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1623),
.B(n_1398),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1547),
.B(n_1492),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1623),
.B(n_1401),
.Y(n_1828)
);

AO22x2_ASAP7_75t_L g1829 ( 
.A1(n_1667),
.A2(n_509),
.B1(n_512),
.B2(n_506),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_SL g1830 ( 
.A(n_1547),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1722),
.B(n_1401),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1672),
.Y(n_1832)
);

OR2x6_ASAP7_75t_SL g1833 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1531),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1538),
.B(n_1322),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1664),
.Y(n_1836)
);

AO22x2_ASAP7_75t_L g1837 ( 
.A1(n_1674),
.A2(n_518),
.B1(n_526),
.B2(n_512),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1680),
.A2(n_526),
.B1(n_527),
.B2(n_518),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_L g1839 ( 
.A(n_1614),
.B(n_1319),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1756),
.B(n_1402),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1526),
.B(n_1322),
.Y(n_1841)
);

OAI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1681),
.A2(n_1728),
.B1(n_1663),
.B2(n_1629),
.C(n_1696),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1685),
.A2(n_528),
.B1(n_529),
.B2(n_527),
.Y(n_1843)
);

AO22x2_ASAP7_75t_L g1844 ( 
.A1(n_1691),
.A2(n_529),
.B1(n_537),
.B2(n_528),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1708),
.B(n_1443),
.Y(n_1845)
);

AO22x2_ASAP7_75t_L g1846 ( 
.A1(n_1693),
.A2(n_546),
.B1(n_552),
.B2(n_537),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1595),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1694),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1595),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1705),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1706),
.Y(n_1851)
);

NAND2x1_ASAP7_75t_L g1852 ( 
.A(n_1566),
.B(n_1324),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1756),
.B(n_1402),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1728),
.A2(n_1471),
.B1(n_1451),
.B2(n_1492),
.Y(n_1854)
);

NAND2x1p5_ASAP7_75t_L g1855 ( 
.A(n_1530),
.B(n_1443),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1856)
);

AO22x2_ASAP7_75t_L g1857 ( 
.A1(n_1736),
.A2(n_552),
.B1(n_562),
.B2(n_546),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1727),
.A2(n_1492),
.B1(n_1443),
.B2(n_1478),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1739),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1671),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1571),
.A2(n_1428),
.B1(n_535),
.B2(n_539),
.C(n_536),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1554),
.B(n_1480),
.Y(n_1863)
);

OAI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1727),
.A2(n_547),
.B1(n_549),
.B2(n_548),
.C(n_531),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1671),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1676),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1676),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1640),
.B(n_1443),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1597),
.Y(n_1869)
);

AO22x2_ASAP7_75t_L g1870 ( 
.A1(n_1556),
.A2(n_572),
.B1(n_573),
.B2(n_562),
.Y(n_1870)
);

AO22x2_ASAP7_75t_L g1871 ( 
.A1(n_1622),
.A2(n_1665),
.B1(n_1677),
.B2(n_1651),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1709),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1561),
.B(n_1480),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1596),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1640),
.B(n_1502),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1640),
.B(n_1502),
.Y(n_1876)
);

BUFx8_ASAP7_75t_L g1877 ( 
.A(n_1546),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1709),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1714),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1714),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1729),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1729),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1732),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1732),
.Y(n_1884)
);

AO22x2_ASAP7_75t_L g1885 ( 
.A1(n_1683),
.A2(n_573),
.B1(n_577),
.B2(n_572),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1735),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1735),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1746),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1682),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1534),
.A2(n_554),
.B1(n_563),
.B2(n_557),
.C(n_553),
.Y(n_1890)
);

CKINVDCx16_ASAP7_75t_R g1891 ( 
.A(n_1544),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1746),
.Y(n_1892)
);

AO22x2_ASAP7_75t_L g1893 ( 
.A1(n_1601),
.A2(n_578),
.B1(n_581),
.B2(n_577),
.Y(n_1893)
);

BUFx8_ASAP7_75t_L g1894 ( 
.A(n_1662),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1547),
.B(n_1319),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1757),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1574),
.B(n_1481),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1738),
.B(n_1243),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1757),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1636),
.B(n_1534),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1618),
.B(n_1488),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1566),
.B(n_1324),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1543),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1543),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1742),
.A2(n_1678),
.B1(n_1679),
.B2(n_1633),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1678),
.A2(n_1341),
.B1(n_1488),
.B2(n_1502),
.Y(n_1906)
);

OAI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1536),
.A2(n_567),
.B1(n_574),
.B2(n_568),
.C(n_565),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1543),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1543),
.Y(n_1909)
);

AND2x6_ASAP7_75t_L g1910 ( 
.A(n_1522),
.B(n_1314),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1536),
.B(n_1502),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1741),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1592),
.B(n_1332),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1711),
.A2(n_1429),
.B1(n_1404),
.B2(n_1445),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1609),
.B(n_908),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1543),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1553),
.B(n_1341),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1711),
.A2(n_1429),
.B1(n_1404),
.B2(n_1422),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1748),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1758),
.Y(n_1920)
);

AO22x2_ASAP7_75t_L g1921 ( 
.A1(n_1525),
.A2(n_581),
.B1(n_601),
.B2(n_578),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1630),
.A2(n_1364),
.B1(n_1361),
.B2(n_1316),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1599),
.Y(n_1923)
);

BUFx8_ASAP7_75t_L g1924 ( 
.A(n_1662),
.Y(n_1924)
);

AO22x2_ASAP7_75t_L g1925 ( 
.A1(n_1522),
.A2(n_604),
.B1(n_607),
.B2(n_601),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1653),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1553),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1572),
.Y(n_1928)
);

AO22x2_ASAP7_75t_L g1929 ( 
.A1(n_1523),
.A2(n_607),
.B1(n_610),
.B2(n_604),
.Y(n_1929)
);

AO22x2_ASAP7_75t_L g1930 ( 
.A1(n_1523),
.A2(n_615),
.B1(n_618),
.B2(n_610),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1531),
.B(n_1332),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1582),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1752),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1572),
.B(n_1341),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1599),
.Y(n_1935)
);

AO22x2_ASAP7_75t_L g1936 ( 
.A1(n_1524),
.A2(n_618),
.B1(n_621),
.B2(n_615),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1573),
.B(n_1510),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1573),
.B(n_908),
.Y(n_1938)
);

AO22x2_ASAP7_75t_L g1939 ( 
.A1(n_1524),
.A2(n_632),
.B1(n_636),
.B2(n_621),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1627),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1627),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1660),
.B(n_1406),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1670),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1594),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1586),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1588),
.B(n_1332),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1594),
.B(n_909),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1753),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1537),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1618),
.B(n_1315),
.Y(n_1950)
);

BUFx12f_ASAP7_75t_L g1951 ( 
.A(n_1548),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1759),
.B(n_1315),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1537),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1658),
.B(n_1143),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1653),
.Y(n_1955)
);

AO22x2_ASAP7_75t_L g1956 ( 
.A1(n_1545),
.A2(n_636),
.B1(n_643),
.B2(n_632),
.Y(n_1956)
);

BUFx8_ASAP7_75t_L g1957 ( 
.A(n_1670),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1754),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1759),
.B(n_1320),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1689),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1690),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1704),
.Y(n_1962)
);

OAI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1723),
.A2(n_579),
.B1(n_586),
.B2(n_582),
.C(n_576),
.Y(n_1963)
);

BUFx8_ASAP7_75t_L g1964 ( 
.A(n_1548),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1772),
.A2(n_1782),
.B1(n_1798),
.B2(n_1786),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1796),
.B(n_1658),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1791),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1932),
.B(n_1587),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1922),
.A2(n_1588),
.B1(n_1577),
.B2(n_1566),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1945),
.B(n_1593),
.Y(n_1970)
);

OAI21xp33_ASAP7_75t_L g1971 ( 
.A1(n_1864),
.A2(n_1555),
.B(n_1549),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1859),
.B(n_1532),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1800),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1761),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1927),
.B(n_1794),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1915),
.B(n_1320),
.Y(n_1976)
);

AO21x2_ASAP7_75t_L g1977 ( 
.A1(n_1901),
.A2(n_1581),
.B(n_1382),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1839),
.A2(n_1578),
.B(n_1576),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1781),
.A2(n_1557),
.B1(n_1612),
.B2(n_1589),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1905),
.A2(n_1382),
.B(n_1652),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_L g1981 ( 
.A(n_1784),
.B(n_1700),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1840),
.A2(n_1578),
.B(n_1576),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1853),
.A2(n_1459),
.B(n_1324),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1938),
.B(n_1947),
.Y(n_1984)
);

A2O1A1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1789),
.A2(n_1652),
.B(n_1698),
.C(n_1684),
.Y(n_1985)
);

OR2x6_ASAP7_75t_SL g1986 ( 
.A(n_1874),
.B(n_587),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1847),
.B(n_1653),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1842),
.A2(n_1579),
.B(n_1540),
.C(n_1650),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1802),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1775),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1897),
.B(n_1326),
.Y(n_1991)
);

O2A1O1Ixp33_ASAP7_75t_L g1992 ( 
.A1(n_1765),
.A2(n_1716),
.B(n_1702),
.C(n_1707),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1849),
.B(n_1700),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1869),
.B(n_1715),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1862),
.A2(n_1707),
.B(n_646),
.C(n_648),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1911),
.B(n_1326),
.Y(n_1996)
);

CKINVDCx10_ASAP7_75t_R g1997 ( 
.A(n_1830),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1900),
.B(n_1333),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1950),
.A2(n_1466),
.B(n_1459),
.Y(n_1999)
);

AO21x1_ASAP7_75t_L g2000 ( 
.A1(n_1803),
.A2(n_1713),
.B(n_1710),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1931),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1792),
.A2(n_1745),
.B1(n_1755),
.B2(n_1730),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1931),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1891),
.B(n_1577),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1783),
.B(n_1715),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1948),
.B(n_1333),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1801),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1858),
.A2(n_1390),
.B(n_1737),
.C(n_1726),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1863),
.A2(n_1466),
.B(n_1459),
.Y(n_2009)
);

NOR2xp67_ASAP7_75t_L g2010 ( 
.A(n_1762),
.B(n_1720),
.Y(n_2010)
);

BUFx12f_ASAP7_75t_L g2011 ( 
.A(n_1964),
.Y(n_2011)
);

AO32x2_ASAP7_75t_L g2012 ( 
.A1(n_1766),
.A2(n_1515),
.A3(n_1340),
.B1(n_1394),
.B2(n_1305),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1873),
.A2(n_1469),
.B(n_1466),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1906),
.A2(n_1560),
.B1(n_1562),
.B2(n_1545),
.Y(n_2014)
);

O2A1O1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1928),
.A2(n_1944),
.B(n_1890),
.C(n_1907),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1804),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1958),
.B(n_1335),
.Y(n_2017)
);

AO32x1_ASAP7_75t_L g2018 ( 
.A1(n_1912),
.A2(n_646),
.A3(n_651),
.B1(n_648),
.B2(n_643),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1933),
.B(n_1424),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1807),
.Y(n_2020)
);

AND2x6_ASAP7_75t_L g2021 ( 
.A(n_1903),
.B(n_1560),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1819),
.B(n_1604),
.Y(n_2022)
);

O2A1O1Ixp33_ASAP7_75t_SL g2023 ( 
.A1(n_1903),
.A2(n_1699),
.B(n_1701),
.C(n_1570),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1799),
.B(n_909),
.Y(n_2024)
);

A2O1A1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1934),
.A2(n_1731),
.B(n_1744),
.C(n_1717),
.Y(n_2025)
);

O2A1O1Ixp33_ASAP7_75t_L g2026 ( 
.A1(n_1963),
.A2(n_654),
.B(n_659),
.C(n_651),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1783),
.B(n_1733),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1933),
.B(n_1418),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1805),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1822),
.A2(n_1513),
.B(n_1469),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1960),
.B(n_1418),
.Y(n_2031)
);

A2O1A1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_1917),
.A2(n_1750),
.B(n_1569),
.C(n_1584),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1828),
.A2(n_1513),
.B(n_1469),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1808),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1797),
.B(n_910),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1856),
.B(n_1604),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1961),
.B(n_1433),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1787),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1962),
.A2(n_1569),
.B(n_1584),
.C(n_1562),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1826),
.A2(n_1513),
.B(n_1344),
.Y(n_2040)
);

BUFx4f_ASAP7_75t_L g2041 ( 
.A(n_1951),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1831),
.A2(n_1288),
.B(n_1468),
.Y(n_2042)
);

AO21x1_ASAP7_75t_L g2043 ( 
.A1(n_1904),
.A2(n_1701),
.B(n_1699),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1787),
.B(n_1590),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1914),
.A2(n_1370),
.B(n_1346),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1918),
.A2(n_1395),
.B(n_1381),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1962),
.B(n_1420),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1954),
.B(n_1719),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_SL g2049 ( 
.A(n_1889),
.B(n_1719),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1825),
.B(n_1570),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1952),
.A2(n_1395),
.B(n_1381),
.Y(n_2051)
);

INVx1_ASAP7_75t_SL g2052 ( 
.A(n_1779),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1841),
.B(n_1412),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1959),
.A2(n_1395),
.B(n_1381),
.Y(n_2054)
);

AO21x1_ASAP7_75t_L g2055 ( 
.A1(n_1904),
.A2(n_1909),
.B(n_1908),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1902),
.A2(n_1423),
.B(n_1400),
.Y(n_2056)
);

OAI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1942),
.A2(n_1388),
.B(n_1600),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1811),
.B(n_1433),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_SL g2059 ( 
.A(n_1955),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1835),
.B(n_1937),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1815),
.A2(n_659),
.B(n_662),
.C(n_654),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1816),
.B(n_1439),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1820),
.B(n_1832),
.Y(n_2063)
);

OAI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1919),
.A2(n_1656),
.B(n_1605),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1848),
.B(n_1439),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1946),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1871),
.A2(n_1423),
.B(n_1400),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1871),
.A2(n_1423),
.B(n_1400),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1850),
.B(n_1422),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1793),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1868),
.B(n_1824),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1817),
.A2(n_1515),
.B(n_1598),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1851),
.B(n_1424),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1852),
.A2(n_1396),
.B(n_1369),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1926),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1946),
.A2(n_1415),
.B(n_1396),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_1792),
.A2(n_1763),
.B1(n_1868),
.B2(n_1875),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1943),
.B(n_1614),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1860),
.B(n_1420),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_1875),
.A2(n_1415),
.B(n_1396),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1870),
.B(n_1435),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1763),
.B(n_910),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_1876),
.A2(n_1415),
.B(n_1396),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1806),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_1898),
.Y(n_2085)
);

OR2x6_ASAP7_75t_SL g2086 ( 
.A(n_1923),
.B(n_588),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1876),
.A2(n_1415),
.B(n_1396),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1855),
.A2(n_1453),
.B(n_1415),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1824),
.B(n_1614),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1870),
.B(n_1427),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1834),
.Y(n_2091)
);

INVxp67_ASAP7_75t_L g2092 ( 
.A(n_1833),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1809),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1949),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1817),
.A2(n_1484),
.B(n_1453),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1920),
.A2(n_1648),
.B(n_1610),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1845),
.B(n_1614),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1812),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1908),
.A2(n_1349),
.B(n_1427),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1854),
.A2(n_1484),
.B(n_1453),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_L g2101 ( 
.A(n_1795),
.B(n_1614),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1773),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1790),
.A2(n_1438),
.B1(n_1435),
.B2(n_1743),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_1909),
.A2(n_1349),
.B(n_1438),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1845),
.B(n_1823),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_1916),
.A2(n_1349),
.B(n_1421),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1861),
.A2(n_1611),
.B(n_1602),
.Y(n_2107)
);

O2A1O1Ixp33_ASAP7_75t_L g2108 ( 
.A1(n_1827),
.A2(n_665),
.B(n_670),
.C(n_662),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1823),
.B(n_1349),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1885),
.B(n_913),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1865),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1916),
.A2(n_1349),
.B(n_1616),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_1885),
.A2(n_1655),
.B1(n_478),
.B2(n_1429),
.Y(n_2113)
);

AND2x2_ASAP7_75t_SL g2114 ( 
.A(n_1818),
.B(n_1590),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1893),
.B(n_913),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1773),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1810),
.A2(n_1624),
.B(n_1617),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1810),
.A2(n_1628),
.B(n_1625),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1764),
.A2(n_1635),
.B(n_1632),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1813),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1814),
.B(n_1490),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1766),
.B(n_1494),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1821),
.Y(n_2123)
);

OAI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_1866),
.A2(n_1639),
.B(n_1637),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_1764),
.A2(n_1647),
.B(n_1642),
.Y(n_2125)
);

A2O1A1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_1935),
.A2(n_1673),
.B(n_1686),
.C(n_1657),
.Y(n_2126)
);

AO21x2_ASAP7_75t_L g2127 ( 
.A1(n_1767),
.A2(n_1760),
.B(n_1687),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1767),
.B(n_1494),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1768),
.B(n_1508),
.Y(n_2129)
);

AOI21x1_ASAP7_75t_L g2130 ( 
.A1(n_1788),
.A2(n_1518),
.B(n_1508),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1836),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1877),
.Y(n_2132)
);

OAI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1867),
.A2(n_1751),
.B(n_1725),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1768),
.A2(n_1760),
.B(n_1293),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1769),
.B(n_1518),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1769),
.A2(n_1294),
.B(n_1287),
.Y(n_2136)
);

AOI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_1771),
.A2(n_1306),
.B(n_1294),
.Y(n_2137)
);

O2A1O1Ixp5_ASAP7_75t_L g2138 ( 
.A1(n_1953),
.A2(n_1751),
.B(n_1725),
.C(n_1634),
.Y(n_2138)
);

A2O1A1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_1940),
.A2(n_1447),
.B(n_1448),
.C(n_1441),
.Y(n_2139)
);

AOI211xp5_ASAP7_75t_L g2140 ( 
.A1(n_1893),
.A2(n_670),
.B(n_676),
.C(n_665),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_1771),
.A2(n_1306),
.B(n_1453),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_1780),
.A2(n_1484),
.B(n_1453),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1780),
.A2(n_1484),
.B(n_1340),
.Y(n_2143)
);

BUFx6f_ASAP7_75t_L g2144 ( 
.A(n_1785),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1941),
.B(n_1621),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_1827),
.A2(n_1655),
.B1(n_1482),
.B2(n_1634),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1878),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1877),
.Y(n_2148)
);

AOI21x1_ASAP7_75t_L g2149 ( 
.A1(n_1788),
.A2(n_1305),
.B(n_1394),
.Y(n_2149)
);

OAI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_1872),
.A2(n_1638),
.B(n_1621),
.Y(n_2150)
);

OAI21xp33_ASAP7_75t_L g2151 ( 
.A1(n_1770),
.A2(n_593),
.B(n_590),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1881),
.B(n_1307),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1830),
.A2(n_1655),
.B1(n_1638),
.B2(n_1644),
.Y(n_2153)
);

A2O1A1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_1879),
.A2(n_1880),
.B(n_1913),
.C(n_1882),
.Y(n_2154)
);

AOI21x1_ASAP7_75t_L g2155 ( 
.A1(n_1777),
.A2(n_1520),
.B(n_1519),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1883),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_1895),
.A2(n_1606),
.B1(n_1645),
.B2(n_1590),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1881),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_1882),
.B(n_915),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1770),
.A2(n_1655),
.B1(n_1695),
.B2(n_1668),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1884),
.A2(n_1484),
.B(n_1391),
.Y(n_2161)
);

O2A1O1Ixp33_ASAP7_75t_L g2162 ( 
.A1(n_1884),
.A2(n_695),
.B(n_696),
.C(n_676),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_1886),
.A2(n_1340),
.B(n_1337),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_1886),
.A2(n_1337),
.B(n_1307),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1887),
.A2(n_1337),
.B(n_1307),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1887),
.Y(n_2166)
);

OR2x6_ASAP7_75t_L g2167 ( 
.A(n_1925),
.B(n_1606),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1888),
.B(n_1367),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_1774),
.A2(n_597),
.B(n_596),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1888),
.A2(n_1391),
.B(n_1319),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1892),
.Y(n_2171)
);

O2A1O1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_1892),
.A2(n_695),
.B(n_703),
.C(n_696),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1896),
.Y(n_2173)
);

OAI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1896),
.A2(n_1645),
.B1(n_1743),
.B2(n_1606),
.Y(n_2174)
);

A2O1A1Ixp33_ASAP7_75t_L g2175 ( 
.A1(n_1899),
.A2(n_1456),
.B(n_1463),
.C(n_1449),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_1894),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_1894),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_1899),
.A2(n_1367),
.B(n_1645),
.Y(n_2178)
);

AOI33xp33_ASAP7_75t_L g2179 ( 
.A1(n_1776),
.A2(n_710),
.A3(n_703),
.B1(n_723),
.B2(n_712),
.B3(n_709),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1777),
.A2(n_1743),
.B1(n_1458),
.B2(n_1506),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1778),
.A2(n_1458),
.B1(n_1506),
.B2(n_1501),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_1778),
.A2(n_1367),
.B(n_1174),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1774),
.B(n_1449),
.Y(n_2183)
);

OAI21x1_ASAP7_75t_L g2184 ( 
.A1(n_1910),
.A2(n_1501),
.B(n_1458),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1829),
.B(n_1456),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_1984),
.A2(n_1829),
.B1(n_1838),
.B2(n_1837),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2024),
.B(n_2035),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1975),
.B(n_1837),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2009),
.A2(n_2013),
.B(n_2030),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2085),
.B(n_1668),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2063),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2060),
.B(n_1924),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_2044),
.B(n_1910),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1972),
.B(n_1838),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2044),
.B(n_1910),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2030),
.A2(n_1391),
.B(n_1319),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1967),
.Y(n_2197)
);

A2O1A1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_2015),
.A2(n_710),
.B(n_712),
.C(n_709),
.Y(n_2198)
);

A2O1A1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_1971),
.A2(n_725),
.B(n_726),
.C(n_723),
.Y(n_2199)
);

AOI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_1983),
.A2(n_1391),
.B(n_1695),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2075),
.B(n_915),
.Y(n_2201)
);

BUFx2_ASAP7_75t_SL g2202 ( 
.A(n_2059),
.Y(n_2202)
);

NOR3xp33_ASAP7_75t_L g2203 ( 
.A(n_2026),
.B(n_922),
.C(n_917),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1968),
.B(n_1843),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1970),
.B(n_1843),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2082),
.B(n_1844),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1965),
.A2(n_2077),
.B1(n_1966),
.B2(n_2053),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1979),
.B(n_1957),
.Y(n_2208)
);

OAI22x1_ASAP7_75t_L g2209 ( 
.A1(n_2092),
.A2(n_2115),
.B1(n_2004),
.B2(n_2050),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2110),
.B(n_2094),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1983),
.A2(n_1391),
.B(n_1655),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1973),
.Y(n_2212)
);

A2O1A1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_1985),
.A2(n_726),
.B(n_728),
.C(n_725),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_1997),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2048),
.B(n_1957),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1976),
.B(n_1964),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1998),
.B(n_1844),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1996),
.B(n_1846),
.Y(n_2218)
);

OAI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2010),
.A2(n_1846),
.B1(n_1857),
.B2(n_1776),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2008),
.A2(n_1749),
.B(n_1465),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1999),
.A2(n_1749),
.B(n_1465),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1987),
.B(n_1749),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2179),
.B(n_1857),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1989),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_2052),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2005),
.B(n_2140),
.Y(n_2226)
);

O2A1O1Ixp33_ASAP7_75t_L g2227 ( 
.A1(n_2108),
.A2(n_735),
.B(n_736),
.C(n_734),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2033),
.A2(n_1749),
.B(n_1470),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_2022),
.B(n_599),
.Y(n_2229)
);

OAI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1988),
.A2(n_1921),
.B1(n_1929),
.B2(n_1925),
.Y(n_2230)
);

AOI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_1978),
.A2(n_1749),
.B(n_1470),
.Y(n_2231)
);

O2A1O1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2121),
.A2(n_744),
.B(n_748),
.C(n_736),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_1978),
.A2(n_2040),
.B(n_2042),
.Y(n_2233)
);

O2A1O1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_2122),
.A2(n_748),
.B(n_762),
.C(n_744),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2016),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2070),
.B(n_1749),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2071),
.B(n_1993),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_2038),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2020),
.Y(n_2239)
);

CKINVDCx16_ASAP7_75t_R g2240 ( 
.A(n_2049),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2040),
.A2(n_1472),
.B(n_1463),
.Y(n_2241)
);

O2A1O1Ixp5_ASAP7_75t_L g2242 ( 
.A1(n_2000),
.A2(n_1473),
.B(n_1475),
.C(n_1472),
.Y(n_2242)
);

AOI21xp33_ASAP7_75t_L g2243 ( 
.A1(n_1995),
.A2(n_1921),
.B(n_1929),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2034),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2114),
.A2(n_2105),
.B1(n_2002),
.B2(n_2167),
.Y(n_2245)
);

AO22x1_ASAP7_75t_L g2246 ( 
.A1(n_2036),
.A2(n_602),
.B1(n_608),
.B2(n_606),
.Y(n_2246)
);

NOR2xp67_ASAP7_75t_SL g2247 ( 
.A(n_2011),
.B(n_917),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2167),
.A2(n_1936),
.B1(n_1939),
.B2(n_1930),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2042),
.A2(n_1475),
.B(n_1473),
.Y(n_2249)
);

AOI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2143),
.A2(n_1495),
.B(n_1487),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2070),
.B(n_478),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2156),
.Y(n_2252)
);

A2O1A1Ixp33_ASAP7_75t_L g2253 ( 
.A1(n_1980),
.A2(n_770),
.B(n_777),
.C(n_762),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1994),
.B(n_1501),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2143),
.A2(n_1495),
.B(n_1487),
.Y(n_2255)
);

INVx4_ASAP7_75t_L g2256 ( 
.A(n_2144),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2111),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1974),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1990),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2038),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2158),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2005),
.B(n_1930),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_SL g2263 ( 
.A(n_2041),
.B(n_2078),
.Y(n_2263)
);

AO21x1_ASAP7_75t_L g2264 ( 
.A1(n_2067),
.A2(n_777),
.B(n_770),
.Y(n_2264)
);

CKINVDCx20_ASAP7_75t_R g2265 ( 
.A(n_2041),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2027),
.B(n_478),
.Y(n_2266)
);

O2A1O1Ixp33_ASAP7_75t_SL g2267 ( 
.A1(n_2081),
.A2(n_1507),
.B(n_1519),
.C(n_1496),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2159),
.B(n_922),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1982),
.A2(n_2046),
.B(n_2025),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_SL g2270 ( 
.A(n_2061),
.B(n_926),
.C(n_925),
.Y(n_2270)
);

A2O1A1Ixp33_ASAP7_75t_L g2271 ( 
.A1(n_1992),
.A2(n_2151),
.B(n_2169),
.C(n_2162),
.Y(n_2271)
);

O2A1O1Ixp5_ASAP7_75t_L g2272 ( 
.A1(n_2067),
.A2(n_1507),
.B(n_1520),
.C(n_1496),
.Y(n_2272)
);

OAI21x1_ASAP7_75t_L g2273 ( 
.A1(n_2170),
.A2(n_1506),
.B(n_1268),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_1982),
.A2(n_1939),
.B(n_1936),
.Y(n_2274)
);

O2A1O1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2183),
.A2(n_926),
.B(n_927),
.C(n_925),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2166),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2007),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2171),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_2038),
.B(n_609),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2102),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2027),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2045),
.A2(n_1956),
.B(n_1910),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_SL g2283 ( 
.A1(n_2116),
.A2(n_612),
.B1(n_614),
.B2(n_611),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_L g2284 ( 
.A(n_2066),
.B(n_619),
.Y(n_2284)
);

A2O1A1Ixp33_ASAP7_75t_L g2285 ( 
.A1(n_2172),
.A2(n_620),
.B(n_623),
.C(n_622),
.Y(n_2285)
);

INVx4_ASAP7_75t_L g2286 ( 
.A(n_2144),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2006),
.B(n_1956),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2101),
.A2(n_1136),
.B(n_1081),
.Y(n_2288)
);

A2O1A1Ixp33_ASAP7_75t_L g2289 ( 
.A1(n_2117),
.A2(n_624),
.B(n_626),
.C(n_625),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_2177),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2167),
.A2(n_631),
.B1(n_633),
.B2(n_628),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2017),
.B(n_634),
.Y(n_2292)
);

A2O1A1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_2117),
.A2(n_635),
.B(n_638),
.C(n_637),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2029),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2031),
.B(n_639),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2084),
.Y(n_2296)
);

A2O1A1Ixp33_ASAP7_75t_L g2297 ( 
.A1(n_2118),
.A2(n_640),
.B(n_644),
.C(n_641),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_SL g2298 ( 
.A1(n_2068),
.A2(n_927),
.B(n_1268),
.C(n_817),
.Y(n_2298)
);

O2A1O1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2032),
.A2(n_820),
.B(n_826),
.C(n_815),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2173),
.Y(n_2300)
);

O2A1O1Ixp5_ASAP7_75t_L g2301 ( 
.A1(n_2068),
.A2(n_820),
.B(n_827),
.C(n_826),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_1991),
.A2(n_1136),
.B(n_1081),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2093),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2113),
.A2(n_717),
.B1(n_753),
.B2(n_691),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2098),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2118),
.A2(n_2057),
.B(n_2072),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2161),
.A2(n_1136),
.B(n_1081),
.Y(n_2307)
);

AOI21xp33_ASAP7_75t_L g2308 ( 
.A1(n_2090),
.A2(n_647),
.B(n_645),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2086),
.B(n_649),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_2066),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2059),
.A2(n_652),
.B1(n_657),
.B2(n_656),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2120),
.Y(n_2312)
);

OA22x2_ASAP7_75t_L g2313 ( 
.A1(n_2153),
.A2(n_660),
.B1(n_666),
.B2(n_658),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_1981),
.B(n_691),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2132),
.A2(n_673),
.B1(n_675),
.B2(n_668),
.Y(n_2315)
);

BUFx12f_ASAP7_75t_L g2316 ( 
.A(n_2148),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2123),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2131),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2160),
.A2(n_679),
.B1(n_682),
.B2(n_677),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2037),
.B(n_683),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2146),
.B(n_717),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2001),
.B(n_685),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2147),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2058),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2144),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2091),
.B(n_717),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2001),
.B(n_2003),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2003),
.B(n_688),
.Y(n_2328)
);

O2A1O1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2185),
.A2(n_828),
.B(n_829),
.C(n_827),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_2021),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2154),
.A2(n_2019),
.B1(n_2047),
.B2(n_2028),
.Y(n_2331)
);

A2O1A1Ixp33_ASAP7_75t_SL g2332 ( 
.A1(n_2072),
.A2(n_829),
.B(n_832),
.C(n_828),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2112),
.A2(n_1136),
.B(n_1081),
.Y(n_2333)
);

O2A1O1Ixp33_ASAP7_75t_L g2334 ( 
.A1(n_2039),
.A2(n_833),
.B(n_836),
.C(n_832),
.Y(n_2334)
);

A2O1A1Ixp33_ASAP7_75t_L g2335 ( 
.A1(n_2100),
.A2(n_692),
.B(n_698),
.C(n_697),
.Y(n_2335)
);

NAND2xp33_ASAP7_75t_R g2336 ( 
.A(n_2109),
.B(n_388),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2089),
.B(n_1332),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2021),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_1986),
.B(n_699),
.Y(n_2339)
);

BUFx3_ASAP7_75t_L g2340 ( 
.A(n_2176),
.Y(n_2340)
);

INVx3_ASAP7_75t_SL g2341 ( 
.A(n_2097),
.Y(n_2341)
);

A2O1A1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_2145),
.A2(n_704),
.B(n_707),
.C(n_705),
.Y(n_2342)
);

BUFx4f_ASAP7_75t_SL g2343 ( 
.A(n_2021),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2103),
.A2(n_715),
.B1(n_719),
.B2(n_708),
.Y(n_2344)
);

O2A1O1Ixp33_ASAP7_75t_L g2345 ( 
.A1(n_2181),
.A2(n_836),
.B(n_837),
.C(n_833),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2062),
.B(n_720),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2065),
.A2(n_721),
.B1(n_727),
.B2(n_724),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2069),
.B(n_729),
.Y(n_2348)
);

BUFx2_ASAP7_75t_L g2349 ( 
.A(n_2021),
.Y(n_2349)
);

INVxp67_ASAP7_75t_L g2350 ( 
.A(n_2073),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2079),
.B(n_2014),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2127),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2128),
.Y(n_2353)
);

BUFx8_ASAP7_75t_SL g2354 ( 
.A(n_2130),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2055),
.B(n_737),
.Y(n_2355)
);

AOI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_1969),
.A2(n_740),
.B1(n_741),
.B2(n_739),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2064),
.B(n_2096),
.Y(n_2357)
);

INVxp67_ASAP7_75t_SL g2358 ( 
.A(n_2163),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2127),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2107),
.B(n_717),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2155),
.B(n_753),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_2095),
.A2(n_742),
.B(n_745),
.C(n_743),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2106),
.A2(n_1171),
.B(n_1169),
.Y(n_2363)
);

OAI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2129),
.A2(n_747),
.B1(n_749),
.B2(n_746),
.Y(n_2364)
);

O2A1O1Ixp33_ASAP7_75t_L g2365 ( 
.A1(n_2023),
.A2(n_838),
.B(n_841),
.C(n_837),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2135),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2157),
.A2(n_752),
.B1(n_754),
.B2(n_751),
.Y(n_2367)
);

A2O1A1Ixp33_ASAP7_75t_L g2368 ( 
.A1(n_2119),
.A2(n_2125),
.B(n_2124),
.C(n_2104),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2152),
.B(n_758),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2168),
.B(n_765),
.Y(n_2370)
);

O2A1O1Ixp5_ASAP7_75t_SL g2371 ( 
.A1(n_2174),
.A2(n_844),
.B(n_845),
.C(n_843),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2180),
.B(n_768),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2021),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2138),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2175),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_2043),
.B(n_769),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2139),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1977),
.B(n_772),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2133),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_1977),
.B(n_775),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2119),
.A2(n_1171),
.B(n_1169),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2012),
.Y(n_2382)
);

NAND2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2184),
.B(n_2080),
.Y(n_2383)
);

BUFx4f_ASAP7_75t_L g2384 ( 
.A(n_2083),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2012),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2125),
.A2(n_753),
.B1(n_760),
.B2(n_776),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2134),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2134),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2150),
.B(n_778),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2182),
.B(n_844),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2136),
.B(n_753),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2136),
.Y(n_2392)
);

A2O1A1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2099),
.A2(n_846),
.B(n_847),
.C(n_845),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2149),
.B(n_1429),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2137),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2012),
.B(n_760),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2099),
.A2(n_1171),
.B(n_1169),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2137),
.B(n_760),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2104),
.A2(n_1171),
.B(n_1169),
.Y(n_2399)
);

O2A1O1Ixp33_ASAP7_75t_L g2400 ( 
.A1(n_2126),
.A2(n_846),
.B(n_848),
.C(n_847),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2087),
.A2(n_2076),
.B1(n_2088),
.B2(n_2142),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2012),
.Y(n_2402)
);

AO32x2_ASAP7_75t_L g2403 ( 
.A1(n_2018),
.A2(n_760),
.A3(n_949),
.B1(n_947),
.B2(n_1429),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2051),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2164),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2051),
.B(n_2054),
.Y(n_2406)
);

O2A1O1Ixp33_ASAP7_75t_L g2407 ( 
.A1(n_2178),
.A2(n_850),
.B(n_851),
.C(n_848),
.Y(n_2407)
);

NAND2x2_ASAP7_75t_L g2408 ( 
.A(n_2018),
.B(n_3),
.Y(n_2408)
);

A2O1A1Ixp33_ASAP7_75t_L g2409 ( 
.A1(n_2142),
.A2(n_850),
.B(n_853),
.C(n_851),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2178),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2054),
.B(n_1429),
.Y(n_2411)
);

BUFx2_ASAP7_75t_L g2412 ( 
.A(n_2182),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2141),
.A2(n_1171),
.B(n_1169),
.Y(n_2413)
);

AOI22x1_ASAP7_75t_SL g2414 ( 
.A1(n_2018),
.A2(n_859),
.B1(n_860),
.B2(n_853),
.Y(n_2414)
);

OR2x6_ASAP7_75t_L g2415 ( 
.A(n_2141),
.B(n_859),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2164),
.B(n_860),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2056),
.B(n_481),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2165),
.B(n_870),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2074),
.Y(n_2419)
);

AOI21xp5_ASAP7_75t_L g2420 ( 
.A1(n_2165),
.A2(n_1182),
.B(n_1177),
.Y(n_2420)
);

OR2x6_ASAP7_75t_L g2421 ( 
.A(n_2167),
.B(n_870),
.Y(n_2421)
);

NOR2xp67_ASAP7_75t_L g2422 ( 
.A(n_2085),
.B(n_391),
.Y(n_2422)
);

INVx2_ASAP7_75t_SL g2423 ( 
.A(n_1997),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1984),
.B(n_871),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_1984),
.A2(n_873),
.B1(n_874),
.B2(n_871),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_1984),
.B(n_3),
.Y(n_2426)
);

A2O1A1Ixp33_ASAP7_75t_L g2427 ( 
.A1(n_2015),
.A2(n_873),
.B(n_874),
.C(n_1018),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2063),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_2044),
.B(n_392),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2024),
.B(n_1018),
.Y(n_2430)
);

AOI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2060),
.A2(n_481),
.B1(n_1517),
.B2(n_1032),
.Y(n_2431)
);

INVx5_ASAP7_75t_L g2432 ( 
.A(n_2144),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_L g2433 ( 
.A(n_1984),
.B(n_947),
.Y(n_2433)
);

AOI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2009),
.A2(n_1182),
.B(n_1177),
.Y(n_2434)
);

A2O1A1Ixp33_ASAP7_75t_L g2435 ( 
.A1(n_2015),
.A2(n_1028),
.B(n_1032),
.C(n_1030),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_1984),
.B(n_481),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2052),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2024),
.B(n_1028),
.Y(n_2438)
);

AO21x1_ASAP7_75t_L g2439 ( 
.A1(n_1965),
.A2(n_966),
.B(n_964),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2085),
.B(n_393),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1967),
.Y(n_2441)
);

NAND2x1p5_ASAP7_75t_L g2442 ( 
.A(n_2004),
.B(n_1177),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2085),
.B(n_396),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_1984),
.A2(n_1182),
.B1(n_1189),
.B2(n_1177),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_1984),
.A2(n_1182),
.B1(n_1189),
.B2(n_1177),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_1984),
.B(n_4),
.Y(n_2446)
);

OAI21x1_ASAP7_75t_L g2447 ( 
.A1(n_2189),
.A2(n_968),
.B(n_966),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2353),
.B(n_481),
.Y(n_2448)
);

AOI22x1_ASAP7_75t_L g2449 ( 
.A1(n_2209),
.A2(n_982),
.B1(n_986),
.B2(n_968),
.Y(n_2449)
);

OAI21x1_ASAP7_75t_L g2450 ( 
.A1(n_2211),
.A2(n_986),
.B(n_982),
.Y(n_2450)
);

A2O1A1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2271),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_2451)
);

BUFx12f_ASAP7_75t_L g2452 ( 
.A(n_2214),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2269),
.A2(n_1189),
.B(n_1182),
.Y(n_2453)
);

OAI21x1_ASAP7_75t_L g2454 ( 
.A1(n_2221),
.A2(n_1002),
.B(n_986),
.Y(n_2454)
);

A2O1A1Ixp33_ASAP7_75t_L g2455 ( 
.A1(n_2389),
.A2(n_9),
.B(n_6),
.C(n_8),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2191),
.B(n_481),
.Y(n_2456)
);

OAI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2289),
.A2(n_1517),
.B(n_1003),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2428),
.B(n_2350),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2210),
.B(n_397),
.Y(n_2459)
);

NOR2xp67_ASAP7_75t_L g2460 ( 
.A(n_2225),
.B(n_399),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2366),
.B(n_2207),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2224),
.Y(n_2462)
);

NAND3xp33_ASAP7_75t_SL g2463 ( 
.A(n_2304),
.B(n_1003),
.C(n_1002),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_L g2464 ( 
.A1(n_2228),
.A2(n_1003),
.B(n_1002),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2281),
.B(n_401),
.Y(n_2465)
);

BUFx10_ASAP7_75t_L g2466 ( 
.A(n_2423),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2261),
.Y(n_2467)
);

INVx4_ASAP7_75t_L g2468 ( 
.A(n_2432),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2350),
.B(n_8),
.Y(n_2469)
);

NAND3x1_ASAP7_75t_L g2470 ( 
.A(n_2192),
.B(n_10),
.C(n_12),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2237),
.B(n_990),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2293),
.A2(n_1517),
.B(n_1004),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2324),
.B(n_10),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2368),
.A2(n_1222),
.B(n_1189),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2187),
.B(n_404),
.Y(n_2475)
);

AOI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2233),
.A2(n_1222),
.B(n_1189),
.Y(n_2476)
);

AOI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2229),
.A2(n_1517),
.B1(n_1030),
.B2(n_1027),
.Y(n_2477)
);

INVx3_ASAP7_75t_SL g2478 ( 
.A(n_2290),
.Y(n_2478)
);

OAI21x1_ASAP7_75t_SL g2479 ( 
.A1(n_2282),
.A2(n_1004),
.B(n_12),
.Y(n_2479)
);

OAI21xp33_ASAP7_75t_L g2480 ( 
.A1(n_2304),
.A2(n_2386),
.B(n_2198),
.Y(n_2480)
);

OAI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2297),
.A2(n_1517),
.B(n_1004),
.Y(n_2481)
);

INVxp67_ASAP7_75t_SL g2482 ( 
.A(n_2318),
.Y(n_2482)
);

AOI21xp33_ASAP7_75t_L g2483 ( 
.A1(n_2380),
.A2(n_2355),
.B(n_2376),
.Y(n_2483)
);

BUFx3_ASAP7_75t_L g2484 ( 
.A(n_2280),
.Y(n_2484)
);

NAND2x1p5_ASAP7_75t_L g2485 ( 
.A(n_2384),
.B(n_2432),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2276),
.Y(n_2486)
);

OAI21xp33_ASAP7_75t_L g2487 ( 
.A1(n_2386),
.A2(n_1030),
.B(n_1027),
.Y(n_2487)
);

AO31x2_ASAP7_75t_L g2488 ( 
.A1(n_2439),
.A2(n_949),
.A3(n_1517),
.B(n_408),
.Y(n_2488)
);

INVx5_ASAP7_75t_L g2489 ( 
.A(n_2421),
.Y(n_2489)
);

A2O1A1Ixp33_ASAP7_75t_L g2490 ( 
.A1(n_2376),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2194),
.B(n_14),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2404),
.B(n_16),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_2237),
.B(n_990),
.Y(n_2493)
);

AO31x2_ASAP7_75t_L g2494 ( 
.A1(n_2264),
.A2(n_949),
.A3(n_409),
.B(n_418),
.Y(n_2494)
);

OAI21x1_ASAP7_75t_L g2495 ( 
.A1(n_2196),
.A2(n_997),
.B(n_985),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2278),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2426),
.B(n_16),
.Y(n_2497)
);

OAI21x1_ASAP7_75t_L g2498 ( 
.A1(n_2249),
.A2(n_997),
.B(n_985),
.Y(n_2498)
);

AO21x1_ASAP7_75t_L g2499 ( 
.A1(n_2360),
.A2(n_17),
.B(n_18),
.Y(n_2499)
);

OAI21x1_ASAP7_75t_L g2500 ( 
.A1(n_2250),
.A2(n_2255),
.B(n_2241),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2300),
.Y(n_2501)
);

AOI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2358),
.A2(n_1246),
.B(n_1222),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2197),
.Y(n_2503)
);

O2A1O1Ixp33_ASAP7_75t_SL g2504 ( 
.A1(n_2213),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2504)
);

OA21x2_ASAP7_75t_L g2505 ( 
.A1(n_2306),
.A2(n_19),
.B(n_21),
.Y(n_2505)
);

OAI21x1_ASAP7_75t_L g2506 ( 
.A1(n_2231),
.A2(n_997),
.B(n_985),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2206),
.B(n_2226),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2426),
.B(n_21),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2358),
.A2(n_1246),
.B(n_1222),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2212),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2235),
.Y(n_2511)
);

BUFx16f_ASAP7_75t_R g2512 ( 
.A(n_2429),
.Y(n_2512)
);

OAI21x1_ASAP7_75t_L g2513 ( 
.A1(n_2381),
.A2(n_1009),
.B(n_985),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2263),
.B(n_990),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_2357),
.A2(n_1246),
.B(n_1222),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_L g2516 ( 
.A1(n_2302),
.A2(n_1009),
.B(n_1027),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2351),
.B(n_22),
.Y(n_2517)
);

NAND3x1_ASAP7_75t_L g2518 ( 
.A(n_2188),
.B(n_23),
.C(n_25),
.Y(n_2518)
);

A2O1A1Ixp33_ASAP7_75t_L g2519 ( 
.A1(n_2372),
.A2(n_28),
.B(n_23),
.C(n_27),
.Y(n_2519)
);

A2O1A1Ixp33_ASAP7_75t_L g2520 ( 
.A1(n_2372),
.A2(n_31),
.B(n_27),
.C(n_29),
.Y(n_2520)
);

NAND3xp33_ASAP7_75t_SL g2521 ( 
.A(n_2309),
.B(n_29),
.C(n_32),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_SL g2522 ( 
.A(n_2343),
.B(n_949),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2325),
.Y(n_2523)
);

AO31x2_ASAP7_75t_L g2524 ( 
.A1(n_2274),
.A2(n_419),
.A3(n_421),
.B(n_406),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2421),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_2525)
);

AO31x2_ASAP7_75t_L g2526 ( 
.A1(n_2401),
.A2(n_424),
.A3(n_426),
.B(n_423),
.Y(n_2526)
);

AO31x2_ASAP7_75t_L g2527 ( 
.A1(n_2374),
.A2(n_429),
.A3(n_430),
.B(n_428),
.Y(n_2527)
);

OAI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2421),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2262),
.B(n_431),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2204),
.B(n_38),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_2288),
.A2(n_1247),
.B(n_1246),
.Y(n_2531)
);

AOI21x1_ASAP7_75t_L g2532 ( 
.A1(n_2208),
.A2(n_1247),
.B(n_1246),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2325),
.Y(n_2533)
);

INVx8_ASAP7_75t_L g2534 ( 
.A(n_2432),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2441),
.Y(n_2535)
);

OAI21x1_ASAP7_75t_L g2536 ( 
.A1(n_2272),
.A2(n_1009),
.B(n_1027),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2422),
.B(n_2240),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2325),
.Y(n_2538)
);

O2A1O1Ixp5_ASAP7_75t_SL g2539 ( 
.A1(n_2417),
.A2(n_1030),
.B(n_1009),
.C(n_42),
.Y(n_2539)
);

A2O1A1Ixp33_ASAP7_75t_L g2540 ( 
.A1(n_2234),
.A2(n_43),
.B(n_39),
.C(n_41),
.Y(n_2540)
);

OAI21x1_ASAP7_75t_L g2541 ( 
.A1(n_2434),
.A2(n_1253),
.B(n_1247),
.Y(n_2541)
);

AOI221x1_ASAP7_75t_L g2542 ( 
.A1(n_2219),
.A2(n_43),
.B1(n_39),
.B2(n_41),
.C(n_44),
.Y(n_2542)
);

BUFx10_ASAP7_75t_L g2543 ( 
.A(n_2279),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2205),
.B(n_45),
.Y(n_2544)
);

BUFx8_ASAP7_75t_L g2545 ( 
.A(n_2316),
.Y(n_2545)
);

OAI21xp33_ASAP7_75t_L g2546 ( 
.A1(n_2380),
.A2(n_1001),
.B(n_990),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_L g2547 ( 
.A(n_2437),
.B(n_2216),
.Y(n_2547)
);

AO32x2_ASAP7_75t_L g2548 ( 
.A1(n_2186),
.A2(n_47),
.A3(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2446),
.B(n_433),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2362),
.A2(n_1247),
.B(n_1253),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2239),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2325),
.Y(n_2552)
);

OAI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2378),
.A2(n_1022),
.B(n_991),
.Y(n_2553)
);

OAI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2331),
.A2(n_1022),
.B(n_991),
.Y(n_2554)
);

OAI21x1_ASAP7_75t_L g2555 ( 
.A1(n_2273),
.A2(n_1253),
.B(n_1247),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2384),
.B(n_990),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2244),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2217),
.B(n_46),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2440),
.B(n_438),
.Y(n_2559)
);

NAND2x1p5_ASAP7_75t_L g2560 ( 
.A(n_2432),
.B(n_1253),
.Y(n_2560)
);

OAI21x1_ASAP7_75t_L g2561 ( 
.A1(n_2406),
.A2(n_1253),
.B(n_444),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_2238),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2335),
.A2(n_1001),
.B(n_990),
.Y(n_2563)
);

OAI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2446),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_2564)
);

AO21x1_ASAP7_75t_L g2565 ( 
.A1(n_2230),
.A2(n_51),
.B(n_52),
.Y(n_2565)
);

OAI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2223),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_2566)
);

AOI21x1_ASAP7_75t_SL g2567 ( 
.A1(n_2396),
.A2(n_54),
.B(n_56),
.Y(n_2567)
);

OAI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2343),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_2568)
);

AO21x1_ASAP7_75t_L g2569 ( 
.A1(n_2319),
.A2(n_59),
.B(n_60),
.Y(n_2569)
);

OAI21x1_ASAP7_75t_L g2570 ( 
.A1(n_2333),
.A2(n_445),
.B(n_439),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2266),
.A2(n_1007),
.B1(n_1012),
.B2(n_1001),
.Y(n_2571)
);

AO32x2_ASAP7_75t_L g2572 ( 
.A1(n_2248),
.A2(n_2245),
.A3(n_2291),
.B1(n_2344),
.B2(n_2444),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2340),
.Y(n_2573)
);

AOI21x1_ASAP7_75t_L g2574 ( 
.A1(n_2391),
.A2(n_2398),
.B(n_2363),
.Y(n_2574)
);

INVxp67_ASAP7_75t_SL g2575 ( 
.A(n_2318),
.Y(n_2575)
);

NOR3xp33_ASAP7_75t_SL g2576 ( 
.A(n_2336),
.B(n_61),
.C(n_62),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2218),
.B(n_61),
.Y(n_2577)
);

OAI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2200),
.A2(n_448),
.B(n_447),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2443),
.B(n_449),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2260),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2257),
.Y(n_2581)
);

NOR2x1_ASAP7_75t_SL g2582 ( 
.A(n_2415),
.B(n_2330),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2238),
.Y(n_2583)
);

NAND3xp33_ASAP7_75t_L g2584 ( 
.A(n_2227),
.B(n_1007),
.C(n_1001),
.Y(n_2584)
);

OAI21x1_ASAP7_75t_L g2585 ( 
.A1(n_2383),
.A2(n_451),
.B(n_450),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2252),
.Y(n_2586)
);

OAI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2253),
.A2(n_1022),
.B(n_991),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2312),
.Y(n_2588)
);

AO31x2_ASAP7_75t_L g2589 ( 
.A1(n_2412),
.A2(n_454),
.A3(n_456),
.B(n_453),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2190),
.B(n_65),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2190),
.B(n_65),
.Y(n_2591)
);

INVx5_ASAP7_75t_L g2592 ( 
.A(n_2330),
.Y(n_2592)
);

O2A1O1Ixp5_ASAP7_75t_SL g2593 ( 
.A1(n_2308),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2408),
.A2(n_69),
.B1(n_66),
.B2(n_68),
.Y(n_2594)
);

AOI21x1_ASAP7_75t_L g2595 ( 
.A1(n_2397),
.A2(n_458),
.B(n_457),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2258),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2259),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2287),
.B(n_69),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2277),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2220),
.A2(n_977),
.B(n_955),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2313),
.B(n_2424),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2294),
.Y(n_2602)
);

OAI21x1_ASAP7_75t_SL g2603 ( 
.A1(n_2232),
.A2(n_70),
.B(n_71),
.Y(n_2603)
);

O2A1O1Ixp5_ASAP7_75t_L g2604 ( 
.A1(n_2243),
.A2(n_2321),
.B(n_2251),
.C(n_2436),
.Y(n_2604)
);

OAI22x1_ASAP7_75t_L g2605 ( 
.A1(n_2341),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_2605)
);

AOI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2415),
.A2(n_977),
.B(n_955),
.Y(n_2606)
);

OAI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2275),
.A2(n_1022),
.B(n_991),
.Y(n_2607)
);

INVx5_ASAP7_75t_L g2608 ( 
.A(n_2330),
.Y(n_2608)
);

OAI21x1_ASAP7_75t_L g2609 ( 
.A1(n_2301),
.A2(n_464),
.B(n_463),
.Y(n_2609)
);

INVx4_ASAP7_75t_SL g2610 ( 
.A(n_2341),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2296),
.Y(n_2611)
);

AO31x2_ASAP7_75t_L g2612 ( 
.A1(n_2352),
.A2(n_470),
.A3(n_472),
.B(n_465),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2411),
.A2(n_977),
.B(n_954),
.Y(n_2613)
);

OAI21x1_ASAP7_75t_L g2614 ( 
.A1(n_2301),
.A2(n_473),
.B(n_1001),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2339),
.B(n_72),
.Y(n_2615)
);

CKINVDCx20_ASAP7_75t_R g2616 ( 
.A(n_2265),
.Y(n_2616)
);

BUFx8_ASAP7_75t_SL g2617 ( 
.A(n_2238),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2242),
.A2(n_977),
.B(n_954),
.Y(n_2618)
);

OAI21x1_ASAP7_75t_L g2619 ( 
.A1(n_2420),
.A2(n_2413),
.B(n_2399),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2313),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2620)
);

AOI21xp33_ASAP7_75t_L g2621 ( 
.A1(n_2234),
.A2(n_74),
.B(n_76),
.Y(n_2621)
);

OAI21x1_ASAP7_75t_L g2622 ( 
.A1(n_2410),
.A2(n_1007),
.B(n_1001),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2379),
.B(n_76),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2254),
.B(n_77),
.Y(n_2624)
);

AO21x2_ASAP7_75t_L g2625 ( 
.A1(n_2332),
.A2(n_77),
.B(n_78),
.Y(n_2625)
);

NAND3x1_ASAP7_75t_L g2626 ( 
.A(n_2311),
.B(n_78),
.C(n_79),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2303),
.Y(n_2627)
);

OAI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2275),
.A2(n_1022),
.B(n_991),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2254),
.B(n_80),
.Y(n_2629)
);

AO31x2_ASAP7_75t_L g2630 ( 
.A1(n_2359),
.A2(n_82),
.A3(n_80),
.B(n_81),
.Y(n_2630)
);

A2O1A1Ixp33_ASAP7_75t_L g2631 ( 
.A1(n_2227),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2410),
.A2(n_2307),
.B(n_2242),
.Y(n_2632)
);

AO21x2_ASAP7_75t_L g2633 ( 
.A1(n_2298),
.A2(n_85),
.B(n_86),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2392),
.B(n_87),
.Y(n_2634)
);

OAI21x1_ASAP7_75t_L g2635 ( 
.A1(n_2365),
.A2(n_1012),
.B(n_1007),
.Y(n_2635)
);

OAI21x1_ASAP7_75t_L g2636 ( 
.A1(n_2365),
.A2(n_1012),
.B(n_1007),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2395),
.B(n_87),
.Y(n_2637)
);

NAND2xp33_ASAP7_75t_L g2638 ( 
.A(n_2215),
.B(n_2310),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_SL g2639 ( 
.A1(n_2285),
.A2(n_1012),
.B(n_1007),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2327),
.B(n_1012),
.Y(n_2640)
);

BUFx2_ASAP7_75t_L g2641 ( 
.A(n_2238),
.Y(n_2641)
);

OAI21x1_ASAP7_75t_L g2642 ( 
.A1(n_2416),
.A2(n_1012),
.B(n_956),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2430),
.B(n_89),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2232),
.B(n_89),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2193),
.B(n_90),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2305),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2438),
.B(n_90),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2193),
.B(n_91),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2195),
.B(n_92),
.Y(n_2649)
);

OAI21x1_ASAP7_75t_L g2650 ( 
.A1(n_2418),
.A2(n_956),
.B(n_991),
.Y(n_2650)
);

AOI21x1_ASAP7_75t_L g2651 ( 
.A1(n_2361),
.A2(n_956),
.B(n_93),
.Y(n_2651)
);

AO31x2_ASAP7_75t_L g2652 ( 
.A1(n_2394),
.A2(n_2388),
.A3(n_2387),
.B(n_2405),
.Y(n_2652)
);

BUFx2_ASAP7_75t_L g2653 ( 
.A(n_2256),
.Y(n_2653)
);

BUFx4f_ASAP7_75t_SL g2654 ( 
.A(n_2256),
.Y(n_2654)
);

AO31x2_ASAP7_75t_L g2655 ( 
.A1(n_2394),
.A2(n_96),
.A3(n_93),
.B(n_94),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2317),
.B(n_96),
.Y(n_2656)
);

INVx5_ASAP7_75t_L g2657 ( 
.A(n_2330),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2268),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2402),
.B(n_2222),
.Y(n_2659)
);

AOI21xp5_ASAP7_75t_L g2660 ( 
.A1(n_2267),
.A2(n_954),
.B(n_940),
.Y(n_2660)
);

OAI21xp33_ASAP7_75t_L g2661 ( 
.A1(n_2356),
.A2(n_97),
.B(n_100),
.Y(n_2661)
);

OR2x2_ASAP7_75t_L g2662 ( 
.A(n_2201),
.B(n_100),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2323),
.Y(n_2663)
);

CKINVDCx11_ASAP7_75t_R g2664 ( 
.A(n_2286),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_2202),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2390),
.B(n_101),
.Y(n_2666)
);

BUFx8_ASAP7_75t_L g2667 ( 
.A(n_2429),
.Y(n_2667)
);

OAI21x1_ASAP7_75t_SL g2668 ( 
.A1(n_2329),
.A2(n_102),
.B(n_104),
.Y(n_2668)
);

OAI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2299),
.A2(n_1022),
.B(n_1048),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2373),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2433),
.B(n_1048),
.Y(n_2671)
);

OAI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2299),
.A2(n_1048),
.B(n_102),
.Y(n_2672)
);

NOR2xp67_ASAP7_75t_L g2673 ( 
.A(n_2286),
.B(n_104),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_L g2674 ( 
.A(n_2195),
.Y(n_2674)
);

INVx5_ASAP7_75t_L g2675 ( 
.A(n_2354),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2419),
.A2(n_954),
.B(n_940),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2369),
.B(n_105),
.Y(n_2677)
);

OA21x2_ASAP7_75t_L g2678 ( 
.A1(n_2382),
.A2(n_105),
.B(n_106),
.Y(n_2678)
);

BUFx3_ASAP7_75t_L g2679 ( 
.A(n_2337),
.Y(n_2679)
);

NAND3x1_ASAP7_75t_L g2680 ( 
.A(n_2328),
.B(n_107),
.C(n_109),
.Y(n_2680)
);

INVx3_ASAP7_75t_L g2681 ( 
.A(n_2338),
.Y(n_2681)
);

NAND2x1p5_ASAP7_75t_L g2682 ( 
.A(n_2338),
.B(n_940),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_2349),
.Y(n_2683)
);

OAI21x1_ASAP7_75t_L g2684 ( 
.A1(n_2400),
.A2(n_956),
.B(n_107),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2385),
.Y(n_2685)
);

OR2x6_ASAP7_75t_L g2686 ( 
.A(n_2442),
.B(n_956),
.Y(n_2686)
);

OAI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2400),
.A2(n_109),
.B(n_110),
.Y(n_2687)
);

OAI21x1_ASAP7_75t_L g2688 ( 
.A1(n_2371),
.A2(n_111),
.B(n_113),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2375),
.Y(n_2689)
);

INVx3_ASAP7_75t_L g2690 ( 
.A(n_2337),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2442),
.B(n_113),
.Y(n_2691)
);

OAI21x1_ASAP7_75t_L g2692 ( 
.A1(n_2407),
.A2(n_114),
.B(n_115),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2407),
.Y(n_2693)
);

OR2x6_ASAP7_75t_L g2694 ( 
.A(n_2329),
.B(n_115),
.Y(n_2694)
);

INVx8_ASAP7_75t_L g2695 ( 
.A(n_2236),
.Y(n_2695)
);

OAI21x1_ASAP7_75t_L g2696 ( 
.A1(n_2334),
.A2(n_116),
.B(n_118),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2445),
.A2(n_954),
.B(n_940),
.Y(n_2697)
);

AO31x2_ASAP7_75t_L g2698 ( 
.A1(n_2377),
.A2(n_121),
.A3(n_119),
.B(n_120),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2393),
.Y(n_2699)
);

A2O1A1Ixp33_ASAP7_75t_L g2700 ( 
.A1(n_2483),
.A2(n_2199),
.B(n_2342),
.C(n_2314),
.Y(n_2700)
);

OAI21x1_ASAP7_75t_SL g2701 ( 
.A1(n_2479),
.A2(n_2345),
.B(n_2334),
.Y(n_2701)
);

OAI21xp5_ASAP7_75t_L g2702 ( 
.A1(n_2483),
.A2(n_2326),
.B(n_2322),
.Y(n_2702)
);

AO21x2_ASAP7_75t_L g2703 ( 
.A1(n_2476),
.A2(n_2270),
.B(n_2345),
.Y(n_2703)
);

OAI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2604),
.A2(n_2328),
.B(n_2284),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2467),
.Y(n_2705)
);

AO31x2_ASAP7_75t_L g2706 ( 
.A1(n_2453),
.A2(n_2409),
.A3(n_2435),
.B(n_2427),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2486),
.Y(n_2707)
);

BUFx2_ASAP7_75t_SL g2708 ( 
.A(n_2675),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2496),
.Y(n_2709)
);

OAI21x1_ASAP7_75t_L g2710 ( 
.A1(n_2500),
.A2(n_2425),
.B(n_2431),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2501),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2652),
.Y(n_2712)
);

OAI21x1_ASAP7_75t_SL g2713 ( 
.A1(n_2565),
.A2(n_2370),
.B(n_2367),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2503),
.Y(n_2714)
);

OA21x2_ASAP7_75t_L g2715 ( 
.A1(n_2474),
.A2(n_2203),
.B(n_2292),
.Y(n_2715)
);

OAI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2490),
.A2(n_2284),
.B(n_2295),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2510),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2616),
.B(n_2246),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2511),
.Y(n_2719)
);

AO21x2_ASAP7_75t_L g2720 ( 
.A1(n_2502),
.A2(n_2270),
.B(n_2203),
.Y(n_2720)
);

HB1xp67_ASAP7_75t_L g2721 ( 
.A(n_2462),
.Y(n_2721)
);

AOI21x1_ASAP7_75t_L g2722 ( 
.A1(n_2651),
.A2(n_2320),
.B(n_2346),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2543),
.B(n_2283),
.Y(n_2723)
);

AO21x2_ASAP7_75t_L g2724 ( 
.A1(n_2509),
.A2(n_2403),
.B(n_2348),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2535),
.Y(n_2725)
);

AOI21x1_ASAP7_75t_L g2726 ( 
.A1(n_2595),
.A2(n_2347),
.B(n_2364),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2670),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2461),
.B(n_2247),
.Y(n_2728)
);

NOR2xp67_ASAP7_75t_L g2729 ( 
.A(n_2675),
.B(n_119),
.Y(n_2729)
);

OR2x2_ASAP7_75t_L g2730 ( 
.A(n_2652),
.B(n_120),
.Y(n_2730)
);

HB1xp67_ASAP7_75t_L g2731 ( 
.A(n_2683),
.Y(n_2731)
);

OAI21x1_ASAP7_75t_L g2732 ( 
.A1(n_2619),
.A2(n_2403),
.B(n_2414),
.Y(n_2732)
);

OAI21x1_ASAP7_75t_L g2733 ( 
.A1(n_2650),
.A2(n_2403),
.B(n_121),
.Y(n_2733)
);

AO21x2_ASAP7_75t_L g2734 ( 
.A1(n_2574),
.A2(n_2403),
.B(n_2315),
.Y(n_2734)
);

BUFx3_ASAP7_75t_L g2735 ( 
.A(n_2617),
.Y(n_2735)
);

OAI21x1_ASAP7_75t_L g2736 ( 
.A1(n_2531),
.A2(n_122),
.B(n_123),
.Y(n_2736)
);

AO21x2_ASAP7_75t_L g2737 ( 
.A1(n_2515),
.A2(n_2600),
.B(n_2613),
.Y(n_2737)
);

OA21x2_ASAP7_75t_L g2738 ( 
.A1(n_2632),
.A2(n_122),
.B(n_123),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2685),
.B(n_124),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2551),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2480),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2557),
.Y(n_2742)
);

AO21x2_ASAP7_75t_L g2743 ( 
.A1(n_2554),
.A2(n_127),
.B(n_128),
.Y(n_2743)
);

OAI21x1_ASAP7_75t_L g2744 ( 
.A1(n_2642),
.A2(n_127),
.B(n_128),
.Y(n_2744)
);

BUFx2_ASAP7_75t_R g2745 ( 
.A(n_2665),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2461),
.B(n_129),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2659),
.B(n_129),
.Y(n_2747)
);

AOI31xp67_ASAP7_75t_L g2748 ( 
.A1(n_2601),
.A2(n_132),
.A3(n_130),
.B(n_131),
.Y(n_2748)
);

INVx1_ASAP7_75t_SL g2749 ( 
.A(n_2664),
.Y(n_2749)
);

AO31x2_ASAP7_75t_L g2750 ( 
.A1(n_2660),
.A2(n_133),
.A3(n_131),
.B(n_132),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2543),
.B(n_136),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2581),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2586),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2588),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2596),
.Y(n_2755)
);

OAI21x1_ASAP7_75t_L g2756 ( 
.A1(n_2541),
.A2(n_136),
.B(n_137),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2478),
.B(n_137),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2547),
.B(n_138),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2681),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2659),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2681),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2554),
.A2(n_940),
.B(n_1048),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2635),
.A2(n_139),
.B(n_140),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2546),
.A2(n_1048),
.B(n_139),
.Y(n_2764)
);

OAI21x1_ASAP7_75t_L g2765 ( 
.A1(n_2636),
.A2(n_140),
.B(n_141),
.Y(n_2765)
);

OR2x6_ASAP7_75t_L g2766 ( 
.A(n_2534),
.B(n_141),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_SL g2767 ( 
.A(n_2452),
.B(n_142),
.Y(n_2767)
);

INVx2_ASAP7_75t_SL g2768 ( 
.A(n_2534),
.Y(n_2768)
);

CKINVDCx11_ASAP7_75t_R g2769 ( 
.A(n_2466),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2482),
.Y(n_2770)
);

OAI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2451),
.A2(n_142),
.B(n_143),
.Y(n_2771)
);

OAI21x1_ASAP7_75t_L g2772 ( 
.A1(n_2495),
.A2(n_146),
.B(n_147),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2678),
.Y(n_2773)
);

A2O1A1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2661),
.A2(n_2615),
.B(n_2576),
.C(n_2455),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2545),
.Y(n_2775)
);

BUFx10_ASAP7_75t_L g2776 ( 
.A(n_2465),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2575),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2683),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2573),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2597),
.Y(n_2780)
);

O2A1O1Ixp33_ASAP7_75t_L g2781 ( 
.A1(n_2519),
.A2(n_2520),
.B(n_2521),
.C(n_2540),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2602),
.Y(n_2782)
);

OAI21x1_ASAP7_75t_L g2783 ( 
.A1(n_2555),
.A2(n_146),
.B(n_147),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2611),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2599),
.Y(n_2785)
);

OAI21x1_ASAP7_75t_L g2786 ( 
.A1(n_2516),
.A2(n_148),
.B(n_149),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2507),
.B(n_149),
.Y(n_2787)
);

OAI21x1_ASAP7_75t_L g2788 ( 
.A1(n_2561),
.A2(n_150),
.B(n_154),
.Y(n_2788)
);

OAI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2675),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2678),
.Y(n_2790)
);

AO32x2_ASAP7_75t_L g2791 ( 
.A1(n_2566),
.A2(n_157),
.A3(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_2791)
);

OAI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2470),
.A2(n_161),
.B1(n_157),
.B2(n_160),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2607),
.A2(n_161),
.B(n_163),
.Y(n_2793)
);

BUFx2_ASAP7_75t_L g2794 ( 
.A(n_2505),
.Y(n_2794)
);

BUFx12f_ASAP7_75t_L g2795 ( 
.A(n_2466),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2627),
.Y(n_2796)
);

OAI21x1_ASAP7_75t_L g2797 ( 
.A1(n_2447),
.A2(n_164),
.B(n_165),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2653),
.Y(n_2798)
);

OAI21x1_ASAP7_75t_L g2799 ( 
.A1(n_2614),
.A2(n_166),
.B(n_167),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2630),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2523),
.Y(n_2801)
);

BUFx3_ASAP7_75t_L g2802 ( 
.A(n_2552),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2630),
.Y(n_2803)
);

HB1xp67_ASAP7_75t_L g2804 ( 
.A(n_2458),
.Y(n_2804)
);

OAI21x1_ASAP7_75t_SL g2805 ( 
.A1(n_2582),
.A2(n_168),
.B(n_169),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2505),
.B(n_387),
.Y(n_2806)
);

AOI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2607),
.A2(n_168),
.B(n_170),
.Y(n_2807)
);

NOR2xp67_ASAP7_75t_L g2808 ( 
.A(n_2469),
.B(n_171),
.Y(n_2808)
);

OA21x2_ASAP7_75t_L g2809 ( 
.A1(n_2684),
.A2(n_172),
.B(n_174),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2630),
.Y(n_2810)
);

OAI21x1_ASAP7_75t_L g2811 ( 
.A1(n_2622),
.A2(n_386),
.B(n_172),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2628),
.A2(n_174),
.B(n_175),
.Y(n_2812)
);

OAI21x1_ASAP7_75t_L g2813 ( 
.A1(n_2513),
.A2(n_386),
.B(n_175),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2634),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2634),
.Y(n_2815)
);

AO31x2_ASAP7_75t_L g2816 ( 
.A1(n_2542),
.A2(n_176),
.A3(n_177),
.B(n_178),
.Y(n_2816)
);

OAI21x1_ASAP7_75t_L g2817 ( 
.A1(n_2609),
.A2(n_385),
.B(n_177),
.Y(n_2817)
);

NAND2x1p5_ASAP7_75t_L g2818 ( 
.A(n_2592),
.B(n_179),
.Y(n_2818)
);

A2O1A1Ixp33_ASAP7_75t_L g2819 ( 
.A1(n_2672),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2637),
.Y(n_2820)
);

OA21x2_ASAP7_75t_L g2821 ( 
.A1(n_2553),
.A2(n_182),
.B(n_185),
.Y(n_2821)
);

OAI21x1_ASAP7_75t_L g2822 ( 
.A1(n_2450),
.A2(n_385),
.B(n_182),
.Y(n_2822)
);

INVx4_ASAP7_75t_L g2823 ( 
.A(n_2534),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2578),
.A2(n_384),
.B(n_185),
.Y(n_2824)
);

BUFx2_ASAP7_75t_L g2825 ( 
.A(n_2641),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2637),
.Y(n_2826)
);

AOI21xp33_ASAP7_75t_L g2827 ( 
.A1(n_2517),
.A2(n_187),
.B(n_188),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2533),
.Y(n_2828)
);

O2A1O1Ixp33_ASAP7_75t_SL g2829 ( 
.A1(n_2631),
.A2(n_188),
.B(n_189),
.C(n_191),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2646),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2620),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_2831)
);

OAI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2621),
.A2(n_192),
.B(n_194),
.Y(n_2832)
);

BUFx2_ASAP7_75t_L g2833 ( 
.A(n_2580),
.Y(n_2833)
);

AO31x2_ASAP7_75t_L g2834 ( 
.A1(n_2594),
.A2(n_194),
.A3(n_195),
.B(n_196),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_L g2835 ( 
.A1(n_2620),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_2835)
);

OR2x6_ASAP7_75t_L g2836 ( 
.A(n_2485),
.B(n_199),
.Y(n_2836)
);

AOI21x1_ASAP7_75t_L g2837 ( 
.A1(n_2532),
.A2(n_200),
.B(n_201),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2663),
.Y(n_2838)
);

AOI21x1_ASAP7_75t_L g2839 ( 
.A1(n_2676),
.A2(n_200),
.B(n_202),
.Y(n_2839)
);

INVx8_ASAP7_75t_L g2840 ( 
.A(n_2592),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2533),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2680),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2492),
.B(n_203),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_SL g2844 ( 
.A(n_2484),
.B(n_205),
.Y(n_2844)
);

AO21x2_ASAP7_75t_L g2845 ( 
.A1(n_2672),
.A2(n_2553),
.B(n_2606),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2517),
.B(n_208),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2624),
.B(n_2629),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_2545),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2624),
.B(n_208),
.Y(n_2849)
);

OAI21x1_ASAP7_75t_L g2850 ( 
.A1(n_2506),
.A2(n_209),
.B(n_211),
.Y(n_2850)
);

AOI22xp33_ASAP7_75t_L g2851 ( 
.A1(n_2566),
.A2(n_209),
.B1(n_212),
.B2(n_214),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2689),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2621),
.A2(n_214),
.B(n_215),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2654),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2698),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2533),
.Y(n_2856)
);

OAI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2536),
.A2(n_384),
.B(n_216),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_L g2858 ( 
.A(n_2492),
.B(n_217),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2698),
.Y(n_2859)
);

OAI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2644),
.A2(n_217),
.B(n_218),
.Y(n_2860)
);

OAI21x1_ASAP7_75t_L g2861 ( 
.A1(n_2454),
.A2(n_383),
.B(n_220),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2538),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_SL g2863 ( 
.A1(n_2644),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_2863)
);

NAND3xp33_ASAP7_75t_SL g2864 ( 
.A(n_2569),
.B(n_2564),
.C(n_2508),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2475),
.B(n_221),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2538),
.Y(n_2866)
);

OAI21x1_ASAP7_75t_L g2867 ( 
.A1(n_2464),
.A2(n_225),
.B(n_226),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2593),
.A2(n_225),
.B(n_226),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2628),
.A2(n_227),
.B(n_229),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2610),
.Y(n_2870)
);

A2O1A1Ixp33_ASAP7_75t_L g2871 ( 
.A1(n_2559),
.A2(n_230),
.B(n_231),
.C(n_232),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2698),
.Y(n_2872)
);

OAI21x1_ASAP7_75t_L g2873 ( 
.A1(n_2498),
.A2(n_383),
.B(n_233),
.Y(n_2873)
);

NOR2xp67_ASAP7_75t_L g2874 ( 
.A(n_2623),
.B(n_235),
.Y(n_2874)
);

OAI21x1_ASAP7_75t_L g2875 ( 
.A1(n_2570),
.A2(n_382),
.B(n_236),
.Y(n_2875)
);

OAI21x1_ASAP7_75t_L g2876 ( 
.A1(n_2697),
.A2(n_382),
.B(n_236),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2618),
.A2(n_381),
.B(n_237),
.Y(n_2877)
);

INVxp67_ASAP7_75t_SL g2878 ( 
.A(n_2471),
.Y(n_2878)
);

AO21x1_ASAP7_75t_L g2879 ( 
.A1(n_2594),
.A2(n_235),
.B(n_237),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2655),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2655),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2564),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2449),
.A2(n_238),
.B(n_241),
.Y(n_2883)
);

HB1xp67_ASAP7_75t_L g2884 ( 
.A(n_2610),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2592),
.B(n_2608),
.Y(n_2885)
);

AO21x2_ASAP7_75t_L g2886 ( 
.A1(n_2550),
.A2(n_243),
.B(n_244),
.Y(n_2886)
);

OAI21x1_ASAP7_75t_L g2887 ( 
.A1(n_2585),
.A2(n_243),
.B(n_244),
.Y(n_2887)
);

AND2x4_ASAP7_75t_L g2888 ( 
.A(n_2608),
.B(n_245),
.Y(n_2888)
);

A2O1A1Ixp33_ASAP7_75t_L g2889 ( 
.A1(n_2579),
.A2(n_2497),
.B(n_2460),
.C(n_2590),
.Y(n_2889)
);

BUFx2_ASAP7_75t_L g2890 ( 
.A(n_2695),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2591),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_2891)
);

OA21x2_ASAP7_75t_L g2892 ( 
.A1(n_2688),
.A2(n_2687),
.B(n_2696),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2629),
.B(n_246),
.Y(n_2893)
);

AO21x2_ASAP7_75t_L g2894 ( 
.A1(n_2493),
.A2(n_249),
.B(n_250),
.Y(n_2894)
);

BUFx2_ASAP7_75t_L g2895 ( 
.A(n_2695),
.Y(n_2895)
);

BUFx2_ASAP7_75t_L g2896 ( 
.A(n_2695),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2669),
.A2(n_250),
.B(n_251),
.Y(n_2897)
);

OAI21x1_ASAP7_75t_L g2898 ( 
.A1(n_2669),
.A2(n_251),
.B(n_252),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2655),
.B(n_252),
.Y(n_2899)
);

AO31x2_ASAP7_75t_L g2900 ( 
.A1(n_2499),
.A2(n_253),
.A3(n_254),
.B(n_255),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2448),
.Y(n_2901)
);

CKINVDCx6p67_ASAP7_75t_R g2902 ( 
.A(n_2489),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2448),
.Y(n_2903)
);

OAI22xp33_ASAP7_75t_SL g2904 ( 
.A1(n_2694),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2589),
.Y(n_2905)
);

AO21x2_ASAP7_75t_L g2906 ( 
.A1(n_2625),
.A2(n_2633),
.B(n_2563),
.Y(n_2906)
);

BUFx3_ASAP7_75t_L g2907 ( 
.A(n_2538),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2639),
.A2(n_2584),
.B(n_2556),
.Y(n_2908)
);

AND2x4_ASAP7_75t_L g2909 ( 
.A(n_2608),
.B(n_256),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2694),
.A2(n_256),
.B1(n_258),
.B2(n_260),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2677),
.B(n_258),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2584),
.A2(n_260),
.B(n_261),
.Y(n_2912)
);

OAI211xp5_ASAP7_75t_L g2913 ( 
.A1(n_2568),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2491),
.B(n_265),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2623),
.Y(n_2915)
);

OAI21x1_ASAP7_75t_SL g2916 ( 
.A1(n_2668),
.A2(n_265),
.B(n_267),
.Y(n_2916)
);

OAI21x1_ASAP7_75t_L g2917 ( 
.A1(n_2692),
.A2(n_381),
.B(n_268),
.Y(n_2917)
);

INVx3_ASAP7_75t_L g2918 ( 
.A(n_2612),
.Y(n_2918)
);

OAI21x1_ASAP7_75t_L g2919 ( 
.A1(n_2539),
.A2(n_267),
.B(n_268),
.Y(n_2919)
);

CKINVDCx11_ASAP7_75t_R g2920 ( 
.A(n_2512),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2491),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2549),
.B(n_269),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2527),
.Y(n_2923)
);

BUFx2_ASAP7_75t_L g2924 ( 
.A(n_2610),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2709),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2709),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2714),
.Y(n_2927)
);

BUFx3_ASAP7_75t_L g2928 ( 
.A(n_2795),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2804),
.B(n_2530),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2714),
.Y(n_2930)
);

BUFx2_ASAP7_75t_R g2931 ( 
.A(n_2775),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2753),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2753),
.Y(n_2933)
);

CKINVDCx6p67_ASAP7_75t_R g2934 ( 
.A(n_2769),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2754),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2754),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2755),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2705),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2721),
.B(n_2530),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2707),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2711),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2717),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2755),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2760),
.B(n_2526),
.Y(n_2944)
);

HB1xp67_ASAP7_75t_L g2945 ( 
.A(n_2731),
.Y(n_2945)
);

CKINVDCx11_ASAP7_75t_R g2946 ( 
.A(n_2769),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2795),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2782),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2719),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2794),
.B(n_2526),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2740),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2742),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2752),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2794),
.B(n_2526),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2864),
.A2(n_2626),
.B1(n_2638),
.B2(n_2537),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2782),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2727),
.B(n_2524),
.Y(n_2957)
);

AND2x4_ASAP7_75t_L g2958 ( 
.A(n_2801),
.B(n_2657),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2784),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2727),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2784),
.Y(n_2961)
);

AOI21x1_ASAP7_75t_L g2962 ( 
.A1(n_2837),
.A2(n_2691),
.B(n_2666),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2770),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2777),
.Y(n_2964)
);

AND2x4_ASAP7_75t_L g2965 ( 
.A(n_2801),
.B(n_2657),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2725),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_SL g2967 ( 
.A1(n_2704),
.A2(n_2568),
.B1(n_2489),
.B2(n_2694),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2780),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2852),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2852),
.Y(n_2970)
);

BUFx2_ASAP7_75t_L g2971 ( 
.A(n_2825),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2727),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2785),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2712),
.B(n_2524),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_SL g2975 ( 
.A1(n_2860),
.A2(n_2489),
.B1(n_2603),
.B2(n_2528),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_L g2976 ( 
.A1(n_2879),
.A2(n_2525),
.B1(n_2528),
.B2(n_2605),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2785),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2712),
.B(n_2524),
.Y(n_2978)
);

INVx5_ASAP7_75t_L g2979 ( 
.A(n_2836),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2796),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2796),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_SL g2982 ( 
.A1(n_2758),
.A2(n_2525),
.B1(n_2658),
.B2(n_2544),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2830),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2830),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2778),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2838),
.Y(n_2986)
);

BUFx2_ASAP7_75t_L g2987 ( 
.A(n_2825),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2759),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2730),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2880),
.B(n_2881),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2730),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2800),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2773),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2803),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2810),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2773),
.Y(n_2996)
);

AOI22xp33_ASAP7_75t_SL g2997 ( 
.A1(n_2771),
.A2(n_2658),
.B1(n_2667),
.B2(n_2512),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2774),
.A2(n_2518),
.B1(n_2571),
.B2(n_2544),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2790),
.Y(n_2999)
);

OA21x2_ASAP7_75t_L g3000 ( 
.A1(n_2855),
.A2(n_2558),
.B(n_2691),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2859),
.Y(n_3001)
);

CKINVDCx20_ASAP7_75t_R g3002 ( 
.A(n_2854),
.Y(n_3002)
);

INVx5_ASAP7_75t_L g3003 ( 
.A(n_2836),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2879),
.A2(n_2667),
.B1(n_2645),
.B2(n_2649),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2872),
.Y(n_3005)
);

BUFx8_ASAP7_75t_L g3006 ( 
.A(n_2888),
.Y(n_3006)
);

OAI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2851),
.A2(n_2558),
.B1(n_2577),
.B2(n_2598),
.Y(n_3007)
);

AO21x2_ASAP7_75t_L g3008 ( 
.A1(n_2905),
.A2(n_2625),
.B(n_2633),
.Y(n_3008)
);

AND2x6_ASAP7_75t_L g3009 ( 
.A(n_2885),
.B(n_2465),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2790),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2759),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2905),
.B(n_2548),
.Y(n_3012)
);

AOI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2832),
.A2(n_2648),
.B1(n_2649),
.B2(n_2645),
.Y(n_3013)
);

CKINVDCx11_ASAP7_75t_R g3014 ( 
.A(n_2854),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2738),
.Y(n_3015)
);

AO21x2_ASAP7_75t_L g3016 ( 
.A1(n_2906),
.A2(n_2666),
.B(n_2640),
.Y(n_3016)
);

CKINVDCx6p67_ASAP7_75t_R g3017 ( 
.A(n_2708),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_2802),
.B(n_2657),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2814),
.Y(n_3019)
);

NAND2x1p5_ASAP7_75t_L g3020 ( 
.A(n_2924),
.B(n_2468),
.Y(n_3020)
);

OAI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_2819),
.A2(n_2648),
.B1(n_2485),
.B2(n_2473),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2815),
.Y(n_3022)
);

OR2x6_ASAP7_75t_L g3023 ( 
.A(n_2840),
.B(n_2708),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2728),
.B(n_2473),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2820),
.Y(n_3025)
);

AO21x1_ASAP7_75t_L g3026 ( 
.A1(n_2899),
.A2(n_2548),
.B(n_2456),
.Y(n_3026)
);

OAI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2910),
.A2(n_2673),
.B1(n_2679),
.B2(n_2690),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2826),
.Y(n_3028)
);

OAI21xp33_ASAP7_75t_SL g3029 ( 
.A1(n_2899),
.A2(n_2548),
.B(n_2514),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2833),
.Y(n_3030)
);

AO21x1_ASAP7_75t_SL g3031 ( 
.A1(n_2806),
.A2(n_2693),
.B(n_2567),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2921),
.B(n_2643),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2923),
.B(n_2589),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2833),
.Y(n_3034)
);

AOI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_2853),
.A2(n_2529),
.B1(n_2463),
.B2(n_2699),
.Y(n_3035)
);

AOI22xp33_ASAP7_75t_L g3036 ( 
.A1(n_2716),
.A2(n_2487),
.B1(n_2647),
.B2(n_2690),
.Y(n_3036)
);

HB1xp67_ASAP7_75t_L g3037 ( 
.A(n_2798),
.Y(n_3037)
);

NAND2x1p5_ASAP7_75t_L g3038 ( 
.A(n_2924),
.B(n_2468),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2915),
.B(n_2662),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2806),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2802),
.Y(n_3041)
);

AO21x2_ASAP7_75t_L g3042 ( 
.A1(n_2906),
.A2(n_2671),
.B(n_2504),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2738),
.Y(n_3043)
);

HB1xp67_ASAP7_75t_L g3044 ( 
.A(n_2798),
.Y(n_3044)
);

OAI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2844),
.A2(n_2674),
.B1(n_2522),
.B2(n_2656),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2738),
.Y(n_3046)
);

OAI22xp5_ASAP7_75t_L g3047 ( 
.A1(n_2831),
.A2(n_2674),
.B1(n_2477),
.B2(n_2459),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_2835),
.A2(n_2674),
.B1(n_2472),
.B2(n_2481),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2903),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2903),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2923),
.B(n_2589),
.Y(n_3051)
);

INVxp33_ASAP7_75t_L g3052 ( 
.A(n_2718),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2901),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2759),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2702),
.A2(n_2457),
.B1(n_2472),
.B2(n_2481),
.Y(n_3055)
);

BUFx8_ASAP7_75t_L g3056 ( 
.A(n_2888),
.Y(n_3056)
);

INVx1_ASAP7_75t_SL g3057 ( 
.A(n_2779),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_2792),
.A2(n_2457),
.B1(n_2562),
.B2(n_2583),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2842),
.A2(n_2583),
.B1(n_2562),
.B2(n_2686),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2843),
.A2(n_2858),
.B1(n_2713),
.B2(n_2863),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_2761),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2918),
.Y(n_3062)
);

BUFx2_ASAP7_75t_L g3063 ( 
.A(n_2870),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2847),
.B(n_2527),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_L g3065 ( 
.A1(n_2871),
.A2(n_2686),
.B1(n_2560),
.B2(n_2682),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_SL g3066 ( 
.A1(n_2913),
.A2(n_2572),
.B1(n_2522),
.B2(n_2686),
.Y(n_3066)
);

INVx6_ASAP7_75t_L g3067 ( 
.A(n_2776),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2747),
.B(n_2527),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_SL g3069 ( 
.A1(n_2713),
.A2(n_2572),
.B1(n_2587),
.B2(n_2682),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2761),
.Y(n_3070)
);

OAI22xp5_ASAP7_75t_SL g3071 ( 
.A1(n_2775),
.A2(n_2572),
.B1(n_2587),
.B2(n_2494),
.Y(n_3071)
);

NAND2x1_ASAP7_75t_L g3072 ( 
.A(n_2885),
.B(n_2494),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2918),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2918),
.Y(n_3074)
);

OAI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2836),
.A2(n_2494),
.B1(n_2488),
.B2(n_273),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2761),
.Y(n_3076)
);

CKINVDCx6p67_ASAP7_75t_R g3077 ( 
.A(n_2735),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2724),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2747),
.Y(n_3079)
);

BUFx10_ASAP7_75t_L g3080 ( 
.A(n_2848),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_L g3081 ( 
.A1(n_2836),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2724),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2878),
.Y(n_3083)
);

OAI21x1_ASAP7_75t_SL g3084 ( 
.A1(n_2793),
.A2(n_2488),
.B(n_276),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2748),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2748),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2735),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2914),
.B(n_2874),
.Y(n_3088)
);

OA21x2_ASAP7_75t_L g3089 ( 
.A1(n_2877),
.A2(n_2488),
.B(n_277),
.Y(n_3089)
);

OAI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2766),
.A2(n_272),
.B1(n_277),
.B2(n_278),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2739),
.Y(n_3091)
);

CKINVDCx16_ASAP7_75t_R g3092 ( 
.A(n_2749),
.Y(n_3092)
);

INVx6_ASAP7_75t_L g3093 ( 
.A(n_2776),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_SL g3094 ( 
.A(n_2766),
.Y(n_3094)
);

CKINVDCx8_ASAP7_75t_R g3095 ( 
.A(n_2848),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2724),
.Y(n_3096)
);

OAI21x1_ASAP7_75t_L g3097 ( 
.A1(n_2710),
.A2(n_279),
.B(n_280),
.Y(n_3097)
);

INVx3_ASAP7_75t_L g3098 ( 
.A(n_2902),
.Y(n_3098)
);

OAI21x1_ASAP7_75t_L g3099 ( 
.A1(n_2710),
.A2(n_281),
.B(n_282),
.Y(n_3099)
);

INVx6_ASAP7_75t_L g3100 ( 
.A(n_2776),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2739),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2897),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_3102)
);

CKINVDCx11_ASAP7_75t_R g3103 ( 
.A(n_2920),
.Y(n_3103)
);

AO21x2_ASAP7_75t_L g3104 ( 
.A1(n_2734),
.A2(n_285),
.B(n_286),
.Y(n_3104)
);

INVx4_ASAP7_75t_L g3105 ( 
.A(n_2902),
.Y(n_3105)
);

AOI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_2807),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_3106)
);

INVx6_ASAP7_75t_L g3107 ( 
.A(n_2840),
.Y(n_3107)
);

BUFx3_ASAP7_75t_L g3108 ( 
.A(n_2828),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2900),
.Y(n_3109)
);

AOI21x1_ASAP7_75t_L g3110 ( 
.A1(n_2837),
.A2(n_287),
.B(n_288),
.Y(n_3110)
);

OAI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_2741),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_3111)
);

OAI21xp5_ASAP7_75t_SL g3112 ( 
.A1(n_3060),
.A2(n_2781),
.B(n_2889),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3010),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_3041),
.B(n_2884),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2993),
.Y(n_3115)
);

AND2x2_ASAP7_75t_SL g3116 ( 
.A(n_2950),
.B(n_2821),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_3041),
.B(n_2890),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2997),
.A2(n_2976),
.B1(n_3066),
.B2(n_2967),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2982),
.A2(n_2882),
.B1(n_2891),
.B2(n_2827),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2930),
.Y(n_3120)
);

OAI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2979),
.A2(n_2812),
.B1(n_2869),
.B2(n_2766),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2993),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_3102),
.A2(n_2904),
.B1(n_2789),
.B2(n_2911),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_3106),
.A2(n_2743),
.B1(n_2922),
.B2(n_2846),
.Y(n_3124)
);

OAI21xp5_ASAP7_75t_SL g3125 ( 
.A1(n_2955),
.A2(n_2700),
.B(n_2723),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_3111),
.A2(n_2743),
.B1(n_2914),
.B2(n_2849),
.Y(n_3126)
);

AOI22xp33_ASAP7_75t_L g3127 ( 
.A1(n_2998),
.A2(n_2743),
.B1(n_2893),
.B2(n_2808),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2975),
.A2(n_2916),
.B1(n_2886),
.B2(n_2821),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2932),
.Y(n_3129)
);

AOI222xp33_ASAP7_75t_L g3130 ( 
.A1(n_3029),
.A2(n_2868),
.B1(n_2767),
.B2(n_2746),
.C1(n_2751),
.C2(n_2865),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2996),
.Y(n_3131)
);

OAI21xp33_ASAP7_75t_L g3132 ( 
.A1(n_3081),
.A2(n_2766),
.B(n_2818),
.Y(n_3132)
);

AOI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_3094),
.A2(n_2920),
.B1(n_2886),
.B2(n_2757),
.Y(n_3133)
);

HB1xp67_ASAP7_75t_L g3134 ( 
.A(n_3040),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_3052),
.B(n_2787),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_3052),
.B(n_2787),
.Y(n_3136)
);

INVx3_ASAP7_75t_L g3137 ( 
.A(n_3098),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2933),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3024),
.B(n_2734),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2935),
.Y(n_3140)
);

OAI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_3004),
.A2(n_2818),
.B1(n_2912),
.B2(n_2909),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2996),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2936),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2971),
.Y(n_3144)
);

BUFx5_ASAP7_75t_L g3145 ( 
.A(n_3033),
.Y(n_3145)
);

CKINVDCx5p33_ASAP7_75t_R g3146 ( 
.A(n_3014),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_3055),
.A2(n_3090),
.B1(n_3007),
.B2(n_3026),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_3026),
.A2(n_2916),
.B1(n_2886),
.B2(n_2821),
.Y(n_3148)
);

OAI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2979),
.A2(n_2818),
.B1(n_2908),
.B2(n_2895),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2979),
.A2(n_2909),
.B1(n_2888),
.B2(n_2896),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2999),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_2971),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2999),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_3030),
.B(n_2890),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_3071),
.A2(n_2845),
.B1(n_2764),
.B2(n_2734),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_3035),
.A2(n_2845),
.B1(n_2715),
.B2(n_2894),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_3024),
.A2(n_3094),
.B1(n_3031),
.B2(n_3036),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2987),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_SL g3159 ( 
.A1(n_2979),
.A2(n_2805),
.B1(n_2845),
.B2(n_2894),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_3094),
.A2(n_3031),
.B1(n_3021),
.B2(n_3003),
.Y(n_3160)
);

INVxp67_ASAP7_75t_L g3161 ( 
.A(n_2945),
.Y(n_3161)
);

INVx3_ASAP7_75t_SL g3162 ( 
.A(n_2934),
.Y(n_3162)
);

OAI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2979),
.A2(n_2895),
.B1(n_2896),
.B2(n_2729),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_3003),
.A2(n_2715),
.B1(n_2894),
.B2(n_2809),
.Y(n_3164)
);

AOI22xp33_ASAP7_75t_SL g3165 ( 
.A1(n_3003),
.A2(n_2805),
.B1(n_2715),
.B2(n_2840),
.Y(n_3165)
);

OAI22xp33_ASAP7_75t_L g3166 ( 
.A1(n_3003),
.A2(n_2823),
.B1(n_2840),
.B2(n_2809),
.Y(n_3166)
);

OAI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_3003),
.A2(n_2909),
.B1(n_2885),
.B2(n_2856),
.Y(n_3167)
);

OAI222xp33_ASAP7_75t_L g3168 ( 
.A1(n_3088),
.A2(n_2722),
.B1(n_2791),
.B2(n_2839),
.C1(n_2726),
.C2(n_2823),
.Y(n_3168)
);

AOI22xp33_ASAP7_75t_L g3169 ( 
.A1(n_3084),
.A2(n_2809),
.B1(n_2898),
.B2(n_2701),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_3014),
.Y(n_3170)
);

INVx3_ASAP7_75t_L g3171 ( 
.A(n_3098),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_3013),
.A2(n_2866),
.B1(n_2856),
.B2(n_2745),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_3059),
.A2(n_2866),
.B1(n_2823),
.B2(n_2768),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2969),
.Y(n_3174)
);

INVx4_ASAP7_75t_L g3175 ( 
.A(n_2934),
.Y(n_3175)
);

OAI22xp33_ASAP7_75t_L g3176 ( 
.A1(n_3017),
.A2(n_2791),
.B1(n_2768),
.B2(n_2839),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_2987),
.Y(n_3177)
);

OAI21xp33_ASAP7_75t_L g3178 ( 
.A1(n_2989),
.A2(n_2722),
.B(n_2736),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_3084),
.A2(n_2898),
.B1(n_2701),
.B2(n_2917),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3037),
.B(n_3044),
.Y(n_3180)
);

OAI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3069),
.A2(n_2907),
.B1(n_2862),
.B2(n_2828),
.Y(n_3181)
);

OAI22xp33_ASAP7_75t_L g3182 ( 
.A1(n_3017),
.A2(n_2791),
.B1(n_2726),
.B2(n_2834),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_SL g3183 ( 
.A1(n_3027),
.A2(n_2917),
.B1(n_2791),
.B2(n_2736),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_3104),
.A2(n_2720),
.B1(n_2892),
.B2(n_2876),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_3079),
.B(n_2862),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2970),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2956),
.Y(n_3187)
);

OAI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_3105),
.A2(n_2791),
.B1(n_2834),
.B2(n_2907),
.Y(n_3188)
);

BUFx12f_ASAP7_75t_L g3189 ( 
.A(n_2946),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_3083),
.B(n_2834),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2959),
.Y(n_3191)
);

OAI21xp33_ASAP7_75t_L g3192 ( 
.A1(n_2991),
.A2(n_2788),
.B(n_2876),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2929),
.B(n_2834),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_3104),
.A2(n_2720),
.B1(n_2892),
.B2(n_2703),
.Y(n_3194)
);

INVx4_ASAP7_75t_L g3195 ( 
.A(n_3077),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3034),
.B(n_2841),
.Y(n_3196)
);

INVx2_ASAP7_75t_SL g3197 ( 
.A(n_3087),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2925),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2925),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2926),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2926),
.Y(n_3201)
);

OAI21xp33_ASAP7_75t_L g3202 ( 
.A1(n_2950),
.A2(n_2788),
.B(n_2887),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_3104),
.A2(n_2720),
.B1(n_2892),
.B2(n_2703),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_3048),
.A2(n_2703),
.B1(n_2919),
.B2(n_2732),
.Y(n_3204)
);

AOI221xp5_ASAP7_75t_L g3205 ( 
.A1(n_3075),
.A2(n_2829),
.B1(n_2841),
.B2(n_2834),
.C(n_2762),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_2985),
.B(n_2732),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2927),
.Y(n_3207)
);

HB1xp67_ASAP7_75t_L g3208 ( 
.A(n_2972),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_3045),
.A2(n_2816),
.B1(n_2900),
.B2(n_2750),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2927),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2966),
.B(n_2737),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_3047),
.A2(n_2919),
.B1(n_2875),
.B2(n_2824),
.Y(n_3212)
);

OAI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_3058),
.A2(n_2816),
.B1(n_2900),
.B2(n_2750),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3063),
.B(n_2988),
.Y(n_3214)
);

AOI211x1_ASAP7_75t_L g3215 ( 
.A1(n_2939),
.A2(n_2816),
.B(n_291),
.C(n_292),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_3065),
.A2(n_2816),
.B1(n_2900),
.B2(n_2750),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3063),
.B(n_2737),
.Y(n_3217)
);

OAI21xp5_ASAP7_75t_SL g3218 ( 
.A1(n_2954),
.A2(n_2816),
.B(n_2900),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_3002),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_3103),
.A2(n_2875),
.B1(n_2824),
.B2(n_2887),
.Y(n_3220)
);

INVx5_ASAP7_75t_L g3221 ( 
.A(n_3080),
.Y(n_3221)
);

OAI21xp33_ASAP7_75t_L g3222 ( 
.A1(n_2954),
.A2(n_3068),
.B(n_3064),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2963),
.B(n_2750),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_3009),
.A2(n_2737),
.B1(n_2744),
.B2(n_2817),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2937),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_3095),
.A2(n_2750),
.B1(n_2883),
.B2(n_2817),
.Y(n_3226)
);

AOI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_3103),
.A2(n_2883),
.B1(n_2799),
.B2(n_2733),
.Y(n_3227)
);

OAI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_3095),
.A2(n_2799),
.B1(n_2811),
.B2(n_2756),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_3002),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3076),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_3000),
.A2(n_2733),
.B1(n_2873),
.B2(n_2850),
.Y(n_3231)
);

OAI21xp5_ASAP7_75t_SL g3232 ( 
.A1(n_3098),
.A2(n_289),
.B(n_293),
.Y(n_3232)
);

OAI21xp33_ASAP7_75t_L g3233 ( 
.A1(n_2974),
.A2(n_2744),
.B(n_2783),
.Y(n_3233)
);

OAI22x1_ASAP7_75t_L g3234 ( 
.A1(n_3091),
.A2(n_2783),
.B1(n_2756),
.B2(n_2765),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2937),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2943),
.Y(n_3236)
);

OAI21xp5_ASAP7_75t_SL g3237 ( 
.A1(n_2974),
.A2(n_293),
.B(n_294),
.Y(n_3237)
);

CKINVDCx20_ASAP7_75t_R g3238 ( 
.A(n_3092),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2943),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2948),
.Y(n_3240)
);

OAI222xp33_ASAP7_75t_L g3241 ( 
.A1(n_3105),
.A2(n_2811),
.B1(n_2772),
.B2(n_2873),
.C1(n_2850),
.C2(n_2813),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2948),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3000),
.A2(n_2867),
.B1(n_2861),
.B2(n_2763),
.Y(n_3243)
);

AOI22xp33_ASAP7_75t_L g3244 ( 
.A1(n_3000),
.A2(n_2867),
.B1(n_2861),
.B2(n_2763),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_3032),
.A2(n_2765),
.B1(n_2822),
.B2(n_2813),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2964),
.B(n_2857),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_SL g3247 ( 
.A(n_3105),
.B(n_2772),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3076),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_3039),
.A2(n_3016),
.B1(n_3101),
.B2(n_3042),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_SL g3250 ( 
.A1(n_3006),
.A2(n_2822),
.B1(n_2786),
.B2(n_2797),
.Y(n_3250)
);

CKINVDCx5p33_ASAP7_75t_R g3251 ( 
.A(n_2946),
.Y(n_3251)
);

AOI222xp33_ASAP7_75t_L g3252 ( 
.A1(n_3012),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.C1(n_299),
.C2(n_300),
.Y(n_3252)
);

AOI222xp33_ASAP7_75t_L g3253 ( 
.A1(n_3012),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.C1(n_299),
.C2(n_300),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_3080),
.Y(n_3254)
);

OAI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3097),
.A2(n_2786),
.B(n_2797),
.Y(n_3255)
);

INVx3_ASAP7_75t_L g3256 ( 
.A(n_2988),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2961),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2988),
.B(n_2857),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_SL g3259 ( 
.A1(n_3006),
.A2(n_3056),
.B1(n_3009),
.B2(n_2978),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_SL g3260 ( 
.A(n_3087),
.B(n_2706),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3077),
.A2(n_2706),
.B1(n_302),
.B2(n_304),
.Y(n_3261)
);

AOI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_3016),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3053),
.B(n_2706),
.Y(n_3263)
);

BUFx5_ASAP7_75t_L g3264 ( 
.A(n_3033),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3016),
.A2(n_2706),
.B(n_307),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_3042),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_2928),
.A2(n_2706),
.B1(n_311),
.B2(n_312),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3042),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_2960),
.Y(n_3269)
);

AOI22xp33_ASAP7_75t_L g3270 ( 
.A1(n_3006),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3011),
.B(n_314),
.Y(n_3271)
);

BUFx2_ASAP7_75t_L g3272 ( 
.A(n_3108),
.Y(n_3272)
);

INVxp67_ASAP7_75t_L g3273 ( 
.A(n_3135),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3113),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3134),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_3221),
.B(n_3023),
.Y(n_3276)
);

AND2x4_ASAP7_75t_L g3277 ( 
.A(n_3221),
.B(n_3023),
.Y(n_3277)
);

XNOR2xp5_ASAP7_75t_L g3278 ( 
.A(n_3238),
.B(n_3057),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_SL g3279 ( 
.A(n_3189),
.B(n_2931),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_3221),
.B(n_3023),
.Y(n_3280)
);

NAND2xp33_ASAP7_75t_R g3281 ( 
.A(n_3251),
.B(n_3023),
.Y(n_3281)
);

CKINVDCx8_ASAP7_75t_R g3282 ( 
.A(n_3146),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_R g3283 ( 
.A(n_3170),
.B(n_3080),
.Y(n_3283)
);

BUFx3_ASAP7_75t_L g3284 ( 
.A(n_3162),
.Y(n_3284)
);

AND2x4_ASAP7_75t_L g3285 ( 
.A(n_3221),
.B(n_3108),
.Y(n_3285)
);

INVx8_ASAP7_75t_L g3286 ( 
.A(n_3219),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3180),
.B(n_3020),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3120),
.Y(n_3288)
);

BUFx3_ASAP7_75t_L g3289 ( 
.A(n_3162),
.Y(n_3289)
);

NAND2xp33_ASAP7_75t_R g3290 ( 
.A(n_3229),
.B(n_2958),
.Y(n_3290)
);

NAND2xp33_ASAP7_75t_R g3291 ( 
.A(n_3137),
.B(n_3171),
.Y(n_3291)
);

NAND2xp33_ASAP7_75t_R g3292 ( 
.A(n_3137),
.B(n_2958),
.Y(n_3292)
);

NAND2xp33_ASAP7_75t_R g3293 ( 
.A(n_3171),
.B(n_2958),
.Y(n_3293)
);

NAND2xp33_ASAP7_75t_R g3294 ( 
.A(n_3272),
.B(n_2965),
.Y(n_3294)
);

NAND2xp33_ASAP7_75t_R g3295 ( 
.A(n_3152),
.B(n_3177),
.Y(n_3295)
);

AND2x4_ASAP7_75t_L g3296 ( 
.A(n_3254),
.B(n_3197),
.Y(n_3296)
);

NAND2xp33_ASAP7_75t_R g3297 ( 
.A(n_3271),
.B(n_2965),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3163),
.B(n_3087),
.Y(n_3298)
);

NOR2xp33_ASAP7_75t_R g3299 ( 
.A(n_3175),
.B(n_3195),
.Y(n_3299)
);

AND2x4_ASAP7_75t_L g3300 ( 
.A(n_3254),
.B(n_2990),
.Y(n_3300)
);

BUFx3_ASAP7_75t_L g3301 ( 
.A(n_3175),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_R g3302 ( 
.A(n_3195),
.B(n_3056),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_R g3303 ( 
.A(n_3270),
.B(n_3056),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3129),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3138),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3139),
.B(n_3193),
.Y(n_3306)
);

CKINVDCx12_ASAP7_75t_R g3307 ( 
.A(n_3117),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3161),
.B(n_3019),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3222),
.B(n_3022),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_R g3310 ( 
.A(n_3270),
.B(n_3087),
.Y(n_3310)
);

AND2x4_ASAP7_75t_L g3311 ( 
.A(n_3114),
.B(n_2990),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3206),
.B(n_3025),
.Y(n_3312)
);

INVxp67_ASAP7_75t_L g3313 ( 
.A(n_3135),
.Y(n_3313)
);

CKINVDCx16_ASAP7_75t_R g3314 ( 
.A(n_3172),
.Y(n_3314)
);

OR2x6_ASAP7_75t_L g3315 ( 
.A(n_3237),
.B(n_3107),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_R g3316 ( 
.A(n_3136),
.B(n_2928),
.Y(n_3316)
);

XNOR2xp5_ASAP7_75t_L g3317 ( 
.A(n_3118),
.B(n_2947),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_3154),
.B(n_3020),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3211),
.B(n_3028),
.Y(n_3319)
);

NAND2xp33_ASAP7_75t_R g3320 ( 
.A(n_3136),
.B(n_2965),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_R g3321 ( 
.A(n_3127),
.B(n_2947),
.Y(n_3321)
);

AND2x4_ASAP7_75t_L g3322 ( 
.A(n_3214),
.B(n_3018),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3190),
.B(n_2977),
.Y(n_3323)
);

AND2x4_ASAP7_75t_L g3324 ( 
.A(n_3258),
.B(n_3018),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_3125),
.B(n_3107),
.Y(n_3325)
);

XNOR2xp5_ASAP7_75t_L g3326 ( 
.A(n_3259),
.B(n_3038),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3140),
.B(n_2986),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_3185),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3143),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3144),
.B(n_3038),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3174),
.B(n_3186),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3187),
.B(n_2944),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_3158),
.B(n_3018),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3191),
.B(n_2944),
.Y(n_3334)
);

BUFx10_ASAP7_75t_L g3335 ( 
.A(n_3116),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3147),
.B(n_2968),
.Y(n_3336)
);

CKINVDCx5p33_ASAP7_75t_R g3337 ( 
.A(n_3150),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_3256),
.B(n_3011),
.Y(n_3338)
);

NAND2xp33_ASAP7_75t_R g3339 ( 
.A(n_3217),
.B(n_3011),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_L g3340 ( 
.A(n_3116),
.Y(n_3340)
);

XNOR2xp5_ASAP7_75t_L g3341 ( 
.A(n_3133),
.B(n_2938),
.Y(n_3341)
);

BUFx10_ASAP7_75t_L g3342 ( 
.A(n_3232),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_3167),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3198),
.Y(n_3344)
);

CKINVDCx5p33_ASAP7_75t_R g3345 ( 
.A(n_3181),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3199),
.Y(n_3346)
);

CKINVDCx5p33_ASAP7_75t_R g3347 ( 
.A(n_3173),
.Y(n_3347)
);

INVxp67_ASAP7_75t_L g3348 ( 
.A(n_3196),
.Y(n_3348)
);

AND2x4_ASAP7_75t_L g3349 ( 
.A(n_3256),
.B(n_3061),
.Y(n_3349)
);

CKINVDCx11_ASAP7_75t_R g3350 ( 
.A(n_3141),
.Y(n_3350)
);

NOR2xp33_ASAP7_75t_R g3351 ( 
.A(n_3127),
.B(n_3107),
.Y(n_3351)
);

NAND2xp33_ASAP7_75t_R g3352 ( 
.A(n_3246),
.B(n_3061),
.Y(n_3352)
);

BUFx3_ASAP7_75t_L g3353 ( 
.A(n_3269),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_R g3354 ( 
.A(n_3157),
.B(n_3107),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_R g3355 ( 
.A(n_3157),
.B(n_3160),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3147),
.B(n_2940),
.Y(n_3356)
);

INVxp67_ASAP7_75t_L g3357 ( 
.A(n_3112),
.Y(n_3357)
);

NAND2xp33_ASAP7_75t_R g3358 ( 
.A(n_3223),
.B(n_3061),
.Y(n_3358)
);

INVxp67_ASAP7_75t_L g3359 ( 
.A(n_3208),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_R g3360 ( 
.A(n_3160),
.B(n_3009),
.Y(n_3360)
);

BUFx10_ASAP7_75t_L g3361 ( 
.A(n_3201),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3188),
.B(n_2941),
.Y(n_3362)
);

BUFx12f_ASAP7_75t_L g3363 ( 
.A(n_3252),
.Y(n_3363)
);

INVxp67_ASAP7_75t_L g3364 ( 
.A(n_3130),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_3149),
.B(n_2960),
.Y(n_3365)
);

BUFx10_ASAP7_75t_L g3366 ( 
.A(n_3210),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_3247),
.B(n_3054),
.Y(n_3367)
);

NAND2xp33_ASAP7_75t_R g3368 ( 
.A(n_3263),
.B(n_3070),
.Y(n_3368)
);

BUFx6f_ASAP7_75t_L g3369 ( 
.A(n_3260),
.Y(n_3369)
);

NAND2xp33_ASAP7_75t_R g3370 ( 
.A(n_3225),
.B(n_2980),
.Y(n_3370)
);

BUFx3_ASAP7_75t_L g3371 ( 
.A(n_3230),
.Y(n_3371)
);

INVxp67_ASAP7_75t_L g3372 ( 
.A(n_3248),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3235),
.B(n_3067),
.Y(n_3373)
);

NAND2xp33_ASAP7_75t_R g3374 ( 
.A(n_3242),
.B(n_2981),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_3228),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3183),
.B(n_2942),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3257),
.B(n_3067),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3200),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_R g3379 ( 
.A(n_3123),
.B(n_3009),
.Y(n_3379)
);

INVxp67_ASAP7_75t_L g3380 ( 
.A(n_3200),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_R g3381 ( 
.A(n_3123),
.B(n_3009),
.Y(n_3381)
);

NAND2xp33_ASAP7_75t_R g3382 ( 
.A(n_3265),
.B(n_2960),
.Y(n_3382)
);

INVxp67_ASAP7_75t_L g3383 ( 
.A(n_3207),
.Y(n_3383)
);

XNOR2xp5_ASAP7_75t_L g3384 ( 
.A(n_3215),
.B(n_2949),
.Y(n_3384)
);

NAND2xp33_ASAP7_75t_R g3385 ( 
.A(n_3255),
.B(n_2973),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3155),
.B(n_2951),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_3121),
.B(n_3049),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3218),
.B(n_3249),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3207),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3236),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_R g3391 ( 
.A(n_3128),
.B(n_3009),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_R g3392 ( 
.A(n_3128),
.B(n_3067),
.Y(n_3392)
);

NAND2xp33_ASAP7_75t_R g3393 ( 
.A(n_3236),
.B(n_2973),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3239),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_R g3395 ( 
.A(n_3126),
.B(n_3067),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3155),
.B(n_2952),
.Y(n_3396)
);

CKINVDCx16_ASAP7_75t_R g3397 ( 
.A(n_3261),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3239),
.Y(n_3398)
);

OR2x2_ASAP7_75t_L g3399 ( 
.A(n_3249),
.B(n_2983),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3148),
.B(n_2953),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3165),
.B(n_3050),
.Y(n_3401)
);

AND2x4_ASAP7_75t_L g3402 ( 
.A(n_3240),
.B(n_3001),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_R g3403 ( 
.A(n_3126),
.B(n_3093),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_R g3404 ( 
.A(n_3266),
.B(n_3093),
.Y(n_3404)
);

AND2x4_ASAP7_75t_L g3405 ( 
.A(n_3240),
.B(n_3005),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_R g3406 ( 
.A(n_3253),
.B(n_2983),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3273),
.B(n_3205),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3288),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3402),
.Y(n_3409)
);

OR2x2_ASAP7_75t_L g3410 ( 
.A(n_3400),
.B(n_3216),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3304),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3402),
.Y(n_3412)
);

INVx2_ASAP7_75t_SL g3413 ( 
.A(n_3284),
.Y(n_3413)
);

BUFx3_ASAP7_75t_L g3414 ( 
.A(n_3289),
.Y(n_3414)
);

NOR2xp67_ASAP7_75t_SL g3415 ( 
.A(n_3397),
.B(n_3093),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3405),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3405),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3305),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3329),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3340),
.B(n_3115),
.Y(n_3420)
);

INVx2_ASAP7_75t_SL g3421 ( 
.A(n_3301),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3274),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3394),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_3299),
.Y(n_3424)
);

NOR2x1p5_ASAP7_75t_L g3425 ( 
.A(n_3363),
.B(n_3072),
.Y(n_3425)
);

OAI221xp5_ASAP7_75t_L g3426 ( 
.A1(n_3364),
.A2(n_3124),
.B1(n_3119),
.B2(n_3132),
.C(n_3148),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3340),
.B(n_3115),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3344),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3335),
.B(n_3145),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3361),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3361),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3346),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3313),
.B(n_3159),
.Y(n_3433)
);

AND2x2_ASAP7_75t_L g3434 ( 
.A(n_3335),
.B(n_3145),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3384),
.B(n_3124),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3366),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3366),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3340),
.B(n_3145),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3378),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3389),
.Y(n_3440)
);

NAND2x1p5_ASAP7_75t_SL g3441 ( 
.A(n_3401),
.B(n_3266),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3331),
.Y(n_3442)
);

HB1xp67_ASAP7_75t_L g3443 ( 
.A(n_3359),
.Y(n_3443)
);

INVxp67_ASAP7_75t_L g3444 ( 
.A(n_3406),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3324),
.B(n_3145),
.Y(n_3445)
);

INVxp67_ASAP7_75t_SL g3446 ( 
.A(n_3295),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3336),
.B(n_3176),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3390),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3356),
.B(n_3182),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3398),
.Y(n_3450)
);

INVxp67_ASAP7_75t_SL g3451 ( 
.A(n_3294),
.Y(n_3451)
);

NOR2x1_ASAP7_75t_L g3452 ( 
.A(n_3298),
.B(n_3166),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3324),
.B(n_3145),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3371),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3283),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3327),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3275),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3309),
.B(n_3156),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_3307),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3399),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3323),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3369),
.Y(n_3462)
);

CKINVDCx20_ASAP7_75t_R g3463 ( 
.A(n_3278),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3332),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3334),
.Y(n_3465)
);

INVx2_ASAP7_75t_SL g3466 ( 
.A(n_3285),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3386),
.B(n_3156),
.Y(n_3467)
);

NOR2xp33_ASAP7_75t_L g3468 ( 
.A(n_3357),
.B(n_3093),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3308),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3391),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3380),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3383),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3319),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3286),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3311),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3311),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_3360),
.Y(n_3477)
);

BUFx2_ASAP7_75t_L g3478 ( 
.A(n_3302),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3322),
.B(n_3145),
.Y(n_3479)
);

AND2x4_ASAP7_75t_L g3480 ( 
.A(n_3276),
.B(n_3122),
.Y(n_3480)
);

INVx1_ASAP7_75t_SL g3481 ( 
.A(n_3286),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3396),
.B(n_3209),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3353),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3322),
.B(n_3264),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3312),
.Y(n_3485)
);

BUFx2_ASAP7_75t_L g3486 ( 
.A(n_3316),
.Y(n_3486)
);

INVx2_ASAP7_75t_SL g3487 ( 
.A(n_3285),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3330),
.B(n_3264),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3372),
.Y(n_3489)
);

OR2x6_ASAP7_75t_L g3490 ( 
.A(n_3276),
.B(n_3226),
.Y(n_3490)
);

INVx2_ASAP7_75t_SL g3491 ( 
.A(n_3296),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3369),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3369),
.B(n_3373),
.Y(n_3493)
);

INVx4_ASAP7_75t_L g3494 ( 
.A(n_3342),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3362),
.Y(n_3495)
);

OA21x2_ASAP7_75t_L g3496 ( 
.A1(n_3388),
.A2(n_3203),
.B(n_3194),
.Y(n_3496)
);

OAI33xp33_ASAP7_75t_L g3497 ( 
.A1(n_3376),
.A2(n_3213),
.A3(n_3267),
.B1(n_3109),
.B2(n_3178),
.B3(n_2992),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3367),
.Y(n_3498)
);

BUFx2_ASAP7_75t_L g3499 ( 
.A(n_3392),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_3370),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3377),
.B(n_3264),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3367),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3300),
.B(n_3264),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3300),
.B(n_3264),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3306),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3333),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3333),
.B(n_3264),
.Y(n_3507)
);

HB1xp67_ASAP7_75t_L g3508 ( 
.A(n_3374),
.Y(n_3508)
);

NOR2xp33_ASAP7_75t_L g3509 ( 
.A(n_3279),
.B(n_3100),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3287),
.B(n_3122),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3387),
.Y(n_3511)
);

BUFx6f_ASAP7_75t_L g3512 ( 
.A(n_3342),
.Y(n_3512)
);

AOI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3350),
.A2(n_3119),
.B1(n_3268),
.B2(n_3262),
.Y(n_3513)
);

BUFx3_ASAP7_75t_L g3514 ( 
.A(n_3282),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3277),
.B(n_3131),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3277),
.B(n_3131),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3348),
.Y(n_3517)
);

BUFx2_ASAP7_75t_L g3518 ( 
.A(n_3280),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3280),
.B(n_3142),
.Y(n_3519)
);

OAI211xp5_ASAP7_75t_SL g3520 ( 
.A1(n_3365),
.A2(n_3268),
.B(n_3262),
.C(n_3202),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3338),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3318),
.B(n_3142),
.Y(n_3522)
);

CKINVDCx16_ASAP7_75t_R g3523 ( 
.A(n_3314),
.Y(n_3523)
);

OA21x2_ASAP7_75t_L g3524 ( 
.A1(n_3375),
.A2(n_3203),
.B(n_3194),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3341),
.B(n_3169),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_3393),
.Y(n_3526)
);

BUFx2_ASAP7_75t_L g3527 ( 
.A(n_3354),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3325),
.B(n_3100),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3296),
.B(n_3151),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3338),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3349),
.Y(n_3531)
);

OR2x2_ASAP7_75t_L g3532 ( 
.A(n_3349),
.B(n_3151),
.Y(n_3532)
);

AOI222xp33_ASAP7_75t_L g3533 ( 
.A1(n_3317),
.A2(n_3168),
.B1(n_3192),
.B2(n_3233),
.C1(n_3169),
.C2(n_3164),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3532),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3460),
.B(n_3315),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_3460),
.B(n_3315),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3532),
.Y(n_3537)
);

CKINVDCx16_ASAP7_75t_R g3538 ( 
.A(n_3523),
.Y(n_3538)
);

INVxp67_ASAP7_75t_L g3539 ( 
.A(n_3527),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3443),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3460),
.B(n_3153),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3408),
.Y(n_3542)
);

INVxp67_ASAP7_75t_SL g3543 ( 
.A(n_3500),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3523),
.B(n_3347),
.Y(n_3544)
);

OR2x2_ASAP7_75t_L g3545 ( 
.A(n_3461),
.B(n_3153),
.Y(n_3545)
);

INVxp67_ASAP7_75t_L g3546 ( 
.A(n_3527),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3495),
.B(n_3345),
.Y(n_3547)
);

INVx5_ASAP7_75t_L g3548 ( 
.A(n_3512),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3451),
.B(n_3337),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3408),
.Y(n_3550)
);

AND2x4_ASAP7_75t_SL g3551 ( 
.A(n_3459),
.B(n_3494),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3420),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3495),
.B(n_3321),
.Y(n_3553)
);

NAND2x1_ASAP7_75t_L g3554 ( 
.A(n_3415),
.B(n_3291),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3420),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3486),
.B(n_3355),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3411),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3411),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3511),
.B(n_3343),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3418),
.Y(n_3560)
);

OAI32xp33_ASAP7_75t_L g3561 ( 
.A1(n_3444),
.A2(n_3385),
.A3(n_3358),
.B1(n_3352),
.B2(n_3368),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3420),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3418),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3511),
.B(n_3379),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3420),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3486),
.B(n_3395),
.Y(n_3566)
);

INVxp67_ASAP7_75t_SL g3567 ( 
.A(n_3508),
.Y(n_3567)
);

OR2x6_ASAP7_75t_L g3568 ( 
.A(n_3512),
.B(n_3097),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3427),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3427),
.Y(n_3570)
);

INVx2_ASAP7_75t_SL g3571 ( 
.A(n_3474),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3427),
.Y(n_3572)
);

BUFx2_ASAP7_75t_L g3573 ( 
.A(n_3455),
.Y(n_3573)
);

HB1xp67_ASAP7_75t_L g3574 ( 
.A(n_3412),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3446),
.B(n_3403),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3447),
.B(n_3381),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3477),
.B(n_3326),
.Y(n_3577)
);

INVx3_ASAP7_75t_L g3578 ( 
.A(n_3474),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3419),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3449),
.B(n_3351),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3419),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3477),
.B(n_3518),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3518),
.B(n_3328),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3422),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3422),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3428),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3470),
.B(n_3404),
.Y(n_3587)
);

INVx2_ASAP7_75t_SL g3588 ( 
.A(n_3474),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3470),
.B(n_2978),
.Y(n_3589)
);

AND2x4_ASAP7_75t_L g3590 ( 
.A(n_3466),
.B(n_2994),
.Y(n_3590)
);

INVxp67_ASAP7_75t_L g3591 ( 
.A(n_3512),
.Y(n_3591)
);

NOR2x1_ASAP7_75t_SL g3592 ( 
.A(n_3490),
.B(n_3491),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3412),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3428),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3427),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3466),
.B(n_2995),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3412),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3435),
.B(n_3310),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3493),
.B(n_3100),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3493),
.B(n_3491),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3432),
.Y(n_3601)
);

OR2x2_ASAP7_75t_L g3602 ( 
.A(n_3461),
.B(n_2984),
.Y(n_3602)
);

OR2x2_ASAP7_75t_L g3603 ( 
.A(n_3461),
.B(n_2984),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3407),
.B(n_3303),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3517),
.B(n_3179),
.Y(n_3605)
);

INVxp67_ASAP7_75t_SL g3606 ( 
.A(n_3415),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3425),
.B(n_3100),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_R g3608 ( 
.A(n_3514),
.B(n_3281),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3432),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3457),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3425),
.B(n_3220),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3455),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3440),
.Y(n_3613)
);

INVxp67_ASAP7_75t_SL g3614 ( 
.A(n_3512),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3440),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3487),
.B(n_3078),
.Y(n_3616)
);

OR2x2_ASAP7_75t_L g3617 ( 
.A(n_3505),
.B(n_2961),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3424),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3457),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3440),
.Y(n_3620)
);

HB1xp67_ASAP7_75t_L g3621 ( 
.A(n_3416),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3526),
.B(n_3220),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3487),
.B(n_3250),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3515),
.B(n_2957),
.Y(n_3624)
);

INVx4_ASAP7_75t_L g3625 ( 
.A(n_3514),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3515),
.B(n_2957),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3517),
.B(n_3179),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3416),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3489),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3505),
.B(n_3078),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3516),
.B(n_3164),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3516),
.B(n_3519),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3448),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3519),
.B(n_3224),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3416),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3409),
.Y(n_3636)
);

NOR2xp67_ASAP7_75t_L g3637 ( 
.A(n_3494),
.B(n_3512),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3448),
.Y(n_3638)
);

INVx3_ASAP7_75t_L g3639 ( 
.A(n_3414),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3452),
.B(n_3184),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3452),
.B(n_3184),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3531),
.B(n_3320),
.Y(n_3642)
);

BUFx3_ASAP7_75t_L g3643 ( 
.A(n_3514),
.Y(n_3643)
);

AND2x4_ASAP7_75t_L g3644 ( 
.A(n_3424),
.B(n_3082),
.Y(n_3644)
);

INVx4_ASAP7_75t_L g3645 ( 
.A(n_3512),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3531),
.B(n_3227),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3490),
.B(n_3227),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_SL g3648 ( 
.A(n_3481),
.B(n_3241),
.Y(n_3648)
);

HB1xp67_ASAP7_75t_L g3649 ( 
.A(n_3414),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3643),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3643),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_3645),
.Y(n_3652)
);

INVx3_ASAP7_75t_L g3653 ( 
.A(n_3645),
.Y(n_3653)
);

NAND2x1p5_ASAP7_75t_L g3654 ( 
.A(n_3554),
.B(n_3494),
.Y(n_3654)
);

INVx1_ASAP7_75t_SL g3655 ( 
.A(n_3573),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3540),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3543),
.B(n_3410),
.Y(n_3657)
);

OR2x2_ASAP7_75t_L g3658 ( 
.A(n_3567),
.B(n_3410),
.Y(n_3658)
);

AND2x4_ASAP7_75t_L g3659 ( 
.A(n_3548),
.B(n_3478),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_L g3660 ( 
.A1(n_3538),
.A2(n_3533),
.B1(n_3520),
.B2(n_3499),
.Y(n_3660)
);

OR2x2_ASAP7_75t_L g3661 ( 
.A(n_3618),
.B(n_3471),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3550),
.Y(n_3662)
);

OR2x6_ASAP7_75t_L g3663 ( 
.A(n_3637),
.B(n_3494),
.Y(n_3663)
);

OR2x6_ASAP7_75t_SL g3664 ( 
.A(n_3598),
.B(n_3467),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3573),
.B(n_3612),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3612),
.B(n_3478),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3618),
.B(n_3499),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3592),
.B(n_3475),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3639),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3592),
.B(n_3475),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3539),
.B(n_3433),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3582),
.B(n_3476),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3550),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3563),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3563),
.Y(n_3675)
);

INVx4_ASAP7_75t_L g3676 ( 
.A(n_3548),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3582),
.B(n_3413),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3579),
.Y(n_3678)
);

OR2x6_ASAP7_75t_L g3679 ( 
.A(n_3645),
.B(n_3414),
.Y(n_3679)
);

AND2x4_ASAP7_75t_SL g3680 ( 
.A(n_3649),
.B(n_3413),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3579),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3581),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3556),
.B(n_3421),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3587),
.B(n_3476),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3581),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3584),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3556),
.B(n_3421),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3546),
.B(n_3469),
.Y(n_3688)
);

AND2x4_ASAP7_75t_L g3689 ( 
.A(n_3548),
.B(n_3639),
.Y(n_3689)
);

BUFx3_ASAP7_75t_L g3690 ( 
.A(n_3639),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3587),
.B(n_3469),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3584),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3551),
.B(n_3490),
.Y(n_3693)
);

HB1xp67_ASAP7_75t_L g3694 ( 
.A(n_3574),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3585),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3585),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3586),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3551),
.B(n_3490),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3614),
.B(n_3525),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3566),
.B(n_3482),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3586),
.Y(n_3701)
);

AND2x4_ASAP7_75t_L g3702 ( 
.A(n_3548),
.B(n_3506),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3549),
.B(n_3490),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3542),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3566),
.B(n_3489),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3549),
.B(n_3506),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3557),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3558),
.Y(n_3708)
);

INVx1_ASAP7_75t_SL g3709 ( 
.A(n_3608),
.Y(n_3709)
);

OR2x2_ASAP7_75t_L g3710 ( 
.A(n_3534),
.B(n_3471),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3625),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3600),
.B(n_3521),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3600),
.B(n_3521),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3591),
.B(n_3483),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_SL g3715 ( 
.A(n_3625),
.B(n_3463),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3606),
.B(n_3530),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3575),
.B(n_3483),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3560),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3583),
.B(n_3530),
.Y(n_3719)
);

OR2x2_ASAP7_75t_L g3720 ( 
.A(n_3534),
.B(n_3472),
.Y(n_3720)
);

INVx4_ASAP7_75t_L g3721 ( 
.A(n_3548),
.Y(n_3721)
);

INVxp67_ASAP7_75t_SL g3722 ( 
.A(n_3554),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3583),
.B(n_3462),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3594),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3601),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_SL g3726 ( 
.A(n_3640),
.B(n_3513),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3575),
.B(n_3462),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3535),
.B(n_3441),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3544),
.B(n_3426),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_3577),
.B(n_3462),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3577),
.B(n_3441),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3632),
.B(n_3492),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3632),
.B(n_3492),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3578),
.B(n_3492),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3642),
.B(n_3498),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3642),
.B(n_3498),
.Y(n_3736)
);

INVxp67_ASAP7_75t_SL g3737 ( 
.A(n_3578),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3625),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3571),
.B(n_3441),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3599),
.B(n_3409),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3571),
.B(n_3458),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3599),
.B(n_3417),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3666),
.B(n_3578),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3694),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3666),
.B(n_3588),
.Y(n_3745)
);

OR2x2_ASAP7_75t_L g3746 ( 
.A(n_3655),
.B(n_3537),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3667),
.B(n_3588),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3665),
.Y(n_3748)
);

INVxp67_ASAP7_75t_SL g3749 ( 
.A(n_3665),
.Y(n_3749)
);

AND2x4_ASAP7_75t_L g3750 ( 
.A(n_3690),
.B(n_3689),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3667),
.B(n_3607),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3657),
.B(n_3537),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3730),
.B(n_3607),
.Y(n_3753)
);

AND2x6_ASAP7_75t_SL g3754 ( 
.A(n_3731),
.B(n_3604),
.Y(n_3754)
);

INVx2_ASAP7_75t_SL g3755 ( 
.A(n_3690),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3676),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3661),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3730),
.B(n_3623),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3657),
.B(n_3597),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3676),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3680),
.B(n_3623),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3661),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3710),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3676),
.Y(n_3764)
);

OR2x2_ASAP7_75t_L g3765 ( 
.A(n_3658),
.B(n_3597),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3710),
.Y(n_3766)
);

NAND4xp25_ASAP7_75t_L g3767 ( 
.A(n_3660),
.B(n_3559),
.C(n_3580),
.D(n_3564),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3720),
.Y(n_3768)
);

OR2x2_ASAP7_75t_L g3769 ( 
.A(n_3658),
.B(n_3656),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3680),
.B(n_3622),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3727),
.B(n_3629),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3721),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3727),
.B(n_3622),
.Y(n_3773)
);

INVxp67_ASAP7_75t_SL g3774 ( 
.A(n_3654),
.Y(n_3774)
);

OR2x2_ASAP7_75t_L g3775 ( 
.A(n_3699),
.B(n_3628),
.Y(n_3775)
);

NAND2x1p5_ASAP7_75t_L g3776 ( 
.A(n_3721),
.B(n_3640),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3720),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3737),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3723),
.B(n_3589),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3662),
.Y(n_3780)
);

NAND2x1_ASAP7_75t_L g3781 ( 
.A(n_3663),
.B(n_3641),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3721),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3689),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3689),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3723),
.B(n_3589),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3650),
.B(n_3641),
.Y(n_3786)
);

AND2x4_ASAP7_75t_L g3787 ( 
.A(n_3659),
.B(n_3652),
.Y(n_3787)
);

OR2x2_ASAP7_75t_L g3788 ( 
.A(n_3728),
.B(n_3628),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3722),
.B(n_3552),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3659),
.B(n_3552),
.Y(n_3790)
);

NOR3xp33_ASAP7_75t_L g3791 ( 
.A(n_3726),
.B(n_3576),
.C(n_3553),
.Y(n_3791)
);

NOR2x1_ASAP7_75t_SL g3792 ( 
.A(n_3663),
.B(n_3535),
.Y(n_3792)
);

INVxp67_ASAP7_75t_SL g3793 ( 
.A(n_3654),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3659),
.B(n_3555),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3652),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3716),
.B(n_3703),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3716),
.B(n_3555),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3703),
.B(n_3562),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3673),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3684),
.B(n_3562),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3684),
.B(n_3565),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3674),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3675),
.Y(n_3803)
);

AND2x4_ASAP7_75t_L g3804 ( 
.A(n_3652),
.B(n_3565),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3672),
.B(n_3569),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3672),
.B(n_3569),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3693),
.B(n_3570),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3650),
.B(n_3547),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3678),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3651),
.B(n_3536),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3651),
.B(n_3536),
.Y(n_3811)
);

AND2x4_ASAP7_75t_L g3812 ( 
.A(n_3653),
.B(n_3570),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3693),
.B(n_3572),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3681),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3698),
.B(n_3572),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3698),
.B(n_3595),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3719),
.B(n_3595),
.Y(n_3817)
);

BUFx2_ASAP7_75t_L g3818 ( 
.A(n_3679),
.Y(n_3818)
);

OR2x2_ASAP7_75t_L g3819 ( 
.A(n_3705),
.B(n_3635),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3706),
.B(n_3719),
.Y(n_3820)
);

NAND2xp33_ASAP7_75t_R g3821 ( 
.A(n_3663),
.B(n_3524),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3726),
.A2(n_3561),
.B(n_3648),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3669),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3732),
.B(n_3646),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3732),
.B(n_3646),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3682),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3653),
.Y(n_3827)
);

HB1xp67_ASAP7_75t_L g3828 ( 
.A(n_3669),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3653),
.Y(n_3829)
);

OR2x2_ASAP7_75t_L g3830 ( 
.A(n_3739),
.B(n_3717),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3679),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3685),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_3715),
.B(n_3611),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3733),
.B(n_3611),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3733),
.B(n_3647),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3759),
.Y(n_3836)
);

HB1xp67_ASAP7_75t_L g3837 ( 
.A(n_3823),
.Y(n_3837)
);

AND2x2_ASAP7_75t_SL g3838 ( 
.A(n_3791),
.B(n_3729),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3796),
.B(n_3709),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3759),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3765),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3747),
.B(n_3706),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3765),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3796),
.B(n_3712),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3747),
.B(n_3711),
.Y(n_3845)
);

INVxp67_ASAP7_75t_L g3846 ( 
.A(n_3792),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3743),
.B(n_3668),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3743),
.B(n_3668),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3773),
.B(n_3670),
.Y(n_3849)
);

OAI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3822),
.A2(n_3833),
.B(n_3793),
.Y(n_3850)
);

NAND3xp33_ASAP7_75t_L g3851 ( 
.A(n_3821),
.B(n_3687),
.C(n_3683),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3773),
.B(n_3670),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3752),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3752),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3758),
.B(n_3712),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3749),
.B(n_3711),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3758),
.B(n_3713),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3755),
.B(n_3738),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3776),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3757),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3757),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3776),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3776),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3762),
.Y(n_3864)
);

INVx2_ASAP7_75t_SL g3865 ( 
.A(n_3787),
.Y(n_3865)
);

INVx1_ASAP7_75t_SL g3866 ( 
.A(n_3770),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3755),
.B(n_3738),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3762),
.Y(n_3868)
);

NAND4xp25_ASAP7_75t_L g3869 ( 
.A(n_3767),
.B(n_3677),
.C(n_3671),
.D(n_3700),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3770),
.B(n_3664),
.Y(n_3870)
);

NAND2x1p5_ASAP7_75t_L g3871 ( 
.A(n_3781),
.B(n_3702),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3824),
.B(n_3713),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3828),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3748),
.B(n_3664),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3792),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3824),
.B(n_3735),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3748),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3825),
.B(n_3735),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3825),
.B(n_3736),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3787),
.Y(n_3880)
);

INVx1_ASAP7_75t_SL g3881 ( 
.A(n_3761),
.Y(n_3881)
);

OR2x2_ASAP7_75t_L g3882 ( 
.A(n_3820),
.B(n_3741),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3789),
.B(n_3714),
.Y(n_3883)
);

HB1xp67_ASAP7_75t_L g3884 ( 
.A(n_3797),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3787),
.B(n_3679),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3778),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3789),
.B(n_3736),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3778),
.Y(n_3888)
);

NAND2x2_ASAP7_75t_L g3889 ( 
.A(n_3808),
.B(n_3830),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3834),
.B(n_3691),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3786),
.B(n_3688),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3761),
.B(n_3740),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3746),
.B(n_3605),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3763),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3834),
.B(n_3734),
.Y(n_3895)
);

BUFx3_ASAP7_75t_L g3896 ( 
.A(n_3750),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3835),
.B(n_3751),
.Y(n_3897)
);

INVx3_ASAP7_75t_L g3898 ( 
.A(n_3787),
.Y(n_3898)
);

OR2x2_ASAP7_75t_L g3899 ( 
.A(n_3746),
.B(n_3627),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3835),
.B(n_3734),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3797),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3750),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3751),
.B(n_3734),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3763),
.Y(n_3904)
);

INVxp67_ASAP7_75t_L g3905 ( 
.A(n_3750),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3754),
.B(n_3663),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3779),
.B(n_3740),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3750),
.B(n_3679),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3766),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3766),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3753),
.B(n_3742),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3779),
.B(n_3742),
.Y(n_3912)
);

HB1xp67_ASAP7_75t_L g3913 ( 
.A(n_3768),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3769),
.B(n_3636),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3768),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3781),
.Y(n_3916)
);

AND2x4_ASAP7_75t_L g3917 ( 
.A(n_3783),
.B(n_3784),
.Y(n_3917)
);

NOR2xp33_ASAP7_75t_L g3918 ( 
.A(n_3769),
.B(n_3702),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3777),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3753),
.B(n_3702),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3777),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3788),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3798),
.B(n_3704),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3788),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3785),
.B(n_3647),
.Y(n_3925)
);

OAI22xp5_ASAP7_75t_L g3926 ( 
.A1(n_3838),
.A2(n_3774),
.B1(n_3830),
.B2(n_3524),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3839),
.B(n_3798),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3892),
.B(n_3807),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3865),
.B(n_3783),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3838),
.B(n_3745),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3913),
.Y(n_3931)
);

BUFx2_ASAP7_75t_SL g3932 ( 
.A(n_3865),
.Y(n_3932)
);

OR2x2_ASAP7_75t_L g3933 ( 
.A(n_3897),
.B(n_3810),
.Y(n_3933)
);

OAI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3906),
.A2(n_3744),
.B(n_3818),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3847),
.B(n_3784),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3892),
.B(n_3807),
.Y(n_3936)
);

OR2x6_ASAP7_75t_L g3937 ( 
.A(n_3875),
.B(n_3756),
.Y(n_3937)
);

INVxp67_ASAP7_75t_SL g3938 ( 
.A(n_3871),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3871),
.Y(n_3939)
);

NOR3xp33_ASAP7_75t_L g3940 ( 
.A(n_3906),
.B(n_3811),
.C(n_3818),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3887),
.B(n_3771),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3898),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3847),
.B(n_3790),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3913),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3876),
.B(n_3813),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3896),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3837),
.Y(n_3947)
);

NAND2x2_ASAP7_75t_L g3948 ( 
.A(n_3896),
.B(n_3775),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3898),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3876),
.B(n_3855),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3848),
.B(n_3790),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3837),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3884),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3898),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3846),
.A2(n_3744),
.B(n_3775),
.Y(n_3955)
);

INVxp33_ASAP7_75t_L g3956 ( 
.A(n_3870),
.Y(n_3956)
);

OAI21xp33_ASAP7_75t_L g3957 ( 
.A1(n_3850),
.A2(n_3815),
.B(n_3813),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3866),
.B(n_3819),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3884),
.B(n_3901),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3848),
.B(n_3794),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3855),
.B(n_3815),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3901),
.Y(n_3962)
);

OR2x2_ASAP7_75t_L g3963 ( 
.A(n_3911),
.B(n_3819),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3857),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3857),
.Y(n_3965)
);

INVxp67_ASAP7_75t_L g3966 ( 
.A(n_3918),
.Y(n_3966)
);

INVx3_ASAP7_75t_L g3967 ( 
.A(n_3885),
.Y(n_3967)
);

OAI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3889),
.A2(n_3524),
.B1(n_3496),
.B2(n_3831),
.Y(n_3968)
);

OAI22xp5_ASAP7_75t_L g3969 ( 
.A1(n_3889),
.A2(n_3524),
.B1(n_3496),
.B2(n_3831),
.Y(n_3969)
);

OR2x2_ASAP7_75t_L g3970 ( 
.A(n_3842),
.B(n_3800),
.Y(n_3970)
);

NOR2xp33_ASAP7_75t_L g3971 ( 
.A(n_3869),
.B(n_3756),
.Y(n_3971)
);

OR2x2_ASAP7_75t_L g3972 ( 
.A(n_3881),
.B(n_3800),
.Y(n_3972)
);

NOR3x1_ASAP7_75t_L g3973 ( 
.A(n_3851),
.B(n_3799),
.C(n_3780),
.Y(n_3973)
);

AOI32xp33_ASAP7_75t_L g3974 ( 
.A1(n_3875),
.A2(n_3852),
.A3(n_3849),
.B1(n_3874),
.B2(n_3907),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3917),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3880),
.Y(n_3976)
);

OR4x1_ASAP7_75t_L g3977 ( 
.A(n_3853),
.B(n_3799),
.C(n_3802),
.D(n_3780),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3917),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3907),
.B(n_3912),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3849),
.B(n_3794),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3917),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3912),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3878),
.A2(n_3496),
.B1(n_3497),
.B2(n_3785),
.Y(n_3983)
);

INVxp67_ASAP7_75t_SL g3984 ( 
.A(n_3918),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3872),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_L g3986 ( 
.A(n_3883),
.B(n_3760),
.Y(n_3986)
);

INVxp67_ASAP7_75t_L g3987 ( 
.A(n_3852),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3879),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3844),
.B(n_3925),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3916),
.Y(n_3990)
);

NOR3xp33_ASAP7_75t_L g3991 ( 
.A(n_3856),
.B(n_3764),
.C(n_3760),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3895),
.B(n_3801),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3914),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3854),
.Y(n_3994)
);

OR2x2_ASAP7_75t_L g3995 ( 
.A(n_3900),
.B(n_3801),
.Y(n_3995)
);

INVxp67_ASAP7_75t_L g3996 ( 
.A(n_3908),
.Y(n_3996)
);

OR2x2_ASAP7_75t_L g3997 ( 
.A(n_3893),
.B(n_3817),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3905),
.B(n_3816),
.Y(n_3998)
);

AND2x4_ASAP7_75t_SL g3999 ( 
.A(n_3908),
.B(n_3885),
.Y(n_3999)
);

INVxp67_ASAP7_75t_L g4000 ( 
.A(n_3908),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3902),
.B(n_3880),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3922),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3924),
.Y(n_4003)
);

INVx1_ASAP7_75t_SL g4004 ( 
.A(n_3885),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3836),
.B(n_3795),
.Y(n_4005)
);

AOI32xp33_ASAP7_75t_L g4006 ( 
.A1(n_3916),
.A2(n_3816),
.A3(n_3920),
.B1(n_3873),
.B2(n_3817),
.Y(n_4006)
);

AO221x1_ASAP7_75t_L g4007 ( 
.A1(n_3902),
.A2(n_3829),
.B1(n_3827),
.B2(n_3795),
.C(n_3764),
.Y(n_4007)
);

OAI32xp33_ASAP7_75t_L g4008 ( 
.A1(n_3899),
.A2(n_3829),
.A3(n_3827),
.B1(n_3772),
.B2(n_3782),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3903),
.B(n_3805),
.Y(n_4009)
);

OAI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3926),
.A2(n_3496),
.B1(n_3845),
.B2(n_3890),
.Y(n_4010)
);

INVxp67_ASAP7_75t_L g4011 ( 
.A(n_3932),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3930),
.A2(n_3926),
.B(n_3934),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3954),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3959),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3959),
.Y(n_4015)
);

OAI31xp33_ASAP7_75t_L g4016 ( 
.A1(n_3968),
.A2(n_3841),
.A3(n_3843),
.B(n_3840),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_SL g4017 ( 
.A1(n_4007),
.A2(n_3561),
.B1(n_3806),
.B2(n_3805),
.Y(n_4017)
);

INVxp67_ASAP7_75t_L g4018 ( 
.A(n_3938),
.Y(n_4018)
);

INVx4_ASAP7_75t_L g4019 ( 
.A(n_3967),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3927),
.B(n_3859),
.Y(n_4020)
);

INVx1_ASAP7_75t_SL g4021 ( 
.A(n_4004),
.Y(n_4021)
);

AOI22xp5_ASAP7_75t_L g4022 ( 
.A1(n_3957),
.A2(n_3806),
.B1(n_3812),
.B2(n_3858),
.Y(n_4022)
);

A2O1A1Ixp33_ASAP7_75t_L g4023 ( 
.A1(n_3934),
.A2(n_3862),
.B(n_3863),
.C(n_3859),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3975),
.Y(n_4024)
);

OAI21xp33_ASAP7_75t_SL g4025 ( 
.A1(n_3983),
.A2(n_3863),
.B(n_3862),
.Y(n_4025)
);

INVx2_ASAP7_75t_SL g4026 ( 
.A(n_3929),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3928),
.B(n_3882),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3978),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3981),
.Y(n_4029)
);

INVx2_ASAP7_75t_SL g4030 ( 
.A(n_3929),
.Y(n_4030)
);

AOI21xp33_ASAP7_75t_L g4031 ( 
.A1(n_3956),
.A2(n_3891),
.B(n_3867),
.Y(n_4031)
);

AOI21xp33_ASAP7_75t_L g4032 ( 
.A1(n_3984),
.A2(n_3923),
.B(n_3888),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3931),
.Y(n_4033)
);

O2A1O1Ixp33_ASAP7_75t_L g4034 ( 
.A1(n_3955),
.A2(n_3861),
.B(n_3864),
.C(n_3860),
.Y(n_4034)
);

XOR2x2_ASAP7_75t_L g4035 ( 
.A(n_3989),
.B(n_3886),
.Y(n_4035)
);

OAI21xp33_ASAP7_75t_L g4036 ( 
.A1(n_3957),
.A2(n_3877),
.B(n_3868),
.Y(n_4036)
);

OAI22xp33_ASAP7_75t_L g4037 ( 
.A1(n_3948),
.A2(n_3972),
.B1(n_3997),
.B2(n_4004),
.Y(n_4037)
);

INVx2_ASAP7_75t_SL g4038 ( 
.A(n_3999),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3944),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3990),
.Y(n_4040)
);

NOR2xp33_ASAP7_75t_L g4041 ( 
.A(n_3996),
.B(n_4000),
.Y(n_4041)
);

INVxp67_ASAP7_75t_L g4042 ( 
.A(n_3936),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3942),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_SL g4044 ( 
.A1(n_3974),
.A2(n_3921),
.B(n_3904),
.Y(n_4044)
);

INVxp67_ASAP7_75t_L g4045 ( 
.A(n_3961),
.Y(n_4045)
);

AOI22x1_ASAP7_75t_L g4046 ( 
.A1(n_3939),
.A2(n_3772),
.B1(n_3782),
.B2(n_3910),
.Y(n_4046)
);

NAND3xp33_ASAP7_75t_L g4047 ( 
.A(n_3940),
.B(n_3909),
.C(n_3894),
.Y(n_4047)
);

AOI31xp33_ASAP7_75t_L g4048 ( 
.A1(n_3987),
.A2(n_3919),
.A3(n_3915),
.B(n_3832),
.Y(n_4048)
);

AOI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3945),
.A2(n_3812),
.B1(n_3804),
.B2(n_3468),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3949),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3950),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3967),
.Y(n_4052)
);

NOR2xp33_ASAP7_75t_L g4053 ( 
.A(n_3966),
.B(n_3802),
.Y(n_4053)
);

AOI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3979),
.A2(n_3812),
.B1(n_3804),
.B2(n_3636),
.Y(n_4054)
);

A2O1A1Ixp33_ASAP7_75t_L g4055 ( 
.A1(n_3955),
.A2(n_3832),
.B(n_3826),
.C(n_3814),
.Y(n_4055)
);

OAI21xp33_ASAP7_75t_L g4056 ( 
.A1(n_3971),
.A2(n_3804),
.B(n_3708),
.Y(n_4056)
);

INVx2_ASAP7_75t_SL g4057 ( 
.A(n_3946),
.Y(n_4057)
);

XOR2x2_ASAP7_75t_L g4058 ( 
.A(n_3980),
.B(n_3509),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3953),
.Y(n_4059)
);

OAI22xp5_ASAP7_75t_L g4060 ( 
.A1(n_3943),
.A2(n_3960),
.B1(n_3951),
.B2(n_3933),
.Y(n_4060)
);

O2A1O1Ixp5_ASAP7_75t_L g4061 ( 
.A1(n_3968),
.A2(n_3804),
.B(n_3814),
.C(n_3809),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3962),
.Y(n_4062)
);

XNOR2xp5_ASAP7_75t_L g4063 ( 
.A(n_4009),
.B(n_3707),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3976),
.Y(n_4064)
);

OAI211xp5_ASAP7_75t_L g4065 ( 
.A1(n_4006),
.A2(n_3826),
.B(n_3809),
.C(n_3803),
.Y(n_4065)
);

OAI21xp5_ASAP7_75t_SL g4066 ( 
.A1(n_3969),
.A2(n_3803),
.B(n_3724),
.Y(n_4066)
);

OAI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_3969),
.A2(n_3725),
.B(n_3718),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3982),
.B(n_3593),
.Y(n_4068)
);

OAI21xp33_ASAP7_75t_L g4069 ( 
.A1(n_3988),
.A2(n_3692),
.B(n_3686),
.Y(n_4069)
);

OAI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3986),
.A2(n_3621),
.B(n_3695),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3992),
.A2(n_3502),
.B1(n_3528),
.B2(n_3437),
.Y(n_4071)
);

AOI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3985),
.A2(n_3631),
.B1(n_3610),
.B2(n_3619),
.Y(n_4072)
);

AOI21xp33_ASAP7_75t_L g4073 ( 
.A1(n_3958),
.A2(n_3635),
.B(n_3696),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3937),
.A2(n_3998),
.B(n_4005),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_4026),
.B(n_3964),
.Y(n_4075)
);

INVx1_ASAP7_75t_SL g4076 ( 
.A(n_4021),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_4030),
.Y(n_4077)
);

AOI222xp33_ASAP7_75t_L g4078 ( 
.A1(n_4047),
.A2(n_3952),
.B1(n_3947),
.B2(n_4003),
.C1(n_4002),
.C2(n_3994),
.Y(n_4078)
);

AOI21xp33_ASAP7_75t_L g4079 ( 
.A1(n_4037),
.A2(n_3993),
.B(n_3963),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_4019),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4019),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_4038),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_4052),
.B(n_3965),
.Y(n_4083)
);

AOI222xp33_ASAP7_75t_L g4084 ( 
.A1(n_4047),
.A2(n_4005),
.B1(n_4008),
.B2(n_4001),
.C1(n_3935),
.C2(n_3973),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4051),
.Y(n_4085)
);

OAI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_4012),
.A2(n_3995),
.B1(n_3970),
.B2(n_3937),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_4011),
.B(n_3941),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_4020),
.Y(n_4088)
);

OAI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_4017),
.A2(n_3937),
.B1(n_3502),
.B2(n_3436),
.Y(n_4089)
);

OAI22xp5_ASAP7_75t_L g4090 ( 
.A1(n_4049),
.A2(n_3437),
.B1(n_3436),
.B2(n_3431),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4027),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4041),
.Y(n_4092)
);

OAI32xp33_ASAP7_75t_L g4093 ( 
.A1(n_4025),
.A2(n_3991),
.A3(n_3701),
.B1(n_3697),
.B2(n_3977),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_4057),
.B(n_3631),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4022),
.B(n_3609),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4013),
.Y(n_4096)
);

XNOR2xp5_ASAP7_75t_L g4097 ( 
.A(n_4058),
.B(n_4035),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4040),
.Y(n_4098)
);

AOI222xp33_ASAP7_75t_L g4099 ( 
.A1(n_4036),
.A2(n_3613),
.B1(n_3638),
.B2(n_3633),
.C1(n_3615),
.C2(n_3620),
.Y(n_4099)
);

AO22x1_ASAP7_75t_L g4100 ( 
.A1(n_4014),
.A2(n_3644),
.B1(n_3590),
.B2(n_3596),
.Y(n_4100)
);

AOI211xp5_ASAP7_75t_L g4101 ( 
.A1(n_4010),
.A2(n_3644),
.B(n_3634),
.C(n_3638),
.Y(n_4101)
);

NAND2xp33_ASAP7_75t_R g4102 ( 
.A(n_4015),
.B(n_315),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_4074),
.B(n_3442),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4063),
.Y(n_4104)
);

AOI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_4042),
.A2(n_3644),
.B1(n_3430),
.B2(n_3431),
.Y(n_4105)
);

OAI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_4044),
.A2(n_3568),
.B1(n_3430),
.B2(n_3633),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4068),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_4046),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_4024),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_SL g4110 ( 
.A1(n_4065),
.A2(n_3634),
.B1(n_3429),
.B2(n_3434),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4018),
.B(n_3442),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_4028),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4029),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4045),
.B(n_3456),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4043),
.Y(n_4115)
);

AOI221xp5_ASAP7_75t_L g4116 ( 
.A1(n_4031),
.A2(n_3620),
.B1(n_3613),
.B2(n_3615),
.C(n_3472),
.Y(n_4116)
);

OAI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_4054),
.A2(n_3290),
.B1(n_3568),
.B2(n_3339),
.Y(n_4117)
);

OAI22xp33_ASAP7_75t_SL g4118 ( 
.A1(n_4050),
.A2(n_4059),
.B1(n_4062),
.B2(n_4064),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_4056),
.B(n_3454),
.Y(n_4119)
);

AOI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_4060),
.A2(n_3438),
.B1(n_3590),
.B2(n_3596),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_4023),
.B(n_3456),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4048),
.Y(n_4122)
);

INVxp67_ASAP7_75t_L g4123 ( 
.A(n_4053),
.Y(n_4123)
);

OAI221xp5_ASAP7_75t_SL g4124 ( 
.A1(n_4016),
.A2(n_3568),
.B1(n_3541),
.B2(n_3438),
.C(n_3434),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_4070),
.B(n_3454),
.Y(n_4125)
);

OAI32xp33_ASAP7_75t_L g4126 ( 
.A1(n_4033),
.A2(n_4039),
.A3(n_4032),
.B1(n_4071),
.B2(n_4067),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4034),
.Y(n_4127)
);

AOI221xp5_ASAP7_75t_L g4128 ( 
.A1(n_4016),
.A2(n_3590),
.B1(n_3596),
.B2(n_3616),
.C(n_3473),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_4061),
.Y(n_4129)
);

INVx1_ASAP7_75t_SL g4130 ( 
.A(n_4073),
.Y(n_4130)
);

OAI32xp33_ASAP7_75t_L g4131 ( 
.A1(n_4069),
.A2(n_3382),
.A3(n_3541),
.B1(n_3429),
.B2(n_3630),
.Y(n_4131)
);

NOR2x1_ASAP7_75t_L g4132 ( 
.A(n_4066),
.B(n_3616),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_4072),
.B(n_3616),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4055),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4066),
.B(n_3479),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4082),
.B(n_3479),
.Y(n_4136)
);

AOI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_4076),
.A2(n_3568),
.B1(n_3293),
.B2(n_3292),
.Y(n_4137)
);

OR2x2_ASAP7_75t_L g4138 ( 
.A(n_4076),
.B(n_4075),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4077),
.B(n_3484),
.Y(n_4139)
);

INVxp67_ASAP7_75t_L g4140 ( 
.A(n_4102),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4091),
.B(n_3484),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_L g4142 ( 
.A(n_4081),
.B(n_3545),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4125),
.B(n_3624),
.Y(n_4143)
);

HB1xp67_ASAP7_75t_L g4144 ( 
.A(n_4129),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4094),
.Y(n_4145)
);

OAI221xp5_ASAP7_75t_L g4146 ( 
.A1(n_4127),
.A2(n_3545),
.B1(n_3297),
.B2(n_3473),
.C(n_3485),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_4080),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4083),
.Y(n_4148)
);

AO22x1_ASAP7_75t_L g4149 ( 
.A1(n_4134),
.A2(n_3507),
.B1(n_3504),
.B2(n_3503),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_4132),
.Y(n_4150)
);

HB1xp67_ASAP7_75t_L g4151 ( 
.A(n_4122),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4119),
.B(n_3624),
.Y(n_4152)
);

OAI32xp33_ASAP7_75t_L g4153 ( 
.A1(n_4108),
.A2(n_3630),
.A3(n_3417),
.B1(n_3465),
.B2(n_3464),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4085),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4088),
.B(n_3626),
.Y(n_4155)
);

AOI21xp33_ASAP7_75t_L g4156 ( 
.A1(n_4086),
.A2(n_3603),
.B(n_3602),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4096),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4092),
.B(n_3626),
.Y(n_4158)
);

AOI22xp33_ASAP7_75t_L g4159 ( 
.A1(n_4079),
.A2(n_3485),
.B1(n_3465),
.B2(n_3464),
.Y(n_4159)
);

OAI21xp33_ASAP7_75t_SL g4160 ( 
.A1(n_4084),
.A2(n_3603),
.B(n_3602),
.Y(n_4160)
);

INVx1_ASAP7_75t_SL g4161 ( 
.A(n_4130),
.Y(n_4161)
);

INVx2_ASAP7_75t_SL g4162 ( 
.A(n_4100),
.Y(n_4162)
);

AOI322xp5_ASAP7_75t_L g4163 ( 
.A1(n_4130),
.A2(n_3503),
.A3(n_3504),
.B1(n_3453),
.B2(n_3445),
.C1(n_3507),
.C2(n_3480),
.Y(n_4163)
);

AOI32xp33_ASAP7_75t_L g4164 ( 
.A1(n_4089),
.A2(n_3453),
.A3(n_3445),
.B1(n_3480),
.B2(n_3529),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4087),
.Y(n_4165)
);

XNOR2x1_ASAP7_75t_L g4166 ( 
.A(n_4097),
.B(n_316),
.Y(n_4166)
);

NAND2xp33_ASAP7_75t_L g4167 ( 
.A(n_4109),
.B(n_3617),
.Y(n_4167)
);

OAI21xp5_ASAP7_75t_SL g4168 ( 
.A1(n_4084),
.A2(n_3480),
.B(n_3501),
.Y(n_4168)
);

INVxp67_ASAP7_75t_L g4169 ( 
.A(n_4078),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4098),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_4093),
.A2(n_4126),
.B(n_4106),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4112),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4135),
.B(n_3480),
.Y(n_4173)
);

OAI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_4110),
.A2(n_3617),
.B1(n_3423),
.B2(n_3450),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_4106),
.A2(n_4078),
.B1(n_4121),
.B2(n_4104),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4113),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_4101),
.B(n_3423),
.Y(n_4177)
);

OAI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_4103),
.A2(n_3423),
.B1(n_3450),
.B2(n_3448),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4123),
.B(n_3488),
.Y(n_4179)
);

AOI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_4117),
.A2(n_3501),
.B1(n_3529),
.B2(n_3488),
.Y(n_4180)
);

XOR2x2_ASAP7_75t_L g4181 ( 
.A(n_4124),
.B(n_316),
.Y(n_4181)
);

INVxp67_ASAP7_75t_L g4182 ( 
.A(n_4115),
.Y(n_4182)
);

OAI21xp33_ASAP7_75t_L g4183 ( 
.A1(n_4105),
.A2(n_3450),
.B(n_3439),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4118),
.B(n_3439),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_L g4185 ( 
.A(n_4140),
.B(n_4095),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4147),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_4138),
.Y(n_4187)
);

AOI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_4169),
.A2(n_4090),
.B1(n_4107),
.B2(n_4133),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4169),
.B(n_4111),
.Y(n_4189)
);

NOR3x1_ASAP7_75t_L g4190 ( 
.A(n_4162),
.B(n_4168),
.C(n_4184),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4147),
.Y(n_4191)
);

NAND3xp33_ASAP7_75t_SL g4192 ( 
.A(n_4161),
.B(n_4114),
.C(n_4116),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_4136),
.B(n_4120),
.Y(n_4193)
);

NOR2xp67_ASAP7_75t_L g4194 ( 
.A(n_4140),
.B(n_317),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_4171),
.A2(n_4160),
.B(n_4166),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4151),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4150),
.Y(n_4197)
);

NOR3xp33_ASAP7_75t_L g4198 ( 
.A(n_4165),
.B(n_4131),
.C(n_4128),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4151),
.Y(n_4199)
);

OAI21xp33_ASAP7_75t_L g4200 ( 
.A1(n_4175),
.A2(n_4099),
.B(n_3510),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_4144),
.B(n_4099),
.Y(n_4201)
);

INVxp67_ASAP7_75t_L g4202 ( 
.A(n_4144),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4152),
.B(n_3510),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4158),
.Y(n_4204)
);

AOI221xp5_ASAP7_75t_L g4205 ( 
.A1(n_4175),
.A2(n_3204),
.B1(n_3244),
.B2(n_3243),
.C(n_3212),
.Y(n_4205)
);

NAND2xp33_ASAP7_75t_L g4206 ( 
.A(n_4139),
.B(n_3522),
.Y(n_4206)
);

BUFx2_ASAP7_75t_L g4207 ( 
.A(n_4141),
.Y(n_4207)
);

AOI21xp5_ASAP7_75t_L g4208 ( 
.A1(n_4167),
.A2(n_3522),
.B(n_3099),
.Y(n_4208)
);

AOI221x1_ASAP7_75t_L g4209 ( 
.A1(n_4157),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.C(n_321),
.Y(n_4209)
);

CKINVDCx16_ASAP7_75t_R g4210 ( 
.A(n_4145),
.Y(n_4210)
);

XNOR2x1_ASAP7_75t_L g4211 ( 
.A(n_4181),
.B(n_318),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4142),
.B(n_319),
.Y(n_4212)
);

OAI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4173),
.A2(n_3099),
.B(n_3110),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_4156),
.B(n_3110),
.Y(n_4214)
);

AOI211xp5_ASAP7_75t_L g4215 ( 
.A1(n_4146),
.A2(n_320),
.B(n_321),
.C(n_322),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_4143),
.B(n_3204),
.Y(n_4216)
);

INVx1_ASAP7_75t_SL g4217 ( 
.A(n_4179),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4155),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_4148),
.B(n_323),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_SL g4220 ( 
.A(n_4142),
.B(n_3085),
.Y(n_4220)
);

NOR3x1_ASAP7_75t_L g4221 ( 
.A(n_4172),
.B(n_4177),
.C(n_4170),
.Y(n_4221)
);

INVx2_ASAP7_75t_L g4222 ( 
.A(n_4176),
.Y(n_4222)
);

OAI221xp5_ASAP7_75t_L g4223 ( 
.A1(n_4200),
.A2(n_4159),
.B1(n_4182),
.B2(n_4154),
.C(n_4183),
.Y(n_4223)
);

NOR3xp33_ASAP7_75t_L g4224 ( 
.A(n_4210),
.B(n_4182),
.C(n_4153),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4194),
.Y(n_4225)
);

AOI21xp33_ASAP7_75t_SL g4226 ( 
.A1(n_4186),
.A2(n_4178),
.B(n_4159),
.Y(n_4226)
);

AOI211xp5_ASAP7_75t_L g4227 ( 
.A1(n_4195),
.A2(n_4178),
.B(n_4149),
.C(n_4174),
.Y(n_4227)
);

OAI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_4188),
.A2(n_4180),
.B1(n_4137),
.B2(n_4164),
.Y(n_4228)
);

NAND4xp25_ASAP7_75t_L g4229 ( 
.A(n_4190),
.B(n_4163),
.C(n_3212),
.D(n_3231),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_4191),
.B(n_3243),
.Y(n_4230)
);

NOR3x1_ASAP7_75t_L g4231 ( 
.A(n_4192),
.B(n_323),
.C(n_324),
.Y(n_4231)
);

AOI222xp33_ASAP7_75t_L g4232 ( 
.A1(n_4205),
.A2(n_3234),
.B1(n_3244),
.B2(n_3231),
.C1(n_3086),
.C2(n_3245),
.Y(n_4232)
);

AOI211xp5_ASAP7_75t_SL g4233 ( 
.A1(n_4202),
.A2(n_324),
.B(n_325),
.C(n_326),
.Y(n_4233)
);

OAI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4185),
.A2(n_2962),
.B(n_3245),
.Y(n_4234)
);

AOI221xp5_ASAP7_75t_L g4235 ( 
.A1(n_4198),
.A2(n_325),
.B1(n_327),
.B2(n_331),
.C(n_332),
.Y(n_4235)
);

AOI211x1_ASAP7_75t_L g4236 ( 
.A1(n_4201),
.A2(n_2962),
.B(n_333),
.C(n_334),
.Y(n_4236)
);

AOI21xp33_ASAP7_75t_L g4237 ( 
.A1(n_4187),
.A2(n_327),
.B(n_334),
.Y(n_4237)
);

NOR4xp25_ASAP7_75t_SL g4238 ( 
.A(n_4207),
.B(n_335),
.C(n_336),
.D(n_337),
.Y(n_4238)
);

OAI221xp5_ASAP7_75t_L g4239 ( 
.A1(n_4197),
.A2(n_3072),
.B1(n_3089),
.B2(n_3046),
.C(n_3043),
.Y(n_4239)
);

NOR3xp33_ASAP7_75t_L g4240 ( 
.A(n_4204),
.B(n_335),
.C(n_336),
.Y(n_4240)
);

OAI21xp33_ASAP7_75t_SL g4241 ( 
.A1(n_4201),
.A2(n_3015),
.B(n_3043),
.Y(n_4241)
);

OAI21xp33_ASAP7_75t_L g4242 ( 
.A1(n_4211),
.A2(n_3096),
.B(n_3082),
.Y(n_4242)
);

AOI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4217),
.A2(n_3096),
.B1(n_3008),
.B2(n_3015),
.Y(n_4243)
);

OAI211xp5_ASAP7_75t_L g4244 ( 
.A1(n_4215),
.A2(n_337),
.B(n_338),
.C(n_339),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_4214),
.A2(n_3008),
.B(n_340),
.Y(n_4245)
);

AOI221xp5_ASAP7_75t_L g4246 ( 
.A1(n_4196),
.A2(n_338),
.B1(n_341),
.B2(n_343),
.C(n_345),
.Y(n_4246)
);

OAI221xp5_ASAP7_75t_SL g4247 ( 
.A1(n_4235),
.A2(n_4199),
.B1(n_4218),
.B2(n_4189),
.C(n_4222),
.Y(n_4247)
);

OAI211xp5_ASAP7_75t_L g4248 ( 
.A1(n_4227),
.A2(n_4189),
.B(n_4212),
.C(n_4209),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_4233),
.B(n_4193),
.Y(n_4249)
);

O2A1O1Ixp5_ASAP7_75t_SL g4250 ( 
.A1(n_4225),
.A2(n_4212),
.B(n_4216),
.C(n_4221),
.Y(n_4250)
);

AOI22xp33_ASAP7_75t_L g4251 ( 
.A1(n_4224),
.A2(n_4205),
.B1(n_4206),
.B2(n_4203),
.Y(n_4251)
);

AOI22xp5_ASAP7_75t_L g4252 ( 
.A1(n_4228),
.A2(n_4203),
.B1(n_4219),
.B2(n_4220),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4231),
.Y(n_4253)
);

OAI22xp5_ASAP7_75t_L g4254 ( 
.A1(n_4223),
.A2(n_4208),
.B1(n_4213),
.B2(n_3046),
.Y(n_4254)
);

AOI221xp5_ASAP7_75t_L g4255 ( 
.A1(n_4226),
.A2(n_4229),
.B1(n_4236),
.B2(n_4242),
.C(n_4230),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4244),
.Y(n_4256)
);

OAI21xp5_ASAP7_75t_SL g4257 ( 
.A1(n_4245),
.A2(n_343),
.B(n_345),
.Y(n_4257)
);

OAI211xp5_ASAP7_75t_SL g4258 ( 
.A1(n_4241),
.A2(n_4237),
.B(n_4246),
.C(n_4232),
.Y(n_4258)
);

NOR4xp25_ASAP7_75t_L g4259 ( 
.A(n_4234),
.B(n_346),
.C(n_347),
.D(n_348),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4238),
.A2(n_346),
.B(n_348),
.Y(n_4260)
);

OAI21xp5_ASAP7_75t_SL g4261 ( 
.A1(n_4240),
.A2(n_349),
.B(n_350),
.Y(n_4261)
);

NOR2x1_ASAP7_75t_L g4262 ( 
.A(n_4239),
.B(n_349),
.Y(n_4262)
);

INVx1_ASAP7_75t_SL g4263 ( 
.A(n_4249),
.Y(n_4263)
);

NOR2xp33_ASAP7_75t_L g4264 ( 
.A(n_4248),
.B(n_4243),
.Y(n_4264)
);

AOI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_4253),
.A2(n_3008),
.B1(n_3051),
.B2(n_3073),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4260),
.B(n_350),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4251),
.A2(n_3074),
.B1(n_3073),
.B2(n_3062),
.Y(n_4267)
);

AOI211xp5_ASAP7_75t_L g4268 ( 
.A1(n_4247),
.A2(n_351),
.B(n_352),
.C(n_353),
.Y(n_4268)
);

OAI211xp5_ASAP7_75t_L g4269 ( 
.A1(n_4252),
.A2(n_4261),
.B(n_4255),
.C(n_4257),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4254),
.A2(n_351),
.B(n_352),
.Y(n_4270)
);

OAI221xp5_ASAP7_75t_L g4271 ( 
.A1(n_4259),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.C(n_357),
.Y(n_4271)
);

O2A1O1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_4256),
.A2(n_355),
.B(n_356),
.C(n_357),
.Y(n_4272)
);

AND4x2_ASAP7_75t_L g4273 ( 
.A(n_4270),
.B(n_4262),
.C(n_4250),
.D(n_4258),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4266),
.B(n_358),
.Y(n_4274)
);

NAND2xp33_ASAP7_75t_L g4275 ( 
.A(n_4263),
.B(n_359),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4268),
.B(n_4272),
.Y(n_4276)
);

NAND3xp33_ASAP7_75t_L g4277 ( 
.A(n_4264),
.B(n_359),
.C(n_361),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4271),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_4278),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4275),
.B(n_4269),
.Y(n_4280)
);

INVxp33_ASAP7_75t_SL g4281 ( 
.A(n_4276),
.Y(n_4281)
);

NAND4xp25_ASAP7_75t_L g4282 ( 
.A(n_4277),
.B(n_4267),
.C(n_4265),
.D(n_363),
.Y(n_4282)
);

INVxp67_ASAP7_75t_SL g4283 ( 
.A(n_4274),
.Y(n_4283)
);

AOI21xp5_ASAP7_75t_SL g4284 ( 
.A1(n_4280),
.A2(n_4273),
.B(n_362),
.Y(n_4284)
);

AOI21xp33_ASAP7_75t_L g4285 ( 
.A1(n_4279),
.A2(n_361),
.B(n_362),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4285),
.B(n_4283),
.Y(n_4286)
);

NAND3xp33_ASAP7_75t_L g4287 ( 
.A(n_4284),
.B(n_4282),
.C(n_4281),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4286),
.Y(n_4288)
);

OAI22x1_ASAP7_75t_SL g4289 ( 
.A1(n_4288),
.A2(n_4287),
.B1(n_364),
.B2(n_365),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4289),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4290),
.Y(n_4291)
);

HB1xp67_ASAP7_75t_L g4292 ( 
.A(n_4291),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4292),
.Y(n_4293)
);

AOI22xp33_ASAP7_75t_L g4294 ( 
.A1(n_4293),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_4294)
);

NOR2x1_ASAP7_75t_L g4295 ( 
.A(n_4294),
.B(n_367),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_4294),
.A2(n_367),
.B(n_368),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4296),
.B(n_368),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_SL g4298 ( 
.A1(n_4295),
.A2(n_369),
.B(n_370),
.Y(n_4298)
);

AOI322xp5_ASAP7_75t_L g4299 ( 
.A1(n_4297),
.A2(n_370),
.A3(n_371),
.B1(n_372),
.B2(n_373),
.C1(n_374),
.C2(n_375),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4298),
.A2(n_371),
.B(n_374),
.Y(n_4300)
);

OR2x6_ASAP7_75t_L g4301 ( 
.A(n_4300),
.B(n_375),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4301),
.A2(n_4299),
.B(n_377),
.Y(n_4302)
);

AOI211xp5_ASAP7_75t_L g4303 ( 
.A1(n_4302),
.A2(n_376),
.B(n_379),
.C(n_380),
.Y(n_4303)
);


endmodule