module fake_jpeg_10709_n_469 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_63),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_18),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_44),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_19),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_62),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_17),
.B(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_0),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_20),
.B1(n_42),
.B2(n_24),
.Y(n_98)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g86 ( 
.A(n_26),
.B(n_1),
.CON(n_86),
.SN(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_26),
.B1(n_41),
.B2(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_89),
.A2(n_93),
.B1(n_128),
.B2(n_136),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_26),
.B1(n_30),
.B2(n_21),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_30),
.B1(n_21),
.B2(n_36),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_97),
.B1(n_69),
.B2(n_102),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_98),
.A2(n_107),
.B1(n_54),
.B2(n_46),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_42),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_103),
.B(n_104),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_134),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_107)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_88),
.B1(n_81),
.B2(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_49),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_34),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_29),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_44),
.B1(n_29),
.B2(n_23),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_80),
.B(n_15),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_44),
.B1(n_23),
.B2(n_22),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_50),
.B(n_22),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_137),
.B(n_145),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_5),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_35),
.B(n_6),
.C(n_7),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_52),
.B(n_15),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_55),
.B(n_5),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_65),
.Y(n_166)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_130),
.B1(n_97),
.B2(n_119),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_149),
.A2(n_124),
.B(n_108),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_153),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_75),
.B1(n_87),
.B2(n_83),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_151),
.A2(n_160),
.B1(n_195),
.B2(n_118),
.Y(n_234)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_158),
.B(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_166),
.B(n_168),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_112),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_169),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_99),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_84),
.B1(n_66),
.B2(n_64),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_173),
.A2(n_175),
.B1(n_202),
.B2(n_124),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_53),
.B1(n_35),
.B2(n_7),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_188),
.B1(n_140),
.B2(n_139),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_109),
.A2(n_35),
.B(n_6),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_177),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_123),
.B(n_131),
.C(n_129),
.Y(n_206)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_5),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_196),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_106),
.B(n_6),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_106),
.B(n_8),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_140),
.C(n_101),
.Y(n_216)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_121),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_194),
.B1(n_125),
.B2(n_116),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_94),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_94),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_138),
.A2(n_11),
.B1(n_14),
.B2(n_144),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_205),
.A2(n_220),
.B1(n_224),
.B2(n_232),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_217),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g208 ( 
.A(n_152),
.B(n_131),
.C(n_141),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_237),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_149),
.A2(n_174),
.B(n_153),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_209),
.A2(n_250),
.B(n_194),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_100),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_213),
.B(n_221),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_216),
.B(n_182),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_175),
.A2(n_100),
.B1(n_139),
.B2(n_109),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_131),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_180),
.B1(n_200),
.B2(n_165),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_230),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_226),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_118),
.C(n_132),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_163),
.B1(n_190),
.B2(n_183),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_155),
.B(n_116),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_159),
.B(n_181),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_171),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_125),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_182),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_257),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_178),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_197),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_R g261 ( 
.A(n_216),
.B(n_179),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_261),
.A2(n_293),
.B(n_163),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_263),
.B(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_148),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_265),
.B(n_273),
.Y(n_313)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_278),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_277),
.Y(n_319)
);

BUFx12_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g273 ( 
.A1(n_209),
.A2(n_162),
.B1(n_201),
.B2(n_191),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_217),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_193),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_279),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_185),
.B1(n_147),
.B2(n_157),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_280),
.B(n_284),
.Y(n_330)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_249),
.A2(n_161),
.B1(n_169),
.B2(n_172),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_188),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_210),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_221),
.B(n_198),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_234),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_234),
.B1(n_237),
.B2(n_223),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_294),
.B1(n_229),
.B2(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_206),
.B(n_243),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_234),
.A2(n_156),
.B1(n_196),
.B2(n_132),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_236),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_266),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_311),
.C(n_314),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_265),
.B(n_260),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_323),
.B1(n_324),
.B2(n_294),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_258),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_331),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_205),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_220),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_223),
.B(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_315),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_321),
.B(n_293),
.C(n_328),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_283),
.A2(n_226),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_322),
.B(n_326),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_219),
.B1(n_211),
.B2(n_239),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_283),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_254),
.C(n_252),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_297),
.C(n_299),
.Y(n_356)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_271),
.Y(n_331)
);

AND2x6_ASAP7_75t_SL g391 ( 
.A(n_334),
.B(n_271),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_357),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_289),
.B1(n_259),
.B2(n_282),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_323),
.A2(n_291),
.B1(n_280),
.B2(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_273),
.B1(n_277),
.B2(n_270),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g385 ( 
.A1(n_341),
.A2(n_262),
.B(n_312),
.C(n_316),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_296),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_342),
.B(n_350),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_257),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_346),
.C(n_356),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_267),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_256),
.Y(n_347)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_348),
.B(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_275),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_353),
.B(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_305),
.B(n_274),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_354),
.B(n_364),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_272),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_316),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_313),
.A2(n_273),
.B1(n_219),
.B2(n_211),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_358),
.A2(n_330),
.B1(n_307),
.B2(n_308),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_326),
.C(n_299),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_292),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_363),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_313),
.B(n_276),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_362),
.B(n_365),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_255),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_242),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_331),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_369),
.B(n_348),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_362),
.A2(n_322),
.B1(n_330),
.B2(n_306),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_372),
.B1(n_374),
.B2(n_368),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_319),
.B(n_315),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

AO22x1_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_306),
.B1(n_321),
.B2(n_325),
.Y(n_373)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_335),
.A2(n_324),
.B1(n_303),
.B2(n_307),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_380),
.C(n_388),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_310),
.Y(n_380)
);

NOR4xp25_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_333),
.C(n_262),
.D(n_310),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_334),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_337),
.A2(n_312),
.B1(n_332),
.B2(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_345),
.B(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_391),
.A2(n_339),
.B1(n_358),
.B2(n_341),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_338),
.B1(n_349),
.B2(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_393),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_381),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_367),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_406),
.Y(n_413)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_356),
.C(n_346),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_403),
.C(n_405),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_399),
.A2(n_400),
.B1(n_391),
.B2(n_371),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_359),
.C(n_363),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_343),
.C(n_361),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_339),
.C(n_355),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_357),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_381),
.Y(n_427)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_378),
.A2(n_357),
.B1(n_318),
.B2(n_239),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_410),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_384),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_366),
.A2(n_318),
.B1(n_240),
.B2(n_233),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_383),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_374),
.B1(n_370),
.B2(n_379),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_414),
.A2(n_424),
.B1(n_430),
.B2(n_399),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_427),
.C(n_428),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_419),
.A2(n_385),
.B1(n_405),
.B2(n_395),
.Y(n_433)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_402),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_422),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_412),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_425),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_404),
.A2(n_383),
.B1(n_390),
.B2(n_366),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_390),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_426),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_373),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_375),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_429),
.B(n_394),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_392),
.A2(n_385),
.B1(n_373),
.B2(n_369),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_433),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_400),
.B1(n_404),
.B2(n_385),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_434),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_398),
.C(n_403),
.Y(n_434)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_424),
.A2(n_229),
.B(n_233),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_246),
.C(n_199),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_442),
.C(n_415),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_441),
.B(n_443),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_SL g442 ( 
.A1(n_430),
.A2(n_419),
.B(n_414),
.C(n_428),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_417),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_440),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_413),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_447),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_416),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_427),
.C(n_440),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_435),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_446),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_454),
.B(n_455),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_433),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_457),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_452),
.A2(n_442),
.B1(n_438),
.B2(n_439),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_448),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_453),
.A2(n_449),
.B(n_444),
.Y(n_459)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_459),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_456),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_448),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_463),
.B(n_462),
.C(n_460),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_466),
.B(n_450),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_455),
.C(n_442),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_458),
.Y(n_469)
);


endmodule