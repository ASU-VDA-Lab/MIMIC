module real_jpeg_27630_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_296, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_296;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_29),
.B1(n_35),
.B2(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_73),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_131),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_131),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_131),
.Y(n_217)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_4),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_143),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_143),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_143),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_6),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_87),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_87),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_90)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_64),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_10),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_46),
.B(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_10),
.B(n_48),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_62),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_62),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_10),
.B(n_102),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_10),
.A2(n_27),
.B1(n_33),
.B2(n_223),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_10),
.A2(n_49),
.B(n_238),
.Y(n_237)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_12),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_12),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_41),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_13),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_105),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_105),
.Y(n_242)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_84)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_17),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_17),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_17),
.A2(n_29),
.B1(n_35),
.B2(n_54),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_121),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_106),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_22),
.B(n_106),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_92),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_23),
.B(n_76),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_56),
.B1(n_57),
.B2(n_75),
.Y(n_23)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_38),
.B(n_56),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_277)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_27),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_33),
.B1(n_96),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_27),
.A2(n_33),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_27),
.A2(n_33),
.B1(n_217),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_27),
.A2(n_33),
.B1(n_212),
.B2(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_28),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_28),
.A2(n_31),
.B1(n_148),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_28),
.A2(n_31),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_35),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_29),
.B(n_69),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_33),
.B(n_140),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_35),
.A2(n_62),
.A3(n_68),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_53),
.B2(n_55),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_40),
.A2(n_45),
.B1(n_48),
.B2(n_104),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_42),
.A2(n_52),
.B(n_140),
.C(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_44),
.A2(n_55),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_45),
.A2(n_48),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_48),
.B1(n_104),
.B2(n_171),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_79),
.B(n_81),
.C(n_84),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_82),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_49),
.A2(n_63),
.A3(n_82),
.B1(n_239),
.B2(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_50),
.B(n_140),
.Y(n_239)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_98),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_62),
.B(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_65),
.A2(n_74),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_65),
.A2(n_74),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_67),
.B(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_67),
.B1(n_98),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_66),
.A2(n_67),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_66),
.A2(n_67),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_66),
.A2(n_67),
.B1(n_136),
.B2(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_67),
.B(n_140),
.Y(n_224)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_89),
.B(n_91),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_84),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_78),
.A2(n_84),
.B1(n_132),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_78),
.A2(n_84),
.B1(n_155),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_107),
.CI(n_119),
.CON(n_106),
.SN(n_106)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_92),
.A2(n_93),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_103),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_94),
.B(n_99),
.CI(n_103),
.CON(n_276),
.SN(n_276)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_97),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_102),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_102),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_106),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_118),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

AOI321xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_274),
.A3(n_282),
.B1(n_287),
.B2(n_292),
.C(n_296),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_176),
.C(n_188),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_159),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_124),
.B(n_159),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_144),
.C(n_151),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_125),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_138),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_134),
.C(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_144),
.A2(n_151),
.B1(n_152),
.B2(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_144),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_147),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_153),
.B(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_156),
.B(n_158),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_157),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_166),
.C(n_167),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_164),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_172),
.C(n_175),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_177),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_178),
.B(n_179),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_181),
.B(n_182),
.C(n_187),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_268),
.B(n_273),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_254),
.B(n_267),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_232),
.B(n_253),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_213),
.B(n_231),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_208),
.C(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B(n_230),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_219),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_229),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_244),
.C(n_252),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_249),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_263),
.C(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_277),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_276),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_288),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);


endmodule