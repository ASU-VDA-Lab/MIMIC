module fake_aes_5969_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_4), .B(n_11), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_1), .B(n_7), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx5_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_15), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_18), .B1(n_20), .B2(n_15), .Y(n_23) );
OAI211xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B(n_20), .C(n_0), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
NOR2xp67_ASAP7_75t_L g26 ( .A(n_24), .B(n_0), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_20), .B1(n_1), .B2(n_6), .C(n_8), .Y(n_27) );
OA21x2_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_3), .B(n_9), .Y(n_28) );
XOR2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_10), .Y(n_29) );
XNOR2xp5_ASAP7_75t_L g30 ( .A(n_29), .B(n_27), .Y(n_30) );
endmodule