module fake_jpeg_1605_n_669 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_669);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_669;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_60),
.B(n_94),
.Y(n_136)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_63),
.Y(n_182)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g219 ( 
.A(n_65),
.Y(n_219)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_72),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_74),
.B(n_119),
.Y(n_174)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_88),
.Y(n_210)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_124),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_104),
.B(n_48),
.Y(n_176)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_0),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_4),
.Y(n_198)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_41),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_113),
.A2(n_55),
.B1(n_43),
.B2(n_35),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

CKINVDCx6p67_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_32),
.B(n_1),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_32),
.B(n_59),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_121),
.B(n_127),
.Y(n_185)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_46),
.Y(n_122)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_122),
.Y(n_133)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_26),
.B(n_1),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_35),
.B(n_3),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_27),
.Y(n_130)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_67),
.A2(n_57),
.B1(n_28),
.B2(n_34),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_138),
.A2(n_146),
.B1(n_154),
.B2(n_155),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_143),
.B(n_148),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_74),
.A2(n_33),
.B1(n_48),
.B2(n_43),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_27),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_28),
.B1(n_34),
.B2(n_52),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_62),
.B1(n_100),
.B2(n_102),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_47),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_162),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_71),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_47),
.B1(n_39),
.B2(n_52),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_164),
.A2(n_18),
.B1(n_221),
.B2(n_200),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_166),
.A2(n_196),
.B1(n_17),
.B2(n_18),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_106),
.A2(n_55),
.B1(n_50),
.B2(n_39),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_167),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_96),
.B(n_57),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_170),
.B(n_198),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_75),
.A2(n_50),
.B(n_46),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_179),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_77),
.A2(n_46),
.B(n_4),
.C(n_5),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_175),
.A2(n_158),
.B(n_206),
.C(n_170),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_176),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_89),
.B(n_48),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_181),
.B(n_197),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_3),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_183),
.B(n_187),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_3),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_131),
.A2(n_129),
.B1(n_70),
.B2(n_79),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_108),
.B(n_4),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_63),
.B(n_46),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_200),
.B(n_205),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_128),
.B(n_6),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_109),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_206),
.A2(n_221),
.B1(n_188),
.B2(n_180),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_84),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_211),
.B(n_136),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_85),
.B(n_8),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_214),
.B(n_133),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_88),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_125),
.B1(n_116),
.B2(n_14),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_229),
.A2(n_251),
.B(n_288),
.Y(n_351)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_230),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_219),
.Y(n_231)
);

INVx4_ASAP7_75t_SL g340 ( 
.A(n_231),
.Y(n_340)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

BUFx2_ASAP7_75t_SL g329 ( 
.A(n_235),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_150),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_236),
.B(n_244),
.Y(n_321)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_178),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_238),
.A2(n_259),
.B1(n_279),
.B2(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_240),
.Y(n_363)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_241)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_150),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_246),
.Y(n_338)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_247),
.Y(n_361)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_248),
.Y(n_349)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_249),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_250),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_190),
.A2(n_212),
.B1(n_204),
.B2(n_220),
.Y(n_251)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_145),
.Y(n_254)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_139),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_255),
.B(n_258),
.Y(n_339)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

BUFx8_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_139),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_262),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_147),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_269),
.Y(n_313)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_135),
.Y(n_264)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_177),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_173),
.Y(n_270)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

NOR2x1_ASAP7_75t_R g272 ( 
.A(n_175),
.B(n_17),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_L g368 ( 
.A1(n_272),
.A2(n_277),
.B(n_286),
.Y(n_368)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_274),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_210),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_224),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_281),
.Y(n_315)
);

NOR2x1_ASAP7_75t_R g277 ( 
.A(n_141),
.B(n_17),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_278),
.A2(n_259),
.B1(n_287),
.B2(n_302),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_201),
.A2(n_18),
.B1(n_203),
.B2(n_213),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_280),
.A2(n_295),
.B(n_305),
.Y(n_336)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_159),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_282),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_137),
.A2(n_156),
.B1(n_174),
.B2(n_159),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_151),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_134),
.A2(n_199),
.B1(n_218),
.B2(n_171),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_151),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_299),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_149),
.A2(n_152),
.B1(n_210),
.B2(n_144),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_284),
.B1(n_294),
.B2(n_292),
.Y(n_347)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_185),
.A2(n_169),
.A3(n_171),
.B1(n_186),
.B2(n_140),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g342 ( 
.A1(n_291),
.A2(n_271),
.A3(n_286),
.B1(n_261),
.B2(n_230),
.Y(n_342)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_156),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_300),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_142),
.B(n_189),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_294),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_160),
.B(n_207),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_193),
.A2(n_222),
.B1(n_169),
.B2(n_209),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_303),
.B1(n_304),
.B2(n_309),
.Y(n_314)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_135),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_298),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_163),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_202),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_301),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_193),
.A2(n_209),
.B1(n_186),
.B2(n_191),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_202),
.Y(n_304)
);

A2O1A1O1Ixp25_ASAP7_75t_L g305 ( 
.A1(n_133),
.A2(n_138),
.B(n_188),
.C(n_224),
.D(n_157),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_153),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_308),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_168),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_180),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_188),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_310),
.A2(n_311),
.B1(n_257),
.B2(n_231),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_265),
.A2(n_224),
.B(n_157),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_325),
.A2(n_355),
.B(n_363),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_287),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_353),
.C(n_366),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_232),
.A2(n_252),
.B1(n_305),
.B2(n_296),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_337),
.A2(n_267),
.B1(n_282),
.B2(n_270),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_343),
.A2(n_329),
.B1(n_319),
.B2(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_293),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_367),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_272),
.A2(n_278),
.B1(n_277),
.B2(n_287),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_350),
.A2(n_354),
.B1(n_355),
.B2(n_333),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_241),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_300),
.A2(n_281),
.B1(n_266),
.B2(n_250),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_240),
.A2(n_241),
.B(n_249),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_SL g359 ( 
.A1(n_257),
.A2(n_243),
.B(n_239),
.C(n_235),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_237),
.B(n_247),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_233),
.B(n_248),
.C(n_245),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_256),
.B(n_262),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_242),
.A2(n_268),
.B(n_276),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_253),
.B(n_264),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_324),
.B(n_274),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_374),
.B(n_381),
.Y(n_442)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_377),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_378),
.A2(n_394),
.B1(n_420),
.B2(n_357),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_379),
.A2(n_387),
.B(n_392),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_324),
.B(n_346),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_234),
.B1(n_304),
.B2(n_301),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_382),
.A2(n_389),
.B1(n_399),
.B2(n_405),
.Y(n_455)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_313),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_406),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_285),
.B(n_289),
.Y(n_387)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_326),
.A2(n_310),
.B1(n_246),
.B2(n_298),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_326),
.B(n_325),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_393),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_327),
.A2(n_314),
.B1(n_353),
.B2(n_331),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_321),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_400),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_371),
.B(n_339),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_396),
.A2(n_398),
.B(n_407),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_363),
.B(n_315),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_354),
.B1(n_334),
.B2(n_369),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_366),
.B(n_352),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_402),
.A2(n_403),
.B(n_412),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_323),
.A2(n_316),
.B(n_312),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_341),
.C(n_358),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_400),
.C(n_386),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_332),
.A2(n_358),
.B1(n_364),
.B2(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_315),
.A2(n_370),
.B(n_312),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_318),
.B(n_345),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_409),
.Y(n_447)
);

AO22x1_ASAP7_75t_SL g409 ( 
.A1(n_322),
.A2(n_315),
.B1(n_349),
.B2(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_413),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_372),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_370),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_391),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_320),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_417),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_340),
.A2(n_356),
.B(n_330),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_416),
.A2(n_396),
.B(n_377),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_330),
.B(n_320),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_365),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_409),
.Y(n_454)
);

INVx11_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_419),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_338),
.A2(n_364),
.B1(n_348),
.B2(n_319),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_421),
.A2(n_372),
.B1(n_349),
.B2(n_365),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_422),
.A2(n_441),
.B1(n_452),
.B2(n_403),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_415),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_436),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_SL g470 ( 
.A1(n_426),
.A2(n_398),
.B(n_416),
.Y(n_470)
);

AOI21x1_ASAP7_75t_SL g476 ( 
.A1(n_427),
.A2(n_407),
.B(n_383),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_378),
.A2(n_394),
.B1(n_401),
.B2(n_384),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_434),
.A2(n_437),
.B1(n_459),
.B2(n_424),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_404),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_401),
.A2(n_399),
.B1(n_382),
.B2(n_390),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_418),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_443),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_401),
.A2(n_381),
.B1(n_390),
.B2(n_411),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_450),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_374),
.B(n_380),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_454),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_380),
.B(n_402),
.Y(n_450)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_451),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_421),
.A2(n_373),
.B1(n_392),
.B2(n_389),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_395),
.B(n_414),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_387),
.B1(n_385),
.B2(n_379),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_376),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_409),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_460),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_462),
.B(n_463),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_433),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_465),
.A2(n_475),
.B1(n_486),
.B2(n_494),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_443),
.B(n_393),
.Y(n_466)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_425),
.Y(n_535)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_471),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_433),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_473),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_453),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_434),
.A2(n_426),
.B1(n_441),
.B2(n_454),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_476),
.A2(n_496),
.B(n_449),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_453),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_477),
.B(n_480),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_444),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_442),
.B(n_435),
.Y(n_481)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_431),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_484),
.B(n_491),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_458),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_485),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_437),
.A2(n_412),
.B1(n_420),
.B2(n_417),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_412),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_450),
.C(n_436),
.Y(n_501)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_447),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_489),
.Y(n_508)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_490),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_451),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_493),
.A2(n_424),
.B1(n_452),
.B2(n_449),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_447),
.A2(n_405),
.B1(n_409),
.B2(n_397),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_423),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_495),
.B(n_422),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_459),
.A2(n_444),
.B(n_427),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_438),
.B(n_410),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_498),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_432),
.B(n_406),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_499),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_501),
.B(n_512),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_506),
.B1(n_493),
.B2(n_535),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_445),
.C(n_446),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_525),
.C(n_533),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_465),
.A2(n_439),
.B1(n_427),
.B2(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_469),
.B(n_429),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_520),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_479),
.B(n_429),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_442),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_527),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_499),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_521),
.A2(n_523),
.B(n_534),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_476),
.A2(n_461),
.B(n_455),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_456),
.C(n_435),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_474),
.B(n_461),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_474),
.B(n_456),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_518),
.Y(n_550)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_464),
.B(n_491),
.C(n_496),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_485),
.A2(n_455),
.B1(n_440),
.B2(n_425),
.Y(n_534)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_486),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_495),
.Y(n_536)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_516),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_537),
.B(n_543),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_538),
.A2(n_554),
.B1(n_558),
.B2(n_566),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_489),
.Y(n_541)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_464),
.C(n_490),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_548),
.C(n_559),
.Y(n_569)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_524),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_547),
.B(n_550),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_501),
.B(n_498),
.C(n_462),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_512),
.B(n_525),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_563),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_478),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_555),
.Y(n_590)
);

NOR2x1_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_556),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_514),
.A2(n_519),
.B1(n_475),
.B2(n_517),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_472),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_473),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_560),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_519),
.A2(n_494),
.B1(n_477),
.B2(n_484),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_463),
.C(n_497),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_500),
.B(n_497),
.C(n_481),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_507),
.C(n_511),
.Y(n_570)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_562),
.B(n_564),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_466),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_508),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_565),
.B(n_529),
.Y(n_583)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_505),
.Y(n_566)
);

FAx1_ASAP7_75t_SL g567 ( 
.A(n_559),
.B(n_531),
.CI(n_521),
.CON(n_567),
.SN(n_567)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_567),
.B(n_570),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_502),
.C(n_523),
.Y(n_571)
);

MAJx2_ASAP7_75t_L g603 ( 
.A(n_571),
.B(n_576),
.C(n_577),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_535),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_544),
.B(n_534),
.C(n_506),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_440),
.C(n_503),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_586),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_546),
.B(n_482),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g607 ( 
.A(n_580),
.B(n_553),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_529),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_585),
.Y(n_604)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_583),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_546),
.B(n_528),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_539),
.B(n_503),
.C(n_513),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_540),
.B(n_467),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_492),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_539),
.B(n_528),
.C(n_513),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_488),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_536),
.Y(n_591)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_591),
.Y(n_597)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_592),
.Y(n_613)
);

CKINVDCx14_ASAP7_75t_R g594 ( 
.A(n_590),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_594),
.B(n_598),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_568),
.A2(n_547),
.B1(n_554),
.B2(n_542),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_595),
.A2(n_599),
.B1(n_601),
.B2(n_584),
.Y(n_624)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_572),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_610),
.Y(n_621)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_570),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_574),
.A2(n_558),
.B1(n_538),
.B2(n_556),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_582),
.A2(n_541),
.B1(n_549),
.B2(n_540),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_573),
.A2(n_561),
.B1(n_566),
.B2(n_563),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_602),
.B(n_606),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_577),
.A2(n_505),
.B1(n_550),
.B2(n_471),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_580),
.Y(n_620)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_589),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_609),
.B(n_611),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_576),
.B(n_483),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_601),
.A2(n_575),
.B(n_571),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_612),
.A2(n_614),
.B(n_617),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_600),
.A2(n_588),
.B(n_567),
.Y(n_614)
);

INVx11_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_615),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_605),
.B(n_569),
.C(n_579),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_SL g640 ( 
.A(n_616),
.B(n_457),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_587),
.B(n_581),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_609),
.A2(n_585),
.B(n_569),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_618),
.A2(n_627),
.B(n_607),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_620),
.B(n_628),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_622),
.A2(n_596),
.B1(n_597),
.B2(n_604),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_586),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_623),
.B(n_624),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_SL g627 ( 
.A(n_605),
.B(n_584),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_603),
.B(n_468),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_616),
.B(n_610),
.C(n_604),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_630),
.B(n_634),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_592),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_632),
.B(n_621),
.Y(n_647)
);

AO21x1_ASAP7_75t_L g646 ( 
.A1(n_633),
.A2(n_614),
.B(n_617),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_625),
.B(n_595),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_611),
.C(n_599),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_635),
.B(n_636),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_619),
.B(n_457),
.Y(n_636)
);

MAJx2_ASAP7_75t_L g648 ( 
.A(n_639),
.B(n_628),
.C(n_624),
.Y(n_648)
);

AOI21x1_ASAP7_75t_SL g650 ( 
.A1(n_640),
.A2(n_615),
.B(n_626),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_618),
.B(n_448),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_641),
.B(n_388),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_448),
.C(n_397),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_642),
.B(n_621),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_645),
.B(n_646),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_647),
.B(n_652),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_648),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_630),
.B(n_626),
.C(n_620),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_649),
.B(n_635),
.C(n_629),
.Y(n_653)
);

AOI21xp33_ASAP7_75t_L g654 ( 
.A1(n_650),
.A2(n_651),
.B(n_631),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_637),
.B(n_629),
.Y(n_651)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_653),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_654),
.A2(n_658),
.B(n_659),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_642),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_641),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_657),
.A2(n_643),
.B(n_644),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_661),
.A2(n_663),
.B(n_656),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_656),
.A2(n_638),
.B(n_419),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_664),
.A2(n_665),
.B1(n_655),
.B2(n_662),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_660),
.Y(n_665)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_666),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_667),
.B(n_638),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_668),
.B(n_419),
.C(n_388),
.Y(n_669)
);


endmodule