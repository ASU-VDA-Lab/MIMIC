module fake_jpeg_1267_n_614 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_614);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_614;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_58),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_59),
.B(n_60),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_22),
.B(n_9),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_61),
.Y(n_181)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_9),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_69),
.Y(n_209)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_73),
.B(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_78),
.B(n_86),
.Y(n_169)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_10),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_93),
.Y(n_220)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_102),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_39),
.A2(n_10),
.B(n_18),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_101),
.B(n_0),
.C(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_103),
.B(n_123),
.Y(n_177)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_104),
.Y(n_221)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_114),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_115),
.B(n_116),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_28),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_118),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_0),
.Y(n_204)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_48),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_51),
.B(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_124),
.B(n_11),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_31),
.Y(n_126)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_43),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_33),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_24),
.Y(n_128)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_77),
.B(n_35),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_131),
.B(n_138),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_46),
.B1(n_44),
.B2(n_31),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_135),
.A2(n_139),
.B1(n_141),
.B2(n_149),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_55),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_72),
.B(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_43),
.B1(n_33),
.B2(n_24),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_46),
.B1(n_24),
.B2(n_57),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_69),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_145),
.B(n_194),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_57),
.B1(n_53),
.B2(n_39),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_72),
.A2(n_57),
.B1(n_55),
.B2(n_35),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_156),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_80),
.A2(n_104),
.B1(n_107),
.B2(n_114),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_71),
.B(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_153),
.B(n_218),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_129),
.B1(n_63),
.B2(n_112),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_90),
.A2(n_33),
.B1(n_57),
.B2(n_21),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_64),
.A2(n_33),
.B1(n_21),
.B2(n_47),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_157),
.A2(n_158),
.B1(n_178),
.B2(n_185),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_74),
.A2(n_47),
.B1(n_26),
.B2(n_50),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_101),
.A2(n_46),
.B1(n_50),
.B2(n_30),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_166),
.B(n_174),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_58),
.A2(n_26),
.B1(n_50),
.B2(n_29),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_50),
.B1(n_29),
.B2(n_54),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_87),
.A2(n_29),
.B1(n_54),
.B2(n_12),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_75),
.A2(n_54),
.B1(n_11),
.B2(n_12),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_192),
.A2(n_196),
.B1(n_198),
.B2(n_205),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_200),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_76),
.B(n_11),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_84),
.A2(n_113),
.B1(n_105),
.B2(n_108),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_93),
.A2(n_7),
.B1(n_18),
.B2(n_17),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_199),
.A2(n_216),
.B(n_185),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_99),
.B(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_6),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_202),
.B(n_212),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_92),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_83),
.B(n_6),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_61),
.A2(n_5),
.B1(n_13),
.B2(n_12),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_4),
.B1(n_13),
.B2(n_218),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_61),
.B(n_5),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_68),
.B(n_19),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_68),
.B(n_7),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_228),
.Y(n_344)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_166),
.A2(n_81),
.A3(n_117),
.B1(n_106),
.B2(n_13),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_250),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_154),
.A2(n_81),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_233),
.A2(n_240),
.B1(n_271),
.B2(n_283),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_174),
.B(n_1),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_234),
.Y(n_335)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_237),
.Y(n_346)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_239),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_149),
.A2(n_4),
.B1(n_158),
.B2(n_140),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_242),
.A2(n_261),
.B1(n_262),
.B2(n_300),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_259),
.Y(n_314)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_245),
.Y(n_319)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_248),
.Y(n_326)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_249),
.B(n_260),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_251),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_194),
.A2(n_4),
.B1(n_191),
.B2(n_186),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_253),
.A2(n_277),
.B1(n_295),
.B2(n_240),
.Y(n_325)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_133),
.A2(n_4),
.B1(n_179),
.B2(n_151),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_257),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_169),
.B(n_144),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_196),
.A2(n_197),
.B1(n_170),
.B2(n_184),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_164),
.A2(n_188),
.B1(n_211),
.B2(n_134),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_161),
.Y(n_265)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_163),
.B(n_132),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_273),
.Y(n_324)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_136),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_288),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_178),
.A2(n_139),
.B1(n_156),
.B2(n_157),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_168),
.Y(n_272)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_147),
.B(n_137),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_275),
.Y(n_352)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_207),
.A2(n_220),
.B1(n_190),
.B2(n_160),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_294),
.Y(n_328)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_162),
.B(n_136),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_281),
.Y(n_357)
);

BUFx4f_ASAP7_75t_L g282 ( 
.A(n_130),
.Y(n_282)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_217),
.A2(n_182),
.B1(n_203),
.B2(n_207),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_179),
.A2(n_151),
.B1(n_176),
.B2(n_183),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_285),
.A2(n_286),
.B1(n_292),
.B2(n_233),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_183),
.A2(n_221),
.B1(n_130),
.B2(n_173),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_293),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_182),
.A2(n_203),
.B1(n_220),
.B2(n_190),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_292),
.B1(n_307),
.B2(n_246),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_152),
.A2(n_221),
.B1(n_143),
.B2(n_213),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_173),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_146),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_143),
.A2(n_210),
.B1(n_146),
.B2(n_201),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_201),
.B(n_210),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_297),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_159),
.B(n_189),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_181),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_299),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_189),
.A2(n_103),
.B1(n_141),
.B2(n_86),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_219),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_303),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_181),
.B(n_199),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_234),
.Y(n_345)
);

INVx6_ASAP7_75t_SL g303 ( 
.A(n_181),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_155),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_155),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_154),
.A2(n_149),
.B1(n_158),
.B2(n_166),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_311),
.A2(n_325),
.B1(n_341),
.B2(n_348),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_244),
.C(n_268),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_318),
.C(n_321),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_243),
.C(n_273),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_243),
.C(n_252),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_234),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_304),
.B1(n_267),
.B2(n_290),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_230),
.B1(n_293),
.B2(n_272),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_260),
.A2(n_278),
.B1(n_263),
.B2(n_253),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_345),
.B(n_303),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_258),
.A2(n_271),
.B1(n_264),
.B2(n_227),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_247),
.B(n_248),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_354),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_277),
.A2(n_295),
.B1(n_259),
.B2(n_288),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_351),
.A2(n_299),
.B1(n_245),
.B2(n_282),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_231),
.B(n_239),
.Y(n_354)
);

OAI32xp33_ASAP7_75t_L g362 ( 
.A1(n_265),
.A2(n_275),
.A3(n_266),
.B1(n_254),
.B2(n_238),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_364),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_284),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_236),
.B1(n_255),
.B2(n_228),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_366),
.A2(n_367),
.B1(n_377),
.B2(n_378),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_311),
.A2(n_237),
.B1(n_289),
.B2(n_235),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_287),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_376),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_230),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_308),
.A2(n_328),
.B1(n_324),
.B2(n_314),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_328),
.A2(n_320),
.B(n_343),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_379),
.A2(n_397),
.B(n_342),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_324),
.B(n_226),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_381),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_306),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_308),
.A2(n_291),
.B1(n_305),
.B2(n_269),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_382),
.A2(n_388),
.B1(n_399),
.B2(n_402),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_232),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_384),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_314),
.B(n_294),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_328),
.A2(n_283),
.B1(n_282),
.B2(n_257),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_389),
.B(n_350),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_279),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_394),
.Y(n_421)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_274),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_392),
.B(n_393),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_318),
.B(n_345),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_251),
.B1(n_298),
.B2(n_325),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_395),
.A2(n_403),
.B1(n_407),
.B2(n_315),
.Y(n_418)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_400),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_317),
.A2(n_310),
.B(n_334),
.Y(n_397)
);

O2A1O1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_355),
.B(n_360),
.C(n_363),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_410),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_334),
.A2(n_335),
.B1(n_338),
.B2(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_401),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_332),
.A2(n_312),
.B1(n_321),
.B2(n_343),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_362),
.A2(n_329),
.B1(n_337),
.B2(n_352),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_409),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_337),
.A2(n_326),
.B1(n_352),
.B2(n_333),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_406),
.B1(n_365),
.B2(n_410),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_327),
.A2(n_333),
.B1(n_331),
.B2(n_329),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_359),
.A2(n_327),
.B1(n_331),
.B2(n_346),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_309),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_360),
.C(n_363),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_330),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_358),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_375),
.B1(n_396),
.B2(n_400),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_411),
.A2(n_429),
.B1(n_438),
.B2(n_442),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_407),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_412),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_330),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_446),
.C(n_437),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_418),
.A2(n_435),
.B1(n_367),
.B2(n_366),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_406),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_426),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_405),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_309),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_428),
.B(n_408),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_375),
.A2(n_315),
.B1(n_346),
.B2(n_356),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_437),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_356),
.B(n_340),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_432),
.A2(n_434),
.B(n_441),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_385),
.A2(n_344),
.B1(n_342),
.B2(n_340),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_370),
.A2(n_319),
.B1(n_365),
.B2(n_361),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_322),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_440),
.B(n_376),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_379),
.A2(n_339),
.B(n_361),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_385),
.A2(n_344),
.B1(n_322),
.B2(n_350),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_369),
.B(n_353),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_384),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_353),
.C(n_358),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_390),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_448),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_451),
.C(n_459),
.Y(n_503)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_381),
.C(n_389),
.Y(n_451)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

OAI22x1_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_403),
.B1(n_395),
.B2(n_393),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_458),
.A2(n_434),
.B(n_441),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_389),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_421),
.B(n_369),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_460),
.B(n_404),
.Y(n_505)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_416),
.Y(n_463)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_431),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_464),
.B(n_466),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_424),
.A2(n_422),
.B1(n_426),
.B2(n_429),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_465),
.A2(n_479),
.B1(n_482),
.B2(n_418),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_431),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_468),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_421),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_474),
.C(n_475),
.Y(n_510)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

AND2x2_ASAP7_75t_SL g492 ( 
.A(n_470),
.B(n_472),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_424),
.A2(n_392),
.B1(n_378),
.B2(n_380),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_471),
.A2(n_483),
.B1(n_410),
.B2(n_387),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_477),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_402),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_419),
.B(n_399),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_430),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_368),
.C(n_408),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_415),
.A2(n_398),
.B1(n_409),
.B2(n_382),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_481),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_415),
.A2(n_398),
.B1(n_397),
.B2(n_391),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_484),
.A2(n_485),
.B1(n_496),
.B2(n_501),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_465),
.A2(n_436),
.B1(n_435),
.B2(n_412),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_456),
.A2(n_436),
.B1(n_448),
.B2(n_439),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_486),
.A2(n_489),
.B1(n_493),
.B2(n_500),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_504),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_455),
.A2(n_423),
.B1(n_438),
.B2(n_425),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_446),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_497),
.C(n_507),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_456),
.A2(n_439),
.B1(n_423),
.B2(n_420),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_494),
.A2(n_416),
.B(n_463),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_458),
.A2(n_442),
.B1(n_420),
.B2(n_443),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_430),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_461),
.A2(n_397),
.B(n_464),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_499),
.B(n_452),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_455),
.A2(n_414),
.B1(n_432),
.B2(n_417),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_414),
.B1(n_388),
.B2(n_444),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_386),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_505),
.B(n_467),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_401),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_482),
.A2(n_444),
.B1(n_416),
.B2(n_410),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_509),
.A2(n_450),
.B1(n_454),
.B2(n_462),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_387),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_459),
.C(n_480),
.Y(n_528)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_515),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_493),
.B(n_477),
.CI(n_510),
.CON(n_516),
.SN(n_516)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_503),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_486),
.A2(n_478),
.B1(n_481),
.B2(n_470),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_517),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_500),
.A2(n_466),
.B1(n_457),
.B2(n_471),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g545 ( 
.A1(n_520),
.A2(n_540),
.B(n_518),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_512),
.A2(n_475),
.B(n_468),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_521),
.A2(n_524),
.B(n_525),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_494),
.A2(n_461),
.B(n_479),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_526),
.A2(n_534),
.B1(n_506),
.B2(n_502),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_487),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g542 ( 
.A(n_527),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_528),
.B(n_503),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_452),
.Y(n_530)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_530),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_472),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_533),
.Y(n_552)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_512),
.Y(n_532)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_532),
.Y(n_550)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_484),
.A2(n_515),
.B1(n_485),
.B2(n_496),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_538),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_539),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_492),
.A2(n_504),
.B(n_501),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_537),
.A2(n_489),
.B(n_514),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_476),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_498),
.B(n_372),
.Y(n_539)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_553),
.C(n_555),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g566 ( 
.A1(n_544),
.A2(n_523),
.B(n_516),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_545),
.A2(n_559),
.B(n_495),
.Y(n_572)
);

OAI21x1_ASAP7_75t_SL g569 ( 
.A1(n_548),
.A2(n_552),
.B(n_550),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_519),
.A2(n_509),
.B1(n_492),
.B2(n_511),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_549),
.A2(n_520),
.B1(n_522),
.B2(n_526),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_534),
.A2(n_510),
.B1(n_498),
.B2(n_511),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_551),
.A2(n_560),
.B1(n_544),
.B2(n_553),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_490),
.C(n_497),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_488),
.Y(n_555)
);

NAND4xp25_ASAP7_75t_L g557 ( 
.A(n_524),
.B(n_518),
.C(n_525),
.D(n_533),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_545),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_SL g559 ( 
.A1(n_532),
.A2(n_519),
.B(n_522),
.C(n_530),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_495),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_521),
.C(n_539),
.Y(n_568)
);

HAxp5_ASAP7_75t_SL g561 ( 
.A(n_556),
.B(n_528),
.CON(n_561),
.SN(n_561)
);

AOI31xp33_ASAP7_75t_L g582 ( 
.A1(n_561),
.A2(n_566),
.A3(n_574),
.B(n_575),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_542),
.B(n_535),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_562),
.B(n_564),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_563),
.A2(n_571),
.B1(n_559),
.B2(n_558),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_550),
.B(n_531),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_546),
.A2(n_540),
.B(n_537),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_565),
.A2(n_570),
.B1(n_573),
.B2(n_541),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_577),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_577),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_546),
.A2(n_527),
.B(n_536),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_549),
.A2(n_554),
.B1(n_548),
.B2(n_552),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_557),
.A2(n_545),
.B(n_547),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_547),
.A2(n_516),
.B(n_372),
.Y(n_575)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_551),
.C(n_543),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_580),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_555),
.C(n_544),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_583),
.B(n_587),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_562),
.B(n_558),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_584),
.B(n_585),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_559),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_559),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g590 ( 
.A(n_588),
.B(n_572),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_569),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_589),
.B(n_574),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_590),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_587),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_593),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_573),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_576),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_598),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_597),
.B(n_586),
.Y(n_599)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_599),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_586),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_602),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_596),
.B(n_579),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_604),
.A2(n_591),
.B(n_580),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_SL g605 ( 
.A(n_601),
.B(n_600),
.C(n_603),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_605),
.B(n_608),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_581),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_591),
.C(n_601),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_610),
.C(n_609),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_570),
.Y(n_613)
);

FAx1_ASAP7_75t_SL g614 ( 
.A(n_613),
.B(n_607),
.CI(n_575),
.CON(n_614),
.SN(n_614)
);


endmodule