module fake_jpeg_23912_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_16),
.Y(n_63)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_20),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_83),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_41),
.B1(n_58),
.B2(n_37),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_55),
.Y(n_90)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_46),
.B(n_52),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_99),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_89),
.B1(n_76),
.B2(n_48),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_41),
.B1(n_25),
.B2(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_41),
.B1(n_46),
.B2(n_54),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_104),
.B1(n_108),
.B2(n_121),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_65),
.B(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_34),
.B1(n_42),
.B2(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_34),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_74),
.B1(n_86),
.B2(n_73),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_64),
.A3(n_45),
.B1(n_20),
.B2(n_35),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_92),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_64),
.B(n_39),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_87),
.Y(n_125)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_80),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_45),
.B1(n_39),
.B2(n_34),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_127),
.B1(n_101),
.B2(n_104),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_134),
.Y(n_171)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_76),
.B1(n_48),
.B2(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_91),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_69),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_144),
.B(n_148),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_140),
.Y(n_159)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_76),
.B1(n_48),
.B2(n_80),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_147),
.B1(n_122),
.B2(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_45),
.C(n_35),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_102),
.C(n_122),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_68),
.B1(n_77),
.B2(n_32),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_173),
.B1(n_135),
.B2(n_124),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_96),
.B(n_119),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_160),
.B(n_162),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_136),
.B1(n_137),
.B2(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_106),
.B1(n_110),
.B2(n_107),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_161),
.B1(n_169),
.B2(n_172),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_107),
.B(n_109),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_109),
.B(n_112),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_133),
.C(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_45),
.B1(n_84),
.B2(n_115),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_113),
.B1(n_115),
.B2(n_105),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_112),
.B1(n_105),
.B2(n_31),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_32),
.B(n_18),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_182),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_134),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_190),
.B(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_198),
.B1(n_200),
.B2(n_158),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_173),
.B1(n_155),
.B2(n_165),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_131),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_188),
.B(n_25),
.Y(n_227)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_189),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_195),
.C(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_146),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_146),
.C(n_93),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_146),
.B1(n_18),
.B2(n_21),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_30),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_30),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_181),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_212),
.C(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_167),
.B1(n_150),
.B2(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_171),
.C(n_161),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_160),
.C(n_152),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_152),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_219),
.C(n_223),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_151),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_157),
.B1(n_18),
.B2(n_21),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_26),
.B(n_33),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_226),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_157),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_93),
.B1(n_79),
.B2(n_24),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_30),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_187),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_228),
.A2(n_241),
.B(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_200),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_225),
.B1(n_215),
.B2(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_181),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_217),
.A2(n_175),
.B(n_182),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_192),
.C(n_186),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_247),
.C(n_24),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_192),
.C(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_30),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_227),
.B(n_210),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_225),
.B(n_219),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_258),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_215),
.B(n_205),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_223),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_30),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_224),
.B1(n_211),
.B2(n_209),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_226),
.B(n_180),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_247),
.A2(n_180),
.B1(n_79),
.B2(n_25),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_243),
.C(n_230),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_32),
.B1(n_23),
.B2(n_27),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_23),
.B1(n_22),
.B2(n_234),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_234),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_233),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_280),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_233),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_255),
.B(n_27),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_262),
.B1(n_251),
.B2(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_28),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_10),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_28),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_256),
.B1(n_269),
.B2(n_257),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_297),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_254),
.CI(n_268),
.CON(n_293),
.SN(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_275),
.Y(n_302)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_261),
.B1(n_260),
.B2(n_11),
.C(n_13),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_0),
.C(n_1),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_285),
.C(n_284),
.Y(n_305)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_9),
.B(n_15),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_299),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_28),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_306),
.B(n_307),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_310),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_9),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_11),
.C2(n_6),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_33),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_28),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_291),
.B1(n_287),
.B2(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_8),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_293),
.B(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_320),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_289),
.B1(n_298),
.B2(n_33),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_318),
.B1(n_311),
.B2(n_309),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_289),
.B1(n_33),
.B2(n_26),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_26),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_0),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_8),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_1),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_325),
.A2(n_329),
.B(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_7),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_9),
.B(n_11),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_326),
.B(n_325),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_330),
.B(n_331),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_317),
.B1(n_12),
.B2(n_5),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_2),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_3),
.C(n_5),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_3),
.C(n_5),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.Y(n_340)
);


endmodule