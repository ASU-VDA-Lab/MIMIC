module fake_jpeg_14627_n_387 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_11),
.CON(n_44),
.SN(n_44)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_0),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_51),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_61),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_74),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_14),
.B1(n_26),
.B2(n_32),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_70),
.A2(n_77),
.B1(n_37),
.B2(n_63),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_14),
.B1(n_26),
.B2(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_14),
.B1(n_26),
.B2(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_78),
.A2(n_92),
.B1(n_96),
.B2(n_110),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_90),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_95),
.B1(n_22),
.B2(n_23),
.Y(n_127)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_109),
.Y(n_124)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_42),
.A2(n_37),
.B1(n_19),
.B2(n_36),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_38),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_102),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_104),
.B(n_1),
.CON(n_154),
.SN(n_154)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_31),
.Y(n_112)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_1),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_53),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_55),
.B1(n_49),
.B2(n_46),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_28),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_118),
.A2(n_162),
.B1(n_133),
.B2(n_123),
.Y(n_208)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_125),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_167),
.B1(n_161),
.B2(n_129),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_127),
.A2(n_118),
.B(n_163),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_131),
.Y(n_185)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_53),
.B1(n_55),
.B2(n_63),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_138),
.B1(n_144),
.B2(n_152),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_60),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_165),
.C(n_99),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_37),
.B1(n_33),
.B2(n_34),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_71),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_139),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_82),
.B(n_1),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_33),
.B(n_34),
.C(n_60),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_154),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_109),
.B(n_33),
.Y(n_148)
);

NOR2x1_ASAP7_75t_R g194 ( 
.A(n_148),
.B(n_76),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_34),
.Y(n_149)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_153),
.Y(n_186)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_71),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_90),
.B1(n_93),
.B2(n_99),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_2),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_164),
.Y(n_198)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_163),
.B1(n_107),
.B2(n_101),
.Y(n_176)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_2),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_6),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_6),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_72),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_201),
.B(n_205),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_208),
.Y(n_227)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_176),
.A2(n_181),
.B1(n_183),
.B2(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_184),
.Y(n_225)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_80),
.B1(n_100),
.B2(n_94),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_170),
.B1(n_184),
.B2(n_194),
.Y(n_220)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_135),
.A2(n_148),
.B1(n_137),
.B2(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_196),
.B1(n_200),
.B2(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_72),
.B1(n_76),
.B2(n_9),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_199),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g247 ( 
.A1(n_194),
.A2(n_148),
.B(n_191),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_126),
.B(n_89),
.CI(n_8),
.CON(n_195),
.SN(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_202),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_155),
.Y(n_200)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_117),
.A2(n_10),
.A3(n_145),
.B1(n_154),
.B2(n_143),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_132),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_120),
.A2(n_10),
.B1(n_142),
.B2(n_156),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_124),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_151),
.C(n_158),
.Y(n_219)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_141),
.B(n_133),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_214),
.A2(n_229),
.B(n_232),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_134),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_236),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_160),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_216),
.B(n_235),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_220),
.A2(n_228),
.B1(n_230),
.B2(n_233),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_174),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_226),
.C(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_208),
.C(n_205),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_200),
.B1(n_169),
.B2(n_176),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_191),
.B(n_189),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_192),
.B1(n_195),
.B2(n_213),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_198),
.B(n_187),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_190),
.B(n_178),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_230),
.B(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_172),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_171),
.B1(n_173),
.B2(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_236),
.B1(n_244),
.B2(n_220),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_241),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_193),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_242),
.B(n_244),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_179),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_225),
.B1(n_239),
.B2(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_168),
.Y(n_248)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_182),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_207),
.B(n_126),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_198),
.B(n_126),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_252),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_182),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_168),
.B(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_278),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_257),
.B(n_259),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_229),
.B1(n_248),
.B2(n_226),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_276),
.B1(n_271),
.B2(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_268),
.C(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_245),
.B1(n_249),
.B2(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_280),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_237),
.C(n_227),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_234),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_231),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_237),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_287),
.C(n_223),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_286),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g286 ( 
.A(n_249),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_218),
.C(n_221),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_218),
.B(n_232),
.CI(n_214),
.CON(n_288),
.SN(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_299),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_262),
.A2(n_222),
.B1(n_253),
.B2(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_217),
.C(n_223),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_310),
.C(n_286),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_262),
.A2(n_249),
.B1(n_282),
.B2(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_302),
.B(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_300),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_311),
.B1(n_297),
.B2(n_314),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_283),
.C(n_275),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_270),
.A2(n_288),
.B1(n_274),
.B2(n_256),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_279),
.B(n_265),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_277),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_322),
.B(n_327),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_303),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_296),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_330),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_304),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_309),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_316),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_333),
.B(n_290),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_292),
.C(n_306),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_336),
.B(n_337),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_334),
.A2(n_290),
.B(n_312),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_350),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_307),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_342),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_329),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_345),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_335),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_324),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_352),
.B(n_323),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_294),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_318),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_292),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_295),
.C(n_337),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_346),
.A2(n_321),
.B1(n_344),
.B2(n_347),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_358),
.B1(n_331),
.B2(n_338),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_336),
.C(n_339),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_361),
.B(n_339),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_344),
.A2(n_321),
.B1(n_338),
.B2(n_347),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_364),
.C(n_351),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_331),
.B(n_326),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_363),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g364 ( 
.A(n_348),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_326),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_371),
.A2(n_359),
.B1(n_357),
.B2(n_366),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_365),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_372),
.A2(n_335),
.B1(n_328),
.B2(n_325),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_373),
.B(n_374),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_368),
.B1(n_320),
.B2(n_325),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_377),
.B(n_379),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_354),
.C(n_356),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_380),
.B(n_376),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_382),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_381),
.Y(n_384)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_384),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_367),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_386),
.Y(n_387)
);


endmodule