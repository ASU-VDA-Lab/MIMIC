module fake_jpeg_17353_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_24),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_16),
.Y(n_30)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_10),
.B1(n_11),
.B2(n_17),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_23),
.B1(n_24),
.B2(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_21),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_38),
.B1(n_20),
.B2(n_31),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_25),
.B(n_21),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_42),
.B1(n_32),
.B2(n_9),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_12),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_24),
.B1(n_19),
.B2(n_11),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_18),
.B(n_15),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.C(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_22),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_22),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_13),
.Y(n_56)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_40),
.B(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_58),
.B1(n_49),
.B2(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_56),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_47),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_48),
.B1(n_46),
.B2(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_58),
.B1(n_48),
.B2(n_56),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_65),
.B1(n_11),
.B2(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_68),
.A3(n_66),
.B1(n_59),
.B2(n_32),
.C1(n_22),
.C2(n_17),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_61),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_71),
.C(n_59),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_75),
.B(n_13),
.C(n_17),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_7),
.A3(n_8),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_16),
.Y(n_76)
);

AOI31xp67_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_8),
.A3(n_4),
.B(n_3),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_78),
.B(n_0),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_1),
.B(n_22),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_1),
.Y(n_81)
);


endmodule