module fake_netlist_6_3746_n_761 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_761);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_761;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_736;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g153 ( 
.A(n_44),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_111),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_73),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_83),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_26),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_86),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_28),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_97),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_32),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_126),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_43),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_55),
.B(n_70),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_69),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_27),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_37),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_25),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_16),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_75),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_14),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_19),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_54),
.B(n_61),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_42),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_20),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_50),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_53),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_66),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_24),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_106),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_18),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_174),
.B(n_0),
.Y(n_213)
);

AOI22x1_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_1),
.Y(n_218)
);

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_2),
.B(n_3),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_21),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_4),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_179),
.A2(n_5),
.B(n_6),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_5),
.B(n_6),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_158),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_184),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_192),
.B(n_172),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_155),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_181),
.B1(n_169),
.B2(n_163),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_161),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

BUFx6f_ASAP7_75t_SL g269 ( 
.A(n_217),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_185),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

BUFx6f_ASAP7_75t_SL g276 ( 
.A(n_217),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_205),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_246),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_248),
.B(n_165),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_166),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_167),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_212),
.B(n_168),
.Y(n_290)
);

CKINVDCx6p67_ASAP7_75t_R g291 ( 
.A(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_170),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_226),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_227),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_257),
.B(n_212),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_173),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_238),
.B1(n_251),
.B2(n_222),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_228),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_278),
.B(n_175),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_238),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_278),
.B(n_271),
.Y(n_313)
);

O2A1O1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_252),
.B(n_237),
.C(n_232),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_252),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_182),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_229),
.B(n_232),
.C(n_236),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_236),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_237),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_242),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_265),
.B(n_189),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_254),
.B(n_242),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_291),
.A2(n_222),
.B1(n_221),
.B2(n_223),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_254),
.B(n_241),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_265),
.B(n_193),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

AO221x1_ASAP7_75t_L g339 ( 
.A1(n_265),
.A2(n_241),
.B1(n_244),
.B2(n_240),
.C(n_230),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_289),
.Y(n_340)
);

AND2x6_ASAP7_75t_SL g341 ( 
.A(n_291),
.B(n_214),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_241),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_280),
.A2(n_223),
.B1(n_247),
.B2(n_244),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_240),
.B(n_244),
.C(n_211),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_285),
.A2(n_247),
.B1(n_223),
.B2(n_250),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_286),
.B(n_230),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_263),
.B(n_201),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

OAI221xp5_ASAP7_75t_L g355 ( 
.A1(n_285),
.A2(n_159),
.B1(n_197),
.B2(n_223),
.C(n_247),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_268),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_269),
.A2(n_276),
.B1(n_204),
.B2(n_247),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_255),
.B(n_273),
.Y(n_360)
);

OR2x6_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_214),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_270),
.Y(n_363)
);

AO32x2_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_250),
.A3(n_230),
.B1(n_239),
.B2(n_11),
.Y(n_364)
);

O2A1O1Ixp5_ASAP7_75t_L g365 ( 
.A1(n_302),
.A2(n_279),
.B(n_277),
.C(n_272),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_281),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_307),
.A2(n_281),
.B(n_279),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_277),
.B(n_272),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_317),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_298),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_308),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_313),
.A2(n_299),
.B(n_294),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_317),
.A2(n_234),
.B(n_215),
.C(n_224),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_313),
.A2(n_234),
.B(n_215),
.C(n_224),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_299),
.B(n_294),
.Y(n_378)
);

INVx11_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_315),
.B(n_250),
.C(n_230),
.Y(n_381)
);

A2O1A1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_315),
.A2(n_233),
.B(n_211),
.C(n_250),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_239),
.B1(n_269),
.B2(n_276),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_301),
.Y(n_384)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_314),
.A2(n_312),
.B(n_316),
.C(n_319),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_340),
.A2(n_233),
.B(n_250),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_230),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_333),
.B(n_276),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_239),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_239),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_333),
.B(n_8),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_80),
.B(n_150),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_341),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_311),
.A2(n_79),
.B(n_149),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_336),
.A2(n_78),
.B(n_148),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_22),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_400)
);

BUFx8_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_305),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_23),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_353),
.A2(n_82),
.B(n_147),
.Y(n_405)
);

BUFx4f_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_353),
.A2(n_81),
.B(n_144),
.Y(n_407)
);

AOI21xp33_ASAP7_75t_L g408 ( 
.A1(n_312),
.A2(n_10),
.B(n_12),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_304),
.B(n_12),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_348),
.A2(n_84),
.B(n_143),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_348),
.A2(n_77),
.B(n_141),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_362),
.B(n_334),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_303),
.A2(n_74),
.B(n_140),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_352),
.B(n_13),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_345),
.A2(n_72),
.B(n_139),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_352),
.A2(n_67),
.B(n_138),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_344),
.A2(n_65),
.B(n_137),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_330),
.B(n_13),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_361),
.B(n_14),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_330),
.A2(n_85),
.B(n_134),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_344),
.A2(n_64),
.B(n_133),
.Y(n_425)
);

A2O1A1Ixp33_ASAP7_75t_L g426 ( 
.A1(n_323),
.A2(n_320),
.B(n_321),
.C(n_356),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_337),
.B(n_15),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_337),
.A2(n_63),
.B(n_132),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_350),
.A2(n_62),
.B(n_131),
.Y(n_429)
);

AO22x1_ASAP7_75t_L g430 ( 
.A1(n_354),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_342),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_365),
.A2(n_368),
.B(n_414),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_305),
.B(n_318),
.Y(n_434)
);

AOI21x1_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_363),
.B(n_358),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_371),
.B(n_305),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_394),
.B(n_305),
.Y(n_437)
);

O2A1O1Ixp5_ASAP7_75t_L g438 ( 
.A1(n_418),
.A2(n_351),
.B(n_29),
.C(n_30),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_351),
.B(n_31),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_375),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_90),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_17),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_370),
.B(n_366),
.Y(n_443)
);

INVx3_ASAP7_75t_SL g444 ( 
.A(n_396),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_33),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_34),
.B(n_35),
.Y(n_446)
);

AOI31xp67_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_36),
.A3(n_38),
.B(n_39),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_374),
.A2(n_40),
.B(n_41),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

BUFx12f_ASAP7_75t_L g451 ( 
.A(n_401),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_420),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_48),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_391),
.B(n_49),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_367),
.A2(n_152),
.B(n_52),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_381),
.B(n_51),
.Y(n_456)
);

HAxp5_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_401),
.CON(n_457),
.SN(n_457)
);

NAND3xp33_ASAP7_75t_SL g458 ( 
.A(n_400),
.B(n_56),
.C(n_57),
.Y(n_458)
);

AOI221x1_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.C(n_87),
.Y(n_459)
);

AOI221x1_ASAP7_75t_L g460 ( 
.A1(n_385),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_378),
.A2(n_95),
.B(n_96),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_98),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_99),
.C(n_100),
.Y(n_463)
);

CKINVDCx8_ASAP7_75t_R g464 ( 
.A(n_379),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_406),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_402),
.A2(n_101),
.B(n_102),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_103),
.C(n_104),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_409),
.B(n_105),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_426),
.A2(n_108),
.B(n_110),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_403),
.A2(n_123),
.B(n_124),
.Y(n_473)
);

AOI221xp5_ASAP7_75t_SL g474 ( 
.A1(n_376),
.A2(n_377),
.B1(n_382),
.B2(n_408),
.C(n_427),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_410),
.A2(n_127),
.B(n_128),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_129),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_413),
.Y(n_477)
);

AOI21xp33_ASAP7_75t_L g478 ( 
.A1(n_421),
.A2(n_400),
.B(n_381),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_386),
.A2(n_424),
.B(n_383),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_422),
.Y(n_482)
);

AO31x2_ASAP7_75t_L g483 ( 
.A1(n_364),
.A2(n_416),
.A3(n_419),
.B(n_428),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_423),
.A2(n_405),
.B(n_407),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_430),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_435),
.A2(n_395),
.B(n_429),
.Y(n_487)
);

OAI21x1_ASAP7_75t_SL g488 ( 
.A1(n_452),
.A2(n_364),
.B(n_454),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_432),
.B(n_482),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_433),
.A2(n_485),
.B(n_480),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_431),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

NAND2x1p5_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_470),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_441),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_484),
.B(n_439),
.Y(n_497)
);

AO21x2_ASAP7_75t_L g498 ( 
.A1(n_462),
.A2(n_471),
.B(n_478),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_468),
.A2(n_452),
.B1(n_459),
.B2(n_458),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_469),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_456),
.B(n_461),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_445),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_468),
.B(n_436),
.Y(n_503)
);

NOR2x1_ASAP7_75t_R g504 ( 
.A(n_451),
.B(n_465),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_453),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_470),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_440),
.B(n_457),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

BUFx5_ASAP7_75t_L g512 ( 
.A(n_447),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_484),
.A2(n_438),
.B(n_446),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_448),
.A2(n_475),
.B(n_455),
.Y(n_514)
);

AOI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_444),
.A2(n_463),
.B(n_467),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_456),
.A2(n_437),
.B(n_476),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_483),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_466),
.B(n_460),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_479),
.A2(n_435),
.B(n_462),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_433),
.A2(n_425),
.B(n_420),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_469),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_468),
.A2(n_400),
.B1(n_213),
.B2(n_452),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_433),
.A2(n_435),
.B(n_485),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_433),
.A2(n_435),
.B(n_485),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_438),
.A2(n_425),
.B(n_420),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_449),
.B(n_470),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_443),
.B(n_369),
.Y(n_532)
);

OA21x2_ASAP7_75t_L g533 ( 
.A1(n_433),
.A2(n_425),
.B(n_420),
.Y(n_533)
);

CKINVDCx6p67_ASAP7_75t_R g534 ( 
.A(n_444),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_495),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_494),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_492),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_525),
.A2(n_526),
.B(n_528),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_524),
.B1(n_499),
.B2(n_528),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_523),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_500),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_496),
.B(n_502),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_508),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_495),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_486),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_514),
.A2(n_497),
.B(n_491),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_513),
.A2(n_520),
.B(n_487),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_493),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_534),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_490),
.B(n_496),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_502),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_490),
.B(n_524),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_531),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_529),
.A2(n_518),
.B(n_488),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_529),
.A2(n_519),
.B(n_517),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_507),
.B(n_511),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_495),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_507),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_517),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_499),
.A2(n_533),
.B(n_522),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_530),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_506),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_515),
.B(n_533),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_516),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_516),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_501),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_510),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_522),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_559),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_564),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_536),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_498),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_559),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_498),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_509),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_512),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_547),
.B(n_512),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_546),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_547),
.B(n_504),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_558),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_538),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_558),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_553),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_567),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_512),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_567),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_542),
.B(n_512),
.Y(n_596)
);

NOR2x1_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_512),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_576),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_512),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_540),
.A2(n_554),
.B1(n_544),
.B2(n_565),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_541),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_543),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_573),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_574),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_544),
.A2(n_554),
.B1(n_571),
.B2(n_545),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_569),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_566),
.B(n_557),
.Y(n_612)
);

AND2x4_ASAP7_75t_SL g613 ( 
.A(n_546),
.B(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_572),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_572),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_566),
.B(n_537),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_535),
.B(n_562),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_550),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_579),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_537),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_614),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_581),
.B(n_579),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_590),
.B(n_570),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_614),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_603),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_605),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_596),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_581),
.B(n_539),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_605),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_587),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_590),
.B(n_546),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_577),
.B(n_539),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_596),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_539),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_577),
.B(n_550),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_616),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_580),
.B(n_546),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_598),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_610),
.B(n_546),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_549),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_608),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_588),
.B(n_552),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_617),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_604),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_584),
.B(n_535),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_584),
.A2(n_552),
.B1(n_562),
.B2(n_549),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_608),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_585),
.B(n_583),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_615),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_630),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_630),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_655),
.B(n_592),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_647),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_621),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_625),
.B(n_599),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_625),
.B(n_599),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_578),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_655),
.B(n_585),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_633),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_633),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_615),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_624),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_632),
.B(n_578),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_641),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_624),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_632),
.B(n_582),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_646),
.B(n_582),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_653),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_628),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_646),
.B(n_591),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_643),
.B(n_594),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_591),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_637),
.B(n_589),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_601),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_638),
.B(n_601),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_637),
.B(n_620),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_660),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_665),
.B(n_627),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_657),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_662),
.B(n_627),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_679),
.B(n_622),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_665),
.B(n_654),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_663),
.B(n_648),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_649),
.Y(n_692)
);

AOI32xp33_ASAP7_75t_L g693 ( 
.A1(n_659),
.A2(n_652),
.A3(n_674),
.B1(n_651),
.B2(n_678),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_659),
.B(n_638),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_664),
.B(n_656),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_661),
.B(n_641),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_674),
.B(n_640),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_675),
.A2(n_602),
.B1(n_609),
.B2(n_611),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_641),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_658),
.Y(n_700)
);

OAI21xp33_ASAP7_75t_L g701 ( 
.A1(n_676),
.A2(n_626),
.B(n_635),
.Y(n_701)
);

NOR2x1p5_ASAP7_75t_L g702 ( 
.A(n_671),
.B(n_642),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_664),
.B(n_656),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_686),
.B(n_673),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_689),
.B(n_673),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_699),
.B(n_670),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_685),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_694),
.B(n_670),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_687),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_698),
.A2(n_593),
.B(n_595),
.C(n_618),
.Y(n_710)
);

OAI222xp33_ASAP7_75t_L g711 ( 
.A1(n_693),
.A2(n_649),
.B1(n_680),
.B2(n_684),
.C1(n_681),
.C2(n_644),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_688),
.B(n_684),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_SL g713 ( 
.A(n_702),
.B(n_593),
.Y(n_713)
);

AOI21xp33_ASAP7_75t_L g714 ( 
.A1(n_710),
.A2(n_701),
.B(n_691),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_709),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_705),
.A2(n_701),
.B(n_690),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_711),
.A2(n_698),
.B(n_692),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_707),
.Y(n_718)
);

OAI211xp5_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_700),
.B(n_697),
.C(n_696),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_707),
.Y(n_720)
);

OAI221xp5_ASAP7_75t_SL g721 ( 
.A1(n_719),
.A2(n_692),
.B1(n_712),
.B2(n_711),
.C(n_703),
.Y(n_721)
);

OAI32xp33_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_713),
.A3(n_695),
.B1(n_681),
.B2(n_680),
.Y(n_722)
);

AOI221xp5_ASAP7_75t_L g723 ( 
.A1(n_714),
.A2(n_704),
.B1(n_666),
.B2(n_667),
.C(n_706),
.Y(n_723)
);

AOI221xp5_ASAP7_75t_L g724 ( 
.A1(n_717),
.A2(n_672),
.B1(n_669),
.B2(n_678),
.C(n_595),
.Y(n_724)
);

AOI211xp5_ASAP7_75t_L g725 ( 
.A1(n_716),
.A2(n_715),
.B(n_720),
.C(n_718),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_714),
.B(n_677),
.C(n_634),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_725),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_723),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_721),
.B(n_726),
.C(n_722),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_724),
.B(n_677),
.C(n_634),
.Y(n_730)
);

NAND4xp25_ASAP7_75t_L g731 ( 
.A(n_727),
.B(n_610),
.C(n_645),
.D(n_623),
.Y(n_731)
);

AND3x2_ASAP7_75t_L g732 ( 
.A(n_729),
.B(n_617),
.C(n_645),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_728),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_733),
.Y(n_734)
);

NOR2x1_ASAP7_75t_L g735 ( 
.A(n_731),
.B(n_730),
.Y(n_735)
);

NOR3x1_ASAP7_75t_L g736 ( 
.A(n_732),
.B(n_629),
.C(n_636),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_SL g737 ( 
.A1(n_735),
.A2(n_708),
.B(n_692),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_734),
.A2(n_677),
.B1(n_649),
.B2(n_645),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_736),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_734),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_734),
.Y(n_741)
);

INVxp33_ASAP7_75t_SL g742 ( 
.A(n_734),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_741),
.B(n_683),
.Y(n_743)
);

XNOR2x1_ASAP7_75t_L g744 ( 
.A(n_739),
.B(n_587),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_683),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

OAI22x1_ASAP7_75t_L g747 ( 
.A1(n_737),
.A2(n_623),
.B1(n_671),
.B2(n_619),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_746),
.B(n_738),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_SL g749 ( 
.A1(n_743),
.A2(n_587),
.B1(n_623),
.B2(n_650),
.Y(n_749)
);

NAND4xp25_ASAP7_75t_L g750 ( 
.A(n_745),
.B(n_612),
.C(n_616),
.D(n_671),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_SL g751 ( 
.A1(n_744),
.A2(n_587),
.B(n_607),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_748),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_SL g753 ( 
.A1(n_749),
.A2(n_747),
.B1(n_607),
.B2(n_616),
.Y(n_753)
);

XNOR2xp5_ASAP7_75t_L g754 ( 
.A(n_750),
.B(n_613),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_752),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_754),
.Y(n_756)
);

OAI22x1_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_751),
.B1(n_616),
.B2(n_660),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_755),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_758),
.B(n_756),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_759),
.B(n_757),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_613),
.B(n_612),
.Y(n_761)
);


endmodule