module fake_netlist_6_1086_n_1700 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1700);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1700;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_2),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_4),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_80),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_34),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_81),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_33),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_15),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_70),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_35),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_58),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_23),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_3),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_60),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_31),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_47),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_83),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_29),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_113),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_149),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_2),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_67),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_30),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_116),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_85),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_74),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_6),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_8),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_44),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_120),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_59),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_66),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_134),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_20),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_135),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_11),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_111),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_118),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_51),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_105),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_123),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_55),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_106),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_61),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_57),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_131),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_52),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_128),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_126),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_26),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_49),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_32),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_91),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_137),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_92),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_148),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_146),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_100),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_121),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_19),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_71),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_97),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_139),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_76),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_42),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_33),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_140),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_54),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_98),
.Y(n_292)
);

BUFx2_ASAP7_75t_SL g293 ( 
.A(n_75),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_65),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_64),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_125),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_110),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_7),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_99),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_142),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_133),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_13),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_28),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_10),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_198),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_173),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_199),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_176),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_200),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_219),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_209),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_203),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_195),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_205),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_263),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_182),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_269),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_208),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_210),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_165),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_211),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_181),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_213),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_186),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_191),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_222),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_194),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_157),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_215),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_217),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_218),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_220),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_157),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_231),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_264),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_224),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_268),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g363 ( 
.A(n_160),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_235),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_160),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_163),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_225),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_227),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_236),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_182),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_249),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_278),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_174),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_174),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_196),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_196),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_237),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_197),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_163),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_312),
.B(n_262),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_311),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_317),
.B(n_262),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_296),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_305),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_313),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_314),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_322),
.B(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_296),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

CKINVDCx11_ASAP7_75t_R g404 ( 
.A(n_315),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_204),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_293),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_335),
.B(n_204),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_318),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_330),
.B(n_182),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_324),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_159),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_158),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_334),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_226),
.B(n_216),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_380),
.B(n_156),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_380),
.B(n_335),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_325),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_337),
.B(n_156),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_337),
.B(n_161),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_342),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_345),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_345),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_319),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_362),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_383),
.A2(n_226),
.B(n_216),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_446),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_326),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_386),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_338),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_446),
.Y(n_461)
);

OAI22x1_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_352),
.B1(n_358),
.B2(n_188),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_416),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_340),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_385),
.B(n_360),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_399),
.B(n_344),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_398),
.B(n_360),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_421),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_406),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_419),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_382),
.B(n_285),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_394),
.B(n_336),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_429),
.A2(n_266),
.B1(n_179),
.B2(n_248),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_343),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_414),
.B(n_347),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_408),
.A2(n_358),
.B1(n_339),
.B2(n_374),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_422),
.B(n_350),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx8_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_430),
.A2(n_363),
.B1(n_169),
.B2(n_177),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_412),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_429),
.B(n_367),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_408),
.B(n_285),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_413),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_SL g503 ( 
.A(n_439),
.B(n_361),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_436),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_439),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_382),
.A2(n_295),
.B1(n_376),
.B2(n_354),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_382),
.A2(n_295),
.B1(n_182),
.B2(n_372),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_389),
.B(n_346),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_426),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_440),
.B(n_369),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_411),
.A2(n_182),
.B1(n_373),
.B2(n_372),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_389),
.B(n_346),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_411),
.A2(n_348),
.B1(n_373),
.B2(n_371),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_393),
.B(n_379),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_384),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_389),
.B(n_348),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_428),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_368),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

BUFx6f_ASAP7_75t_SL g533 ( 
.A(n_442),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_384),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_401),
.B(n_170),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_441),
.B(n_162),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_401),
.B(n_238),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_409),
.B(n_168),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_411),
.A2(n_371),
.B1(n_364),
.B2(n_359),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_409),
.B(n_241),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_427),
.B(n_242),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_393),
.B(n_161),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_387),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_420),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_430),
.A2(n_228),
.B1(n_193),
.B2(n_202),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_387),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_387),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_438),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_441),
.B(n_364),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_427),
.B(n_251),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_391),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_427),
.B(n_254),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_416),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_403),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_434),
.B(n_359),
.C(n_357),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_391),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_427),
.B(n_259),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_397),
.A2(n_289),
.B1(n_309),
.B2(n_308),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_428),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_428),
.Y(n_567)
);

BUFx6f_ASAP7_75t_SL g568 ( 
.A(n_442),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_396),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_396),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_396),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_404),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_434),
.B(n_164),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_403),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_444),
.B(n_164),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_405),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_405),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_435),
.B(n_349),
.Y(n_581)
);

BUFx4f_ASAP7_75t_L g582 ( 
.A(n_420),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_383),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_443),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_431),
.B(n_349),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_444),
.B(n_166),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_418),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_418),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_427),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_461),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_470),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_453),
.B(n_166),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_471),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_461),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_553),
.B(n_172),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_467),
.B(n_234),
.C(n_201),
.Y(n_602)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_492),
.B(n_445),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_539),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_553),
.B(n_175),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_452),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_459),
.B(n_167),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_388),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_581),
.A2(n_388),
.B(n_390),
.C(n_432),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_543),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_584),
.B(n_167),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_390),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_447),
.B(n_183),
.Y(n_613)
);

INVxp33_ASAP7_75t_L g614 ( 
.A(n_486),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_464),
.B(n_178),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_169),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_403),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_531),
.B(n_178),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_591),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_447),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_180),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_475),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_475),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_447),
.B(n_190),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_535),
.B(n_180),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_463),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_558),
.B(n_169),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_533),
.B(n_188),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_448),
.B(n_454),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_448),
.B(n_454),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_458),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_477),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_455),
.B(n_395),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_477),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_487),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_543),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_455),
.B(n_395),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_536),
.B(n_184),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_458),
.B(n_192),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_457),
.B(n_472),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_184),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_487),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_457),
.B(n_395),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_587),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_496),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_515),
.B(n_351),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_587),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_495),
.B(n_206),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_496),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_472),
.B(n_395),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_504),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_533),
.A2(n_177),
.B1(n_272),
.B2(n_288),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_515),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_536),
.A2(n_267),
.B1(n_247),
.B2(n_240),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_497),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_473),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_473),
.Y(n_661)
);

BUFx8_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_514),
.B(n_207),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_514),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_560),
.B(n_488),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_497),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_482),
.B(n_425),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_482),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_537),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_491),
.B(n_493),
.Y(n_670)
);

BUFx8_ASAP7_75t_L g671 ( 
.A(n_576),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_514),
.B(n_232),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_500),
.A2(n_252),
.B1(n_256),
.B2(n_260),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_489),
.B(n_351),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_581),
.B(n_507),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_536),
.B(n_189),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_353),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_501),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_514),
.B(n_261),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_510),
.B(n_425),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_521),
.B(n_353),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_528),
.B(n_356),
.Y(n_682)
);

AO221x1_ASAP7_75t_L g683 ( 
.A1(n_462),
.A2(n_302),
.B1(n_276),
.B2(n_290),
.C(n_292),
.Y(n_683)
);

INVx8_ASAP7_75t_L g684 ( 
.A(n_533),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_510),
.B(n_418),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_568),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_511),
.B(n_431),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_500),
.B(n_265),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_560),
.B(n_432),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_582),
.B(n_479),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_574),
.B(n_189),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_511),
.B(n_271),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_463),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_512),
.B(n_274),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_500),
.A2(n_272),
.B1(n_288),
.B2(n_301),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_503),
.B(n_404),
.C(n_356),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_512),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_479),
.A2(n_500),
.B1(n_528),
.B2(n_568),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_516),
.B(n_274),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_514),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_523),
.B(n_275),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_517),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_541),
.B(n_275),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_501),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_479),
.B(n_277),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_479),
.B(n_277),
.Y(n_708)
);

OAI22x1_ASAP7_75t_SL g709 ( 
.A1(n_573),
.A2(n_309),
.B1(n_308),
.B2(n_306),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_543),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_559),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_502),
.Y(n_712)
);

BUFx8_ASAP7_75t_L g713 ( 
.A(n_568),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_486),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_559),
.B(n_279),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_559),
.B(n_280),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_502),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_571),
.B(n_280),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_480),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_523),
.B(n_281),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_571),
.B(n_281),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_523),
.B(n_282),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_506),
.B(n_357),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_523),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_523),
.B(n_282),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_505),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_577),
.B(n_588),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_582),
.B(n_284),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_505),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_571),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_513),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_513),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_520),
.A2(n_286),
.B(n_307),
.C(n_287),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_500),
.A2(n_301),
.B1(n_306),
.B2(n_212),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_524),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_506),
.B(n_304),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_583),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_506),
.B(n_233),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_506),
.B(n_230),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_583),
.B(n_297),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_500),
.A2(n_257),
.B1(n_221),
.B2(n_229),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_582),
.B(n_286),
.Y(n_743)
);

INVx8_ASAP7_75t_L g744 ( 
.A(n_494),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_520),
.A2(n_554),
.B(n_542),
.C(n_557),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_547),
.B(n_304),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_529),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_529),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_569),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_532),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_480),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_538),
.B(n_299),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_538),
.B(n_298),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_544),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_465),
.B(n_214),
.C(n_239),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_562),
.B(n_508),
.Y(n_756)
);

AND2x4_ASAP7_75t_SL g757 ( 
.A(n_655),
.B(n_483),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_596),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_665),
.B(n_603),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_664),
.B(n_550),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_723),
.B(n_563),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_598),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_598),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_719),
.A2(n_483),
.B1(n_573),
.B2(n_563),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_595),
.B(n_600),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_664),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_597),
.B(n_468),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_599),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_597),
.B(n_526),
.Y(n_769)
);

AO22x1_ASAP7_75t_L g770 ( 
.A1(n_618),
.A2(n_538),
.B1(n_255),
.B2(n_253),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_599),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_657),
.B(n_519),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_664),
.B(n_550),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_618),
.B(n_575),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_621),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_622),
.B(n_575),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_627),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_664),
.B(n_556),
.Y(n_778)
);

AND2x2_ASAP7_75t_SL g779 ( 
.A(n_695),
.B(n_522),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_700),
.B(n_556),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_700),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_606),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_623),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_700),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_624),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_624),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_700),
.B(n_565),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_693),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_724),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_657),
.B(n_575),
.Y(n_790)
);

NOR2x2_ASAP7_75t_L g791 ( 
.A(n_652),
.B(n_462),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_724),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_634),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_634),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_635),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_724),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_575),
.Y(n_797)
);

BUFx5_ASAP7_75t_L g798 ( 
.A(n_690),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_635),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_684),
.B(n_686),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

AO22x1_ASAP7_75t_L g802 ( 
.A1(n_746),
.A2(n_538),
.B1(n_244),
.B2(n_246),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_669),
.A2(n_538),
.B1(n_579),
.B2(n_586),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_754),
.B(n_287),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_724),
.B(n_565),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_620),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_674),
.A2(n_250),
.B1(n_258),
.B2(n_538),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_638),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_638),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_620),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_639),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_639),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_604),
.B(n_540),
.Y(n_813)
);

BUFx8_ASAP7_75t_L g814 ( 
.A(n_628),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_646),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_616),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_650),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_675),
.B(n_579),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_669),
.B(n_585),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_607),
.B(n_291),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_649),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_611),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_690),
.B(n_546),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_711),
.B(n_585),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_684),
.B(n_686),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_649),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_653),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_650),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_615),
.A2(n_538),
.B1(n_586),
.B2(n_494),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_663),
.A2(n_450),
.B(n_590),
.C(n_589),
.Y(n_831)
);

AO22x1_ASAP7_75t_L g832 ( 
.A1(n_746),
.A2(n_297),
.B1(n_294),
.B2(n_291),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_610),
.B(n_294),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_677),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_653),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_659),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_648),
.B(n_564),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_738),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_677),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_681),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_659),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_666),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_608),
.B(n_593),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_666),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_682),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_615),
.B(n_546),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_678),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_662),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_611),
.B(n_451),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_727),
.B(n_546),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_651),
.B(n_564),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_678),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_712),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_671),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_SL g855 ( 
.A(n_684),
.B(n_494),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_712),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_612),
.B(n_570),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_695),
.A2(n_494),
.B1(n_469),
.B2(n_466),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_671),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_633),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_726),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_601),
.A2(n_605),
.B(n_725),
.C(n_720),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_631),
.B(n_570),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_714),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_632),
.B(n_593),
.Y(n_865)
);

OR2x6_ASAP7_75t_L g866 ( 
.A(n_686),
.B(n_494),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_735),
.A2(n_456),
.B1(n_466),
.B2(n_469),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_727),
.A2(n_566),
.B1(n_567),
.B2(n_481),
.Y(n_868)
);

INVx5_ASAP7_75t_L g869 ( 
.A(n_744),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_726),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_644),
.B(n_572),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_670),
.B(n_572),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_SL g873 ( 
.A(n_691),
.B(n_456),
.C(n_590),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_713),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_732),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_689),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_732),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_619),
.B(n_578),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_660),
.B(n_578),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_706),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_739),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_626),
.B(n_546),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_717),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_734),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_633),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_729),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_731),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_661),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_740),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_668),
.B(n_580),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_629),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_R g892 ( 
.A(n_630),
.B(n_450),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_735),
.A2(n_742),
.B1(n_676),
.B2(n_642),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_626),
.B(n_580),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_698),
.B(n_566),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_745),
.A2(n_567),
.B(n_481),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_697),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_701),
.B(n_703),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_749),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_704),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_594),
.B(n_589),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_640),
.B(n_530),
.Y(n_902)
);

AND2x2_ASAP7_75t_SL g903 ( 
.A(n_696),
.B(n_530),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_736),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_702),
.A2(n_474),
.B1(n_481),
.B2(n_460),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_609),
.B(n_499),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_749),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_747),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_702),
.A2(n_499),
.B1(n_474),
.B2(n_460),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_751),
.B(n_0),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_710),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_748),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_750),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_614),
.B(n_0),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_601),
.B(n_499),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_605),
.B(n_687),
.Y(n_916)
);

NOR2x2_ASAP7_75t_L g917 ( 
.A(n_656),
.B(n_7),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_685),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_642),
.A2(n_645),
.B1(n_676),
.B2(n_755),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_637),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_602),
.B(n_451),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_645),
.B(n_592),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_737),
.B(n_451),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_756),
.B(n_663),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_672),
.B(n_474),
.Y(n_925)
);

NOR2x2_ASAP7_75t_L g926 ( 
.A(n_709),
.B(n_9),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_694),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_641),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_744),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_672),
.B(n_460),
.Y(n_930)
);

OR2x2_ASAP7_75t_SL g931 ( 
.A(n_914),
.B(n_713),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_860),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_792),
.A2(n_744),
.B(n_679),
.Y(n_933)
);

BUFx4f_ASAP7_75t_L g934 ( 
.A(n_826),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_840),
.B(n_699),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_777),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_893),
.A2(n_679),
.B1(n_715),
.B2(n_741),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_792),
.A2(n_797),
.B(n_776),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_SL g939 ( 
.A(n_769),
.B(n_691),
.C(n_733),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_782),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_758),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_888),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_823),
.B(n_705),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_924),
.A2(n_720),
.B(n_722),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_862),
.A2(n_725),
.B(n_722),
.C(n_708),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_821),
.A2(n_658),
.B(n_692),
.C(n_625),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_774),
.A2(n_721),
.B1(n_716),
.B2(n_718),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_862),
.A2(n_707),
.B(n_643),
.C(n_613),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_829),
.B(n_613),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_792),
.A2(n_688),
.B(n_673),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_779),
.A2(n_743),
.B1(n_728),
.B2(n_625),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_834),
.B(n_643),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_916),
.A2(n_743),
.B1(n_728),
.B2(n_617),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_839),
.B(n_654),
.Y(n_955)
);

BUFx12f_ASAP7_75t_L g956 ( 
.A(n_854),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_761),
.A2(n_680),
.B(n_667),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_864),
.B(n_647),
.Y(n_958)
);

OAI22xp33_ASAP7_75t_L g959 ( 
.A1(n_845),
.A2(n_683),
.B1(n_752),
.B2(n_753),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_478),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_927),
.B(n_561),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_881),
.B(n_816),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_860),
.B(n_478),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_762),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_916),
.A2(n_478),
.B1(n_484),
.B2(n_485),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_788),
.B(n_478),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_885),
.B(n_484),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_814),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_792),
.A2(n_490),
.B(n_485),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_924),
.A2(n_484),
.B1(n_485),
.B2(n_490),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_766),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_901),
.A2(n_490),
.B(n_509),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_889),
.B(n_525),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_901),
.A2(n_509),
.B(n_530),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_846),
.A2(n_545),
.B(n_561),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_800),
.B(n_82),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_814),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_838),
.A2(n_509),
.B1(n_530),
.B2(n_525),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_L g979 ( 
.A1(n_807),
.A2(n_527),
.B(n_534),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_763),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_817),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_918),
.B(n_527),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_929),
.B(n_509),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_813),
.B(n_534),
.Y(n_984)
);

AND2x2_ASAP7_75t_SL g985 ( 
.A(n_757),
.B(n_9),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_781),
.Y(n_986)
);

O2A1O1Ixp5_ASAP7_75t_L g987 ( 
.A1(n_759),
.A2(n_548),
.B(n_555),
.C(n_551),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_897),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_838),
.A2(n_592),
.B(n_546),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_760),
.A2(n_552),
.B(n_546),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_813),
.B(n_555),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_832),
.A2(n_548),
.B1(n_549),
.B2(n_551),
.C(n_20),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_11),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_898),
.B(n_843),
.Y(n_994)
);

INVx5_ASAP7_75t_L g995 ( 
.A(n_826),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_900),
.Y(n_996)
);

AO32x1_ASAP7_75t_L g997 ( 
.A1(n_894),
.A2(n_12),
.A3(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_910),
.B(n_12),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_781),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_848),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_791),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_911),
.B(n_21),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_843),
.B(n_22),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_849),
.B(n_24),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_859),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_807),
.A2(n_552),
.B(n_25),
.C(n_26),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_765),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_798),
.B(n_552),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_781),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_802),
.B(n_552),
.C(n_27),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_826),
.B(n_62),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_904),
.B(n_908),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_820),
.A2(n_552),
.B1(n_73),
.B2(n_87),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_874),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_784),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_912),
.B(n_24),
.Y(n_1016)
);

AOI22x1_ASAP7_75t_L g1017 ( 
.A1(n_920),
.A2(n_420),
.B1(n_56),
.B2(n_147),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_772),
.A2(n_420),
.B1(n_552),
.B2(n_32),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_820),
.A2(n_48),
.B1(n_132),
.B2(n_130),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_928),
.B(n_28),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_919),
.A2(n_420),
.B1(n_46),
.B2(n_89),
.Y(n_1021)
);

OAI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_764),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.C(n_40),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_760),
.A2(n_420),
.B(n_102),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_857),
.B(n_36),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_784),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_806),
.A2(n_119),
.B1(n_127),
.B2(n_124),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_911),
.B(n_41),
.Y(n_1027)
);

AO32x2_ASAP7_75t_L g1028 ( 
.A1(n_896),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_90),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_768),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_911),
.B(n_45),
.Y(n_1030)
);

OAI22x1_ASAP7_75t_L g1031 ( 
.A1(n_917),
.A2(n_420),
.B1(n_810),
.B2(n_806),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_771),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_773),
.A2(n_780),
.B(n_787),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_810),
.A2(n_913),
.B1(n_906),
.B2(n_858),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_866),
.B(n_891),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_837),
.B(n_851),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_837),
.B(n_851),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_880),
.B(n_883),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_863),
.B(n_865),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_784),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_863),
.B(n_865),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_789),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_789),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_773),
.A2(n_805),
.B(n_787),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_798),
.B(n_891),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_871),
.B(n_872),
.Y(n_1046)
);

AO32x2_ASAP7_75t_L g1047 ( 
.A1(n_896),
.A2(n_873),
.A3(n_906),
.B1(n_895),
.B2(n_892),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_886),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_775),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_789),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_887),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_804),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_884),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_830),
.A2(n_825),
.B1(n_778),
.B2(n_805),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_833),
.B(n_770),
.C(n_790),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_866),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_818),
.A2(n_915),
.B(n_890),
.C(n_878),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_818),
.A2(n_800),
.B(n_923),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_825),
.B(n_785),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_944),
.A2(n_831),
.B(n_803),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1038),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_942),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_975),
.A2(n_831),
.B(n_780),
.Y(n_1063)
);

AOI221x1_ASAP7_75t_L g1064 ( 
.A1(n_939),
.A2(n_873),
.B1(n_921),
.B2(n_778),
.C(n_930),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_994),
.B(n_798),
.Y(n_1065)
);

AOI221x1_ASAP7_75t_L g1066 ( 
.A1(n_952),
.A2(n_930),
.B1(n_925),
.B2(n_915),
.C(n_878),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_1004),
.A2(n_882),
.B(n_922),
.C(n_850),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_972),
.A2(n_929),
.B(n_890),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1039),
.B(n_798),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_974),
.A2(n_879),
.B(n_842),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_946),
.A2(n_903),
.B(n_868),
.C(n_879),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_988),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_945),
.A2(n_867),
.B(n_905),
.Y(n_1073)
);

AOI21x1_ASAP7_75t_L g1074 ( 
.A1(n_938),
.A2(n_902),
.B(n_835),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_947),
.A2(n_869),
.B(n_796),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1041),
.B(n_798),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_996),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_937),
.A2(n_909),
.B(n_895),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1012),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_954),
.A2(n_895),
.B(n_877),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_995),
.B(n_866),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_943),
.A2(n_895),
.B1(n_902),
.B2(n_855),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1029),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_SL g1084 ( 
.A(n_1022),
.B(n_926),
.C(n_809),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1032),
.Y(n_1085)
);

OAI22x1_ASAP7_75t_L g1086 ( 
.A1(n_1021),
.A2(n_875),
.B1(n_861),
.B2(n_793),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_985),
.B(n_783),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1033),
.A2(n_1044),
.B(n_987),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_1056),
.B(n_869),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1046),
.A2(n_869),
.B(n_855),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_935),
.B(n_907),
.Y(n_1091)
);

CKINVDCx16_ASAP7_75t_R g1092 ( 
.A(n_1014),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_951),
.A2(n_856),
.B(n_853),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_957),
.A2(n_822),
.B(n_852),
.C(n_795),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_998),
.B(n_786),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_959),
.A2(n_1024),
.B(n_949),
.C(n_1003),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_995),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_933),
.A2(n_815),
.B(n_847),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_SL g1099 ( 
.A1(n_1019),
.A2(n_1045),
.B(n_1013),
.C(n_1054),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1057),
.A2(n_796),
.B(n_902),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_969),
.A2(n_812),
.B(n_799),
.Y(n_1101)
);

NOR2x1_ASAP7_75t_L g1102 ( 
.A(n_936),
.B(n_1015),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_968),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1056),
.Y(n_1104)
);

INVx3_ASAP7_75t_SL g1105 ( 
.A(n_977),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1059),
.B(n_808),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_970),
.A2(n_794),
.B(n_801),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_983),
.A2(n_811),
.B(n_819),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1000),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1034),
.A2(n_841),
.B(n_827),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1058),
.A2(n_828),
.B(n_836),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_981),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_995),
.B(n_899),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_958),
.B(n_1001),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1056),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1048),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_1027),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1036),
.B(n_870),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_SL g1119 ( 
.A1(n_963),
.A2(n_824),
.B(n_844),
.C(n_967),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_965),
.A2(n_978),
.A3(n_1006),
.B(n_960),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_984),
.B(n_991),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_982),
.B(n_1020),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_962),
.B(n_1051),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1021),
.A2(n_1018),
.B1(n_1035),
.B2(n_1016),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1008),
.A2(n_979),
.B(n_989),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_950),
.B(n_953),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1055),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_983),
.A2(n_990),
.B(n_1017),
.Y(n_1128)
);

AOI22x1_ASAP7_75t_L g1129 ( 
.A1(n_1031),
.A2(n_980),
.B1(n_1049),
.B2(n_964),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_955),
.B(n_941),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_956),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_955),
.B(n_961),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1007),
.B(n_1052),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1011),
.B(n_948),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_971),
.A2(n_1043),
.B(n_986),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_950),
.A2(n_953),
.B(n_992),
.C(n_993),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_986),
.A2(n_1043),
.B(n_1026),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_966),
.A2(n_1053),
.B(n_1002),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1030),
.A2(n_934),
.B(n_1047),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1047),
.A2(n_1011),
.B(n_934),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_999),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_1005),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1047),
.A2(n_1028),
.A3(n_997),
.B(n_1015),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_940),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_999),
.A2(n_1009),
.B(n_1042),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_976),
.A2(n_1028),
.B(n_1050),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_932),
.B(n_948),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_1025),
.B(n_1042),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1009),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_997),
.A2(n_1050),
.B(n_1009),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1025),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_948),
.B(n_1025),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_SL g1153 ( 
.A1(n_1028),
.A2(n_997),
.B(n_931),
.Y(n_1153)
);

NAND3x1_ASAP7_75t_L g1154 ( 
.A(n_1040),
.B(n_1042),
.C(n_1050),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_1040),
.A2(n_769),
.B(n_446),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1040),
.A2(n_945),
.B(n_944),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_935),
.B(n_461),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_938),
.A2(n_797),
.B(n_776),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_994),
.B(n_1039),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_938),
.A2(n_797),
.B(n_776),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1056),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1022),
.B(n_769),
.C(n_618),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_994),
.B(n_1039),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1038),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_958),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_994),
.B(n_1039),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_947),
.A2(n_797),
.B(n_776),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_994),
.B(n_1039),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1035),
.B(n_826),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_942),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_994),
.B(n_1039),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_973),
.B(n_761),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_947),
.A2(n_797),
.B(n_776),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1178)
);

BUFx4_ASAP7_75t_SL g1179 ( 
.A(n_1014),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_938),
.A2(n_954),
.B(n_937),
.Y(n_1180)
);

INVxp67_ASAP7_75t_SL g1181 ( 
.A(n_1037),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_939),
.A2(n_769),
.B(n_597),
.C(n_618),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_939),
.A2(n_769),
.B1(n_597),
.B2(n_618),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_942),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_994),
.B(n_1039),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_973),
.B(n_761),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1035),
.B(n_826),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_936),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_971),
.B(n_766),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_975),
.A2(n_974),
.B(n_972),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1156),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1188),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1144),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1077),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_1092),
.B(n_1142),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1174),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1109),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1133),
.A2(n_1155),
.B(n_1105),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1184),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_1164),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1079),
.B(n_1176),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1112),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1072),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1161),
.A2(n_1170),
.B(n_1178),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1186),
.B(n_1159),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1134),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1070),
.A2(n_1068),
.B(n_1088),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1081),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1156),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1083),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1075),
.A2(n_1090),
.B(n_1086),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_1097),
.B(n_1104),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1128),
.A2(n_1093),
.B(n_1125),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1140),
.A2(n_1122),
.B(n_1150),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1085),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1159),
.B(n_1165),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1167),
.B(n_1157),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1126),
.A2(n_1124),
.B1(n_1117),
.B2(n_1087),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1101),
.A2(n_1098),
.B(n_1107),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1165),
.B(n_1169),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1136),
.A2(n_1124),
.B(n_1096),
.C(n_1084),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1173),
.B(n_1187),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1173),
.B(n_1187),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1179),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1097),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1175),
.B(n_1185),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_1073),
.B1(n_1122),
.B2(n_1153),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1074),
.A2(n_1063),
.B(n_1110),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1167),
.A2(n_1114),
.B1(n_1082),
.B2(n_1123),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1061),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1132),
.B(n_1091),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1102),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1075),
.A2(n_1158),
.B(n_1162),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1132),
.B(n_1181),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1103),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_1173),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1080),
.A2(n_1064),
.B(n_1073),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_1180),
.B(n_1071),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1089),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1166),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1111),
.A2(n_1108),
.B(n_1119),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_SL g1245 ( 
.A(n_1131),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1118),
.B(n_1095),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1104),
.B(n_1163),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1065),
.B(n_1069),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1130),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1121),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1137),
.A2(n_1099),
.B(n_1129),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1116),
.B(n_1138),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1187),
.B(n_1115),
.Y(n_1253)
);

OAI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_1127),
.A2(n_1121),
.B1(n_1067),
.B2(n_1069),
.C(n_1076),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1152),
.B(n_1149),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1127),
.A2(n_1150),
.B(n_1060),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1106),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1060),
.A2(n_1066),
.B(n_1135),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1139),
.A2(n_1146),
.B(n_1089),
.Y(n_1259)
);

INVx8_ASAP7_75t_L g1260 ( 
.A(n_1113),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1115),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1145),
.A2(n_1148),
.B(n_1163),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1189),
.A2(n_1154),
.B(n_1147),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1094),
.A2(n_1120),
.B(n_1141),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1151),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1120),
.A2(n_1190),
.B(n_1161),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1143),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1143),
.B(n_1056),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_769),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1176),
.B(n_1186),
.Y(n_1272)
);

AOI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1100),
.A2(n_1075),
.B(n_1090),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1062),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1062),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1062),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1173),
.B(n_1187),
.Y(n_1277)
);

AOI21xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1092),
.A2(n_480),
.B(n_486),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1164),
.A2(n_1183),
.B1(n_769),
.B2(n_1022),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1144),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1062),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_SL g1283 ( 
.A1(n_1164),
.A2(n_1006),
.B(n_939),
.C(n_1182),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1164),
.B(n_769),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1176),
.B(n_1186),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1062),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1171),
.A2(n_1177),
.A3(n_1071),
.B(n_1086),
.Y(n_1287)
);

NAND2x1_ASAP7_75t_L g1288 ( 
.A(n_1081),
.B(n_1035),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1096),
.A2(n_1177),
.B(n_1171),
.Y(n_1289)
);

INVx8_ASAP7_75t_L g1290 ( 
.A(n_1173),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1112),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1096),
.A2(n_1177),
.B(n_1171),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1171),
.A2(n_1177),
.B(n_1078),
.Y(n_1294)
);

OAI211xp5_ASAP7_75t_L g1295 ( 
.A1(n_1183),
.A2(n_1164),
.B(n_769),
.C(n_1182),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1164),
.A2(n_1183),
.B1(n_769),
.B2(n_1022),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1164),
.A2(n_1006),
.B(n_939),
.C(n_1182),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1062),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1142),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1164),
.A2(n_1006),
.B(n_939),
.C(n_1182),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1183),
.A2(n_769),
.B1(n_597),
.B2(n_893),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1079),
.B(n_1176),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_SL g1304 ( 
.A1(n_1164),
.A2(n_1006),
.B(n_939),
.C(n_1182),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1171),
.A2(n_1177),
.B(n_1078),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1168),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1062),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1234),
.B(n_1217),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1192),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1211),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1280),
.A2(n_1297),
.B1(n_1284),
.B2(n_1219),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1234),
.B(n_1221),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1222),
.A2(n_1229),
.B(n_1223),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1211),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1237),
.B(n_1206),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1191),
.B(n_1210),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1216),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1237),
.B(n_1284),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1271),
.A2(n_1201),
.B(n_1295),
.C(n_1283),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1283),
.A2(n_1304),
.B(n_1301),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1298),
.A2(n_1304),
.B(n_1301),
.C(n_1297),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1249),
.B(n_1250),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1280),
.A2(n_1239),
.B1(n_1300),
.B2(n_1277),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1250),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1232),
.B(n_1246),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1287),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1192),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1191),
.B(n_1210),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1198),
.A2(n_1224),
.B1(n_1303),
.B2(n_1202),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1204),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1195),
.Y(n_1332)
);

O2A1O1Ixp5_ASAP7_75t_L g1333 ( 
.A1(n_1212),
.A2(n_1264),
.B(n_1273),
.C(n_1248),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1272),
.B(n_1285),
.Y(n_1334)
);

OAI31xp33_ASAP7_75t_L g1335 ( 
.A1(n_1254),
.A2(n_1225),
.A3(n_1226),
.B(n_1218),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1195),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1235),
.B(n_1227),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1294),
.A2(n_1305),
.B(n_1257),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1275),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1277),
.A2(n_1230),
.B1(n_1203),
.B2(n_1291),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1209),
.B(n_1252),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1275),
.B(n_1276),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1240),
.B(n_1230),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_L g1344 ( 
.A1(n_1248),
.A2(n_1236),
.B(n_1288),
.C(n_1253),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1209),
.B(n_1255),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1278),
.A2(n_1197),
.B1(n_1281),
.B2(n_1193),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1197),
.A2(n_1233),
.B1(n_1243),
.B2(n_1290),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1290),
.A2(n_1207),
.B1(n_1265),
.B2(n_1199),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1276),
.B(n_1307),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1244),
.A2(n_1256),
.B(n_1251),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1245),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1282),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1282),
.B(n_1307),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1207),
.B(n_1286),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1290),
.A2(n_1194),
.B1(n_1196),
.B2(n_1299),
.Y(n_1355)
);

NAND4xp25_ASAP7_75t_L g1356 ( 
.A(n_1274),
.B(n_1286),
.C(n_1213),
.D(n_1261),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1300),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1287),
.B(n_1240),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_SL g1359 ( 
.A1(n_1215),
.A2(n_1268),
.B(n_1263),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1260),
.B(n_1247),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1228),
.A2(n_1260),
.B1(n_1240),
.B2(n_1242),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1228),
.A2(n_1260),
.B1(n_1242),
.B2(n_1241),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1262),
.B(n_1259),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1267),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1287),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1289),
.B(n_1293),
.Y(n_1367)
);

CKINVDCx12_ASAP7_75t_R g1368 ( 
.A(n_1238),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1262),
.B(n_1259),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1238),
.A2(n_1258),
.B1(n_1266),
.B2(n_1231),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1214),
.Y(n_1371)
);

BUFx2_ASAP7_75t_R g1372 ( 
.A(n_1208),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1200),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1205),
.B(n_1269),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1205),
.A2(n_1269),
.B(n_1270),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1270),
.A2(n_1279),
.B(n_1292),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_1306),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1296),
.B(n_1306),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1284),
.A2(n_1164),
.B1(n_1302),
.B2(n_1280),
.C(n_1297),
.Y(n_1380)
);

INVx3_ASAP7_75t_SL g1381 ( 
.A(n_1245),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1280),
.A2(n_1297),
.B1(n_1183),
.B2(n_769),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_L g1383 ( 
.A1(n_1302),
.A2(n_1295),
.B(n_1271),
.C(n_1201),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1234),
.B(n_1217),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1211),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1272),
.B(n_1285),
.Y(n_1386)
);

O2A1O1Ixp5_ASAP7_75t_L g1387 ( 
.A1(n_1302),
.A2(n_1295),
.B(n_1271),
.C(n_1201),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1302),
.A2(n_1182),
.B(n_1284),
.C(n_1224),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1191),
.B(n_1210),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1280),
.A2(n_1297),
.B1(n_1183),
.B2(n_769),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1338),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1369),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1363),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_SL g1394 ( 
.A(n_1332),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1343),
.B(n_1358),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1364),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1319),
.B(n_1316),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1317),
.B(n_1329),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1366),
.B(n_1327),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1363),
.B(n_1369),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1369),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1343),
.B(n_1365),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1367),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1317),
.B(n_1329),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1315),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1318),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1354),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1389),
.B(n_1325),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1385),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1389),
.B(n_1350),
.Y(n_1411)
);

XNOR2xp5_ASAP7_75t_L g1412 ( 
.A(n_1311),
.B(n_1382),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1371),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1370),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1373),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1349),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1371),
.B(n_1375),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1378),
.B(n_1379),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1374),
.Y(n_1422)
);

INVxp67_ASAP7_75t_R g1423 ( 
.A(n_1362),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_1324),
.B1(n_1321),
.B2(n_1326),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1339),
.B(n_1341),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1377),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1352),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1377),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1314),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1333),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1388),
.B(n_1314),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1376),
.A2(n_1320),
.B(n_1361),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1340),
.B(n_1313),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1353),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1312),
.B(n_1384),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1355),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1342),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1415),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1420),
.B(n_1411),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1415),
.Y(n_1440)
);

CKINVDCx6p67_ASAP7_75t_R g1441 ( 
.A(n_1416),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1416),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1399),
.B(n_1309),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1434),
.B(n_1322),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1426),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1434),
.B(n_1418),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1399),
.B(n_1328),
.Y(n_1447)
);

OAI222xp33_ASAP7_75t_L g1448 ( 
.A1(n_1412),
.A2(n_1383),
.B1(n_1387),
.B2(n_1347),
.C1(n_1348),
.C2(n_1323),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1395),
.B(n_1404),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1334),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1395),
.B(n_1345),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1395),
.B(n_1386),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1404),
.B(n_1356),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1396),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1404),
.B(n_1372),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1433),
.B(n_1359),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1403),
.B(n_1344),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1392),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1426),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1403),
.B(n_1335),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1428),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1421),
.B(n_1346),
.C(n_1360),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1393),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1419),
.B(n_1381),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1393),
.B(n_1337),
.Y(n_1465)
);

NOR4xp25_ASAP7_75t_SL g1466 ( 
.A(n_1391),
.B(n_1332),
.C(n_1336),
.D(n_1351),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1419),
.B(n_1381),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1405),
.B(n_1351),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1428),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1392),
.B(n_1336),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1413),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1445),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1462),
.B(n_1398),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1449),
.B(n_1409),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1392),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1462),
.A2(n_1421),
.B1(n_1412),
.B2(n_1441),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1439),
.B(n_1392),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1442),
.B(n_1412),
.C(n_1424),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1448),
.A2(n_1433),
.B(n_1424),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1442),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1471),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1458),
.B(n_1392),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1448),
.A2(n_1398),
.B1(n_1435),
.B2(n_1414),
.C(n_1391),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1460),
.A2(n_1431),
.B1(n_1433),
.B2(n_1435),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1444),
.B(n_1414),
.C(n_1436),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1450),
.B(n_1408),
.Y(n_1486)
);

NOR4xp25_ASAP7_75t_SL g1487 ( 
.A(n_1463),
.B(n_1413),
.C(n_1422),
.D(n_1423),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1441),
.A2(n_1431),
.B1(n_1436),
.B2(n_1432),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1439),
.B(n_1401),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1443),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1460),
.A2(n_1456),
.B1(n_1431),
.B2(n_1432),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1465),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1453),
.Y(n_1493)
);

OAI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1460),
.A2(n_1444),
.B(n_1457),
.C(n_1453),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1468),
.A2(n_1429),
.B1(n_1409),
.B2(n_1408),
.C(n_1402),
.Y(n_1495)
);

OAI211xp5_ASAP7_75t_L g1496 ( 
.A1(n_1457),
.A2(n_1357),
.B(n_1430),
.C(n_1410),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1441),
.A2(n_1423),
.B1(n_1429),
.B2(n_1430),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1466),
.A2(n_1394),
.B1(n_1429),
.B2(n_1430),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1468),
.A2(n_1394),
.B1(n_1406),
.B2(n_1407),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1454),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1443),
.A2(n_1407),
.B1(n_1406),
.B2(n_1410),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1454),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1453),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1450),
.B(n_1425),
.Y(n_1505)
);

AOI222xp33_ASAP7_75t_L g1506 ( 
.A1(n_1457),
.A2(n_1357),
.B1(n_1425),
.B2(n_1427),
.C1(n_1437),
.C2(n_1397),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1447),
.A2(n_1427),
.B1(n_1400),
.B2(n_1417),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1446),
.A2(n_1402),
.B1(n_1393),
.B2(n_1437),
.C(n_1400),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1459),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1509),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1450),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1501),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1504),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1449),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1491),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1478),
.B(n_1440),
.C(n_1438),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1501),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1472),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1470),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1503),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1485),
.B(n_1465),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1481),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1492),
.B(n_1479),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1492),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1488),
.A2(n_1461),
.B(n_1469),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1496),
.Y(n_1528)
);

NOR2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1470),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1526),
.B(n_1492),
.Y(n_1530)
);

AND2x4_ASAP7_75t_SL g1531 ( 
.A(n_1525),
.B(n_1464),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1513),
.B(n_1494),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1519),
.B(n_1368),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1513),
.B(n_1505),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1525),
.Y(n_1535)
);

AOI211x1_ASAP7_75t_L g1536 ( 
.A1(n_1516),
.A2(n_1495),
.B(n_1508),
.C(n_1498),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1519),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1522),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1529),
.A2(n_1476),
.B1(n_1432),
.B2(n_1500),
.Y(n_1545)
);

NOR2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1516),
.B(n_1470),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1510),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_SL g1552 ( 
.A(n_1521),
.B(n_1499),
.C(n_1507),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1486),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1521),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1515),
.B(n_1502),
.C(n_1467),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1526),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1452),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1518),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1524),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1526),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1475),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1528),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

OAI21xp33_ASAP7_75t_L g1568 ( 
.A1(n_1524),
.A2(n_1506),
.B(n_1455),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1567),
.B(n_1477),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1532),
.B(n_1517),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1560),
.B(n_1544),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1541),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1567),
.B(n_1489),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1532),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1547),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1548),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1447),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1559),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1536),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1452),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1553),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1557),
.B(n_1464),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1565),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1531),
.B(n_1527),
.Y(n_1587)
);

AOI32xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1552),
.A2(n_1533),
.A3(n_1553),
.B1(n_1555),
.B2(n_1546),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1562),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1464),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1566),
.B(n_1520),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1545),
.A2(n_1487),
.B(n_1527),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1554),
.B(n_1451),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1535),
.B(n_1527),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1547),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1535),
.B(n_1527),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1520),
.Y(n_1598)
);

OAI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1545),
.A2(n_1527),
.B1(n_1528),
.B2(n_1455),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1546),
.B(n_1467),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1550),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1550),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1535),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1579),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1572),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1572),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1592),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1539),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1581),
.A2(n_1528),
.B1(n_1568),
.B2(n_1558),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1577),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1592),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1595),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1595),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1589),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1583),
.B(n_1368),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1588),
.A2(n_1534),
.B1(n_1455),
.B2(n_1540),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1598),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1597),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1590),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1623),
.A2(n_1599),
.B(n_1571),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1606),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1606),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1611),
.B(n_1598),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1623),
.A2(n_1599),
.B1(n_1573),
.B2(n_1593),
.Y(n_1633)
);

NAND2x1_ASAP7_75t_L g1634 ( 
.A(n_1621),
.B(n_1563),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1622),
.A2(n_1573),
.B1(n_1598),
.B2(n_1528),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1614),
.Y(n_1636)
);

INVxp33_ASAP7_75t_L g1637 ( 
.A(n_1611),
.Y(n_1637)
);

OAI322xp33_ASAP7_75t_L g1638 ( 
.A1(n_1607),
.A2(n_1570),
.A3(n_1585),
.B1(n_1602),
.B2(n_1596),
.C1(n_1601),
.C2(n_1580),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1608),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1578),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1610),
.B(n_1624),
.Y(n_1641)
);

NAND2x1_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1563),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1627),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1575),
.Y(n_1645)
);

OAI32xp33_ASAP7_75t_L g1646 ( 
.A1(n_1612),
.A2(n_1563),
.A3(n_1587),
.B1(n_1597),
.B2(n_1538),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1647)
);

CKINVDCx16_ASAP7_75t_R g1648 ( 
.A(n_1639),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1637),
.B(n_1616),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1639),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1608),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1632),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1633),
.A2(n_1604),
.B1(n_1609),
.B2(n_1616),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1636),
.B(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1628),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1630),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1657),
.B(n_1629),
.C(n_1635),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1648),
.B(n_1643),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1655),
.A2(n_1646),
.B(n_1642),
.C(n_1634),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1647),
.A2(n_1604),
.B1(n_1609),
.B2(n_1625),
.Y(n_1662)
);

AOI322xp5_ASAP7_75t_L g1663 ( 
.A1(n_1649),
.A2(n_1631),
.A3(n_1609),
.B1(n_1605),
.B2(n_1603),
.C1(n_1613),
.C2(n_1620),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1651),
.A2(n_1638),
.B(n_1625),
.C(n_1614),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1653),
.A2(n_1645),
.B(n_1603),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1647),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1667),
.Y(n_1668)
);

OAI322xp33_ASAP7_75t_L g1669 ( 
.A1(n_1660),
.A2(n_1653),
.A3(n_1666),
.B1(n_1654),
.B2(n_1662),
.C1(n_1665),
.C2(n_1658),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1664),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1656),
.B1(n_1650),
.B2(n_1652),
.C(n_1645),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_SL g1672 ( 
.A1(n_1661),
.A2(n_1658),
.B(n_1603),
.C(n_1605),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1668),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1672),
.B(n_1652),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1671),
.B(n_1605),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1669),
.Y(n_1676)
);

XOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1670),
.B(n_1604),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1672),
.A2(n_1663),
.B(n_1604),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1673),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1675),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1678),
.A2(n_1618),
.B(n_1613),
.C(n_1620),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1677),
.Y(n_1682)
);

XOR2xp5_ASAP7_75t_L g1683 ( 
.A(n_1676),
.B(n_1604),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_L g1684 ( 
.A(n_1683),
.B(n_1674),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1681),
.A2(n_1618),
.B(n_1619),
.C(n_1621),
.Y(n_1685)
);

OAI22x1_ASAP7_75t_L g1686 ( 
.A1(n_1679),
.A2(n_1621),
.B1(n_1619),
.B2(n_1615),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1684),
.B(n_1682),
.Y(n_1687)
);

AOI322xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1680),
.A3(n_1617),
.B1(n_1626),
.B2(n_1615),
.C1(n_1685),
.C2(n_1686),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1626),
.B1(n_1617),
.B2(n_1615),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1617),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1690),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1626),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1691),
.B(n_1575),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1587),
.B(n_1591),
.Y(n_1694)
);

XOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1692),
.B(n_1594),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1538),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1694),
.A2(n_1530),
.B1(n_1549),
.B2(n_1558),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1696),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1697),
.B1(n_1561),
.B2(n_1551),
.Y(n_1699)
);

AOI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1561),
.B(n_1551),
.C(n_1530),
.Y(n_1700)
);


endmodule