module fake_netlist_5_2362_n_1023 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1023);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1023;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_568;
wire n_509;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_969;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_795;
wire n_710;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_40),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_166),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_16),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_47),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_159),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_37),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_187),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_181),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_32),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_42),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_88),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_137),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_162),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_60),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_173),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_126),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_160),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_149),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_101),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_62),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_193),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_124),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_213),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_24),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_130),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_123),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_17),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_157),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_96),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_139),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_104),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_36),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_84),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_85),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_117),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_146),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_150),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_76),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_103),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_31),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_54),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_17),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_48),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_64),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_121),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_20),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_111),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_90),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_28),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_114),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_86),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_113),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_30),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_275),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_218),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_221),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_226),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_231),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_234),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_236),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_223),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_240),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_239),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_0),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_219),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_224),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_225),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_233),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_243),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_244),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_230),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_238),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_1),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_235),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_253),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_245),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_249),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_220),
.B(n_259),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_242),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_247),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_262),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_246),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_250),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_263),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_268),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_268),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_273),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_274),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_265),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_310),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_361),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_344),
.B(n_302),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_312),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_330),
.B(n_273),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_320),
.A2(n_282),
.B(n_277),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_288),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_302),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_349),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_308),
.B(n_222),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_290),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_315),
.B(n_292),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_317),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_294),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_362),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_321),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_345),
.B(n_301),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_318),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_325),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_318),
.B(n_254),
.Y(n_423)
);

OR2x6_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_248),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_405),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_252),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_269),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_305),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_415),
.A2(n_295),
.B1(n_279),
.B2(n_271),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_365),
.B(n_279),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_385),
.B(n_255),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_413),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_295),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_385),
.B(n_389),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_385),
.B(n_257),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_366),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_289),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_293),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_385),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_410),
.B(n_258),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_410),
.B(n_411),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_365),
.B(n_260),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_410),
.B(n_261),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_264),
.Y(n_466)
);

INVx3_ASAP7_75t_R g467 ( 
.A(n_409),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_373),
.B(n_382),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_392),
.B(n_272),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_407),
.B(n_296),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_276),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_412),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_418),
.B(n_278),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_410),
.B(n_281),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_418),
.B(n_222),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_411),
.B(n_297),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_406),
.B(n_283),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_422),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_227),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_411),
.B(n_284),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_366),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_299),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_374),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_227),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_374),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

BUFx6f_ASAP7_75t_SL g497 ( 
.A(n_419),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_375),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_411),
.B(n_300),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_454),
.B(n_406),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_454),
.B(n_406),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_420),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_397),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_397),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_461),
.A2(n_372),
.B1(n_383),
.B2(n_414),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_445),
.B(n_387),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_461),
.B(n_397),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_372),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_383),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_444),
.A2(n_367),
.B1(n_414),
.B2(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_464),
.B(n_367),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_476),
.B(n_408),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_464),
.B(n_388),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

AO22x1_ASAP7_75t_L g520 ( 
.A1(n_435),
.A2(n_307),
.B1(n_409),
.B2(n_306),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_494),
.C(n_449),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_432),
.B(n_401),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_428),
.B(n_388),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_437),
.B(n_377),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_436),
.B(n_388),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_401),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_430),
.B(n_402),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_460),
.B(n_450),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_500),
.B(n_390),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_328),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_SL g532 ( 
.A(n_438),
.B(n_306),
.C(n_287),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_460),
.B(n_375),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_466),
.A2(n_390),
.B(n_375),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_457),
.B(n_480),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_500),
.A2(n_402),
.B1(n_399),
.B2(n_370),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

NAND2x1_ASAP7_75t_L g540 ( 
.A(n_431),
.B(n_453),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_475),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_328),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_448),
.B(n_402),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_494),
.B(n_285),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_434),
.B(n_304),
.C(n_291),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_444),
.A2(n_371),
.B(n_379),
.C(n_369),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_475),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_493),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_499),
.B(n_375),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_379),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_473),
.A2(n_363),
.B1(n_334),
.B2(n_347),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_486),
.B(n_379),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_458),
.B(n_364),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_331),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_463),
.B(n_364),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_478),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_473),
.B(n_422),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_433),
.A2(n_376),
.B1(n_369),
.B2(n_364),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_433),
.A2(n_376),
.B1(n_384),
.B2(n_355),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_479),
.B(n_331),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_438),
.B(n_462),
.Y(n_564)
);

AND2x6_ASAP7_75t_L g565 ( 
.A(n_462),
.B(n_384),
.Y(n_565)
);

NOR2x2_ASAP7_75t_L g566 ( 
.A(n_424),
.B(n_334),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_487),
.B(n_347),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_459),
.B(n_1),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_453),
.B(n_384),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_459),
.B(n_348),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_424),
.B(n_348),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_465),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_483),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_482),
.B(n_355),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_483),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_465),
.Y(n_578)
);

AND2x6_ASAP7_75t_SL g579 ( 
.A(n_490),
.B(n_421),
.Y(n_579)
);

CKINVDCx11_ASAP7_75t_R g580 ( 
.A(n_479),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_483),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_482),
.B(n_477),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_505),
.B(n_474),
.Y(n_584)
);

CKINVDCx11_ASAP7_75t_R g585 ( 
.A(n_579),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_569),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_512),
.B(n_467),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_SL g589 ( 
.A(n_564),
.B(n_497),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_528),
.B(n_474),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_528),
.B(n_489),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_515),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_577),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_568),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_558),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_525),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_569),
.Y(n_597)
);

AND2x6_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_492),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_536),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_543),
.B(n_489),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_L g603 ( 
.A(n_521),
.B(n_472),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_512),
.B(n_497),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_577),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_542),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_492),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_560),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_541),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_565),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_580),
.B(n_360),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_511),
.B(n_360),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_574),
.B(n_456),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_519),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_535),
.B(n_495),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_543),
.B(n_433),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_522),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_SL g624 ( 
.A(n_555),
.B(n_363),
.C(n_471),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_537),
.B(n_433),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_511),
.B(n_496),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_574),
.B(n_433),
.Y(n_628)
);

O2A1O1Ixp5_ASAP7_75t_L g629 ( 
.A1(n_523),
.A2(n_481),
.B(n_495),
.C(n_441),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_562),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_522),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_578),
.B(n_439),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_508),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_578),
.B(n_506),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_527),
.B(n_439),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_550),
.B(n_441),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_516),
.B(n_456),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_581),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_565),
.B(n_456),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_570),
.B(n_440),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_526),
.B(n_452),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_518),
.B(n_529),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_539),
.B(n_452),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_565),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_527),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_552),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_544),
.B(n_440),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_549),
.B(n_440),
.Y(n_649)
);

NAND2x1p5_ASAP7_75t_L g650 ( 
.A(n_646),
.B(n_559),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_517),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_624),
.B(n_531),
.C(n_513),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_640),
.A2(n_504),
.B(n_501),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_584),
.A2(n_533),
.B(n_547),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_590),
.A2(n_534),
.B(n_538),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_646),
.B(n_509),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_607),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_627),
.B(n_507),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_629),
.A2(n_530),
.B(n_582),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_591),
.A2(n_546),
.B(n_545),
.C(n_510),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_646),
.B(n_576),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_643),
.A2(n_456),
.B(n_530),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_602),
.A2(n_583),
.A3(n_554),
.B(n_556),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_627),
.B(n_588),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_613),
.A2(n_538),
.B1(n_561),
.B2(n_562),
.Y(n_665)
);

OAI21x1_ASAP7_75t_SL g666 ( 
.A1(n_645),
.A2(n_561),
.B(n_553),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_613),
.A2(n_551),
.B(n_571),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_595),
.B(n_563),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_596),
.B(n_572),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_622),
.A2(n_557),
.B(n_560),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_609),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_629),
.A2(n_540),
.B(n_532),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_646),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_599),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_618),
.B(n_573),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_641),
.A2(n_447),
.B1(n_483),
.B2(n_498),
.Y(n_676)
);

AO21x2_ASAP7_75t_L g677 ( 
.A1(n_625),
.A2(n_532),
.B(n_520),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_447),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g679 ( 
.A1(n_614),
.A2(n_566),
.B(n_447),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_637),
.A2(n_498),
.B(n_496),
.Y(n_680)
);

AO31x2_ASAP7_75t_L g681 ( 
.A1(n_642),
.A2(n_447),
.A3(n_3),
.B(n_4),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_638),
.A2(n_39),
.B(n_38),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_638),
.A2(n_44),
.B(n_43),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_616),
.A2(n_46),
.B(n_45),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_628),
.A2(n_633),
.A3(n_644),
.B(n_588),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_608),
.B(n_50),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_594),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_648),
.A2(n_53),
.B(n_51),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_619),
.A2(n_56),
.B(n_55),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_604),
.B(n_2),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_604),
.B(n_3),
.Y(n_691)
);

OAI21x1_ASAP7_75t_SL g692 ( 
.A1(n_645),
.A2(n_58),
.B(n_57),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_4),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_620),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_641),
.A2(n_589),
.B(n_624),
.C(n_632),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_598),
.B(n_5),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_619),
.A2(n_109),
.B(n_216),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_586),
.B(n_6),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_649),
.A2(n_110),
.B(n_215),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_616),
.A2(n_108),
.B1(n_214),
.B2(n_212),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_587),
.A2(n_106),
.B(n_211),
.Y(n_703)
);

AO31x2_ASAP7_75t_L g704 ( 
.A1(n_601),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_616),
.A2(n_105),
.B1(n_210),
.B2(n_207),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_655),
.A2(n_616),
.B(n_606),
.Y(n_706)
);

NAND2x1p5_ASAP7_75t_L g707 ( 
.A(n_673),
.B(n_593),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_652),
.A2(n_598),
.B1(n_603),
.B2(n_589),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_680),
.A2(n_639),
.B(n_600),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_658),
.A2(n_598),
.B(n_611),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_668),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_651),
.B(n_623),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_696),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_659),
.A2(n_639),
.B(n_600),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_653),
.A2(n_597),
.B(n_587),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_672),
.A2(n_597),
.B(n_592),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_652),
.A2(n_598),
.B1(n_611),
.B2(n_621),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_673),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_SL g720 ( 
.A1(n_697),
.A2(n_586),
.B(n_605),
.C(n_631),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_662),
.A2(n_606),
.B(n_593),
.Y(n_721)
);

OA21x2_ASAP7_75t_L g722 ( 
.A1(n_654),
.A2(n_630),
.B(n_615),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_694),
.B(n_636),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_695),
.A2(n_605),
.B1(n_647),
.B2(n_631),
.Y(n_724)
);

AO21x2_ASAP7_75t_L g725 ( 
.A1(n_666),
.A2(n_621),
.B(n_636),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_664),
.B(n_598),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_656),
.B(n_610),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_660),
.A2(n_626),
.B(n_610),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_626),
.B(n_617),
.C(n_585),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_671),
.B(n_675),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_703),
.A2(n_612),
.B(n_599),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_682),
.A2(n_612),
.B(n_599),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_665),
.A2(n_612),
.B1(n_599),
.B2(n_617),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_693),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_691),
.A2(n_585),
.B1(n_612),
.B2(n_9),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_698),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_663),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

BUFx2_ASAP7_75t_R g740 ( 
.A(n_677),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_704),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_704),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_667),
.A2(n_107),
.B(n_205),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_668),
.B(n_674),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

AO21x2_ASAP7_75t_L g746 ( 
.A1(n_670),
.A2(n_102),
.B(n_203),
.Y(n_746)
);

AO31x2_ASAP7_75t_L g747 ( 
.A1(n_676),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_668),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_704),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_687),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_663),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_677),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_669),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_688),
.A2(n_118),
.B(n_202),
.Y(n_754)
);

AOI21xp33_ASAP7_75t_L g755 ( 
.A1(n_661),
.A2(n_16),
.B(n_18),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_701),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_683),
.A2(n_119),
.B(n_201),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_750),
.B(n_687),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_736),
.Y(n_759)
);

AOI21x1_ASAP7_75t_L g760 ( 
.A1(n_721),
.A2(n_686),
.B(n_689),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_730),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_741),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_723),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_744),
.B(n_650),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_744),
.B(n_679),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_750),
.B(n_679),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_708),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_744),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_714),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_R g770 ( 
.A(n_723),
.B(n_700),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_713),
.B(n_724),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_719),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_692),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_739),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_719),
.B(n_684),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_SL g776 ( 
.A(n_735),
.B(n_699),
.C(n_702),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_735),
.B(n_681),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_757),
.A2(n_705),
.B1(n_685),
.B2(n_681),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_748),
.B(n_685),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_742),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_745),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_724),
.A2(n_685),
.B1(n_663),
.B2(n_21),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_734),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_712),
.B(n_19),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_711),
.A2(n_19),
.B(n_20),
.Y(n_785)
);

INVx8_ASAP7_75t_L g786 ( 
.A(n_745),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_709),
.B(n_22),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_745),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_706),
.A2(n_217),
.B(n_122),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_745),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_726),
.B(n_59),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_709),
.B(n_23),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_737),
.B(n_23),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_R g795 ( 
.A(n_727),
.B(n_61),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_707),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_749),
.Y(n_797)
);

NOR2x1_ASAP7_75t_L g798 ( 
.A(n_728),
.B(n_24),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_746),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_SL g801 ( 
.A1(n_752),
.A2(n_28),
.B(n_29),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_737),
.B(n_29),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_729),
.B(n_30),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_755),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_804)
);

OAI221xp5_ASAP7_75t_L g805 ( 
.A1(n_753),
.A2(n_34),
.B1(n_35),
.B2(n_63),
.C(n_65),
.Y(n_805)
);

OAI211xp5_ASAP7_75t_SL g806 ( 
.A1(n_752),
.A2(n_35),
.B(n_66),
.C(n_67),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_718),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_807)
);

OAI211xp5_ASAP7_75t_SL g808 ( 
.A1(n_720),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_808)
);

AOI211xp5_ASAP7_75t_L g809 ( 
.A1(n_720),
.A2(n_75),
.B(n_77),
.C(n_78),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_738),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_200),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_740),
.B(n_79),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_746),
.A2(n_725),
.B1(n_722),
.B2(n_743),
.Y(n_813)
);

OAI211xp5_ASAP7_75t_SL g814 ( 
.A1(n_803),
.A2(n_738),
.B(n_751),
.C(n_747),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_SL g815 ( 
.A1(n_785),
.A2(n_732),
.B(n_754),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_782),
.A2(n_717),
.B(n_776),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_762),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_794),
.A2(n_725),
.B1(n_722),
.B2(n_751),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_802),
.A2(n_805),
.B1(n_801),
.B2(n_812),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_707),
.B1(n_756),
.B2(n_747),
.Y(n_820)
);

OAI221xp5_ASAP7_75t_SL g821 ( 
.A1(n_804),
.A2(n_747),
.B1(n_754),
.B2(n_82),
.C(n_83),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_806),
.A2(n_756),
.B1(n_716),
.B2(n_731),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_787),
.A2(n_756),
.B1(n_716),
.B2(n_731),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_766),
.A2(n_756),
.B1(n_747),
.B2(n_732),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_777),
.A2(n_710),
.B1(n_715),
.B2(n_717),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_801),
.A2(n_715),
.B1(n_81),
.B2(n_89),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_780),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_792),
.A2(n_80),
.B1(n_91),
.B2(n_93),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_761),
.B(n_94),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_761),
.B(n_771),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_780),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_769),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_798),
.A2(n_198),
.B1(n_97),
.B2(n_98),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_798),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_797),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_SL g837 ( 
.A1(n_807),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_759),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_799),
.A2(n_770),
.B1(n_765),
.B2(n_811),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_784),
.B(n_125),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_800),
.A2(n_127),
.B1(n_128),
.B2(n_131),
.Y(n_841)
);

AOI21xp33_ASAP7_75t_L g842 ( 
.A1(n_778),
.A2(n_809),
.B(n_773),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_132),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_765),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_808),
.A2(n_196),
.B1(n_141),
.B2(n_142),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_789),
.B(n_138),
.C(n_143),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_779),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_758),
.A2(n_764),
.B1(n_763),
.B2(n_773),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_781),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_797),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_813),
.A2(n_775),
.B(n_793),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_810),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_791),
.A2(n_144),
.B1(n_145),
.B2(n_148),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_791),
.A2(n_763),
.B1(n_768),
.B2(n_764),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_796),
.A2(n_152),
.B(n_154),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_772),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_760),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.C(n_163),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_791),
.A2(n_195),
.B1(n_168),
.B2(n_169),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_817),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_828),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_832),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_836),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_831),
.B(n_850),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_852),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_856),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_825),
.B(n_791),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_816),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_818),
.B(n_826),
.Y(n_869)
);

NOR2x1_ASAP7_75t_L g870 ( 
.A(n_814),
.B(n_774),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_816),
.B(n_772),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_838),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_822),
.B(n_833),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_843),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_851),
.B(n_788),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_849),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_819),
.B(n_793),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_815),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_824),
.B(n_793),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_788),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_848),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_821),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_854),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_830),
.B(n_788),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_857),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_846),
.Y(n_888)
);

OA21x2_ASAP7_75t_L g889 ( 
.A1(n_827),
.A2(n_164),
.B(n_171),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_840),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_854),
.B(n_781),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_844),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_884),
.A2(n_839),
.B1(n_842),
.B2(n_845),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_875),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_862),
.Y(n_895)
);

OAI221xp5_ASAP7_75t_L g896 ( 
.A1(n_884),
.A2(n_841),
.B1(n_858),
.B2(n_853),
.C(n_835),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_862),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_872),
.Y(n_898)
);

OAI211xp5_ASAP7_75t_L g899 ( 
.A1(n_880),
.A2(n_845),
.B(n_841),
.C(n_834),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_869),
.B(n_827),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_887),
.A2(n_858),
.B1(n_853),
.B2(n_834),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_863),
.Y(n_902)
);

NOR4xp25_ASAP7_75t_SL g903 ( 
.A(n_876),
.B(n_855),
.C(n_835),
.D(n_829),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_865),
.Y(n_904)
);

NAND4xp25_ASAP7_75t_L g905 ( 
.A(n_876),
.B(n_837),
.C(n_774),
.D(n_790),
.Y(n_905)
);

AO21x2_ASAP7_75t_L g906 ( 
.A1(n_868),
.A2(n_880),
.B(n_871),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_875),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_863),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_865),
.Y(n_909)
);

OAI211xp5_ASAP7_75t_SL g910 ( 
.A1(n_872),
.A2(n_790),
.B(n_786),
.C(n_781),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_887),
.A2(n_786),
.B1(n_174),
.B2(n_175),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_861),
.Y(n_912)
);

OAI211xp5_ASAP7_75t_SL g913 ( 
.A1(n_879),
.A2(n_172),
.B(n_177),
.C(n_179),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_859),
.B(n_180),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_906),
.B(n_859),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_912),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_895),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_894),
.B(n_871),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_904),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_894),
.B(n_871),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_907),
.B(n_875),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_907),
.B(n_869),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_906),
.B(n_869),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_904),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_906),
.B(n_868),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_909),
.B(n_885),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_909),
.B(n_885),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_921),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_916),
.B(n_898),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_917),
.Y(n_931)
);

AND2x4_ASAP7_75t_SL g932 ( 
.A(n_921),
.B(n_875),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_925),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_919),
.Y(n_934)
);

AND2x4_ASAP7_75t_SL g935 ( 
.A(n_921),
.B(n_891),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_922),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_927),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_919),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_936),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_936),
.B(n_899),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_931),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_933),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_934),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_932),
.B(n_929),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_932),
.B(n_923),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_930),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_SL g947 ( 
.A(n_930),
.B(n_903),
.C(n_893),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_SL g948 ( 
.A1(n_946),
.A2(n_901),
.B1(n_896),
.B2(n_900),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_947),
.B(n_885),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_940),
.A2(n_900),
.B1(n_923),
.B2(n_867),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_941),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_948),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_949),
.B(n_940),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_950),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_954),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_952),
.B(n_951),
.Y(n_956)
);

XOR2x2_ASAP7_75t_L g957 ( 
.A(n_953),
.B(n_939),
.Y(n_957)
);

AOI21xp33_ASAP7_75t_L g958 ( 
.A1(n_952),
.A2(n_940),
.B(n_942),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_940),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_L g960 ( 
.A(n_958),
.B(n_913),
.C(n_911),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_943),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_945),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_955),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_955),
.B(n_945),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_958),
.B(n_889),
.C(n_914),
.Y(n_965)
);

XNOR2x1_ASAP7_75t_L g966 ( 
.A(n_957),
.B(n_914),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_SL g967 ( 
.A1(n_966),
.A2(n_962),
.B(n_959),
.Y(n_967)
);

OAI211xp5_ASAP7_75t_L g968 ( 
.A1(n_963),
.A2(n_889),
.B(n_888),
.C(n_944),
.Y(n_968)
);

OAI211xp5_ASAP7_75t_SL g969 ( 
.A1(n_964),
.A2(n_887),
.B(n_879),
.C(n_915),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_961),
.B(n_944),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_965),
.A2(n_905),
.B(n_910),
.Y(n_971)
);

NOR3x1_ASAP7_75t_L g972 ( 
.A(n_960),
.B(n_915),
.C(n_890),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_963),
.B(n_922),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_973),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_970),
.Y(n_975)
);

NAND4xp25_ASAP7_75t_L g976 ( 
.A(n_967),
.B(n_972),
.C(n_968),
.D(n_971),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_969),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_970),
.Y(n_978)
);

NAND4xp75_ASAP7_75t_L g979 ( 
.A(n_972),
.B(n_926),
.C(n_889),
.D(n_870),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_937),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_SL g981 ( 
.A1(n_970),
.A2(n_926),
.B(n_938),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_978),
.A2(n_935),
.B1(n_888),
.B2(n_885),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_975),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_976),
.A2(n_888),
.B(n_889),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_980),
.B(n_182),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_977),
.B(n_890),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_928),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_981),
.B(n_885),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_978),
.A2(n_889),
.B(n_867),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_975),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_978),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_992),
.Y(n_993)
);

AOI211xp5_ASAP7_75t_L g994 ( 
.A1(n_991),
.A2(n_928),
.B(n_927),
.C(n_886),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_982),
.A2(n_920),
.B1(n_918),
.B2(n_890),
.Y(n_995)
);

INVxp67_ASAP7_75t_SL g996 ( 
.A(n_983),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_984),
.A2(n_875),
.B1(n_883),
.B2(n_892),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_987),
.A2(n_883),
.B1(n_892),
.B2(n_891),
.Y(n_998)
);

OAI221xp5_ASAP7_75t_L g999 ( 
.A1(n_989),
.A2(n_886),
.B1(n_874),
.B2(n_892),
.C(n_881),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_985),
.B(n_920),
.Y(n_1000)
);

NOR4xp25_ASAP7_75t_L g1001 ( 
.A(n_988),
.B(n_918),
.C(n_902),
.D(n_908),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_990),
.A2(n_883),
.B1(n_891),
.B2(n_874),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_993),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_1000),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_1001),
.B(n_986),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_996),
.B(n_924),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_999),
.A2(n_886),
.B1(n_924),
.B2(n_902),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_995),
.A2(n_897),
.B1(n_881),
.B2(n_864),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1003),
.A2(n_997),
.B1(n_1002),
.B2(n_1005),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1006),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_1004),
.B(n_998),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1010),
.B(n_994),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1011),
.A2(n_1008),
.B1(n_1007),
.B2(n_891),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_1012),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_1013),
.A2(n_1009),
.B1(n_878),
.B2(n_877),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_183),
.B(n_184),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1015),
.B(n_873),
.Y(n_1017)
);

AOI222xp33_ASAP7_75t_L g1018 ( 
.A1(n_1017),
.A2(n_1016),
.B1(n_891),
.B2(n_878),
.C1(n_877),
.C2(n_882),
.Y(n_1018)
);

AOI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_1017),
.A2(n_878),
.B1(n_877),
.B2(n_873),
.C(n_874),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_1017),
.A2(n_882),
.B1(n_870),
.B2(n_866),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_866),
.B1(n_864),
.B2(n_860),
.Y(n_1021)
);

OAI221xp5_ASAP7_75t_R g1022 ( 
.A1(n_1021),
.A2(n_1019),
.B1(n_1018),
.B2(n_189),
.C(n_190),
.Y(n_1022)
);

AOI211xp5_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_186),
.B(n_188),
.C(n_192),
.Y(n_1023)
);


endmodule