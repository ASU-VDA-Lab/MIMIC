module fake_jpeg_11671_n_306 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_273;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_300;
wire n_294;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_29),
.B(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_4),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_9),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_67),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_1),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_15),
.B(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_69),
.B(n_76),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_73),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_10),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_40),
.B1(n_31),
.B2(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_91),
.B1(n_57),
.B2(n_62),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_31),
.B1(n_38),
.B2(n_37),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_82),
.A2(n_111),
.B(n_106),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_96),
.B1(n_117),
.B2(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_119),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_35),
.B1(n_18),
.B2(n_17),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_18),
.B1(n_17),
.B2(n_2),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_108),
.B(n_122),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_12),
.B1(n_19),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_42),
.A2(n_60),
.B1(n_44),
.B2(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_116),
.Y(n_147)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_2),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_45),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_48),
.B(n_2),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_3),
.B1(n_22),
.B2(n_30),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_59),
.A2(n_3),
.B1(n_30),
.B2(n_74),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_3),
.B1(n_78),
.B2(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_100),
.B1(n_127),
.B2(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_56),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_113),
.Y(n_149)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_145),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_139),
.Y(n_173)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_139),
.C(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_95),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_115),
.B1(n_85),
.B2(n_86),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_158),
.B1(n_162),
.B2(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_83),
.B1(n_113),
.B2(n_129),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_159),
.Y(n_205)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_97),
.B(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_168),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_83),
.A2(n_106),
.B1(n_102),
.B2(n_92),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_101),
.B1(n_87),
.B2(n_109),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_165),
.B1(n_131),
.B2(n_145),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_101),
.A2(n_109),
.B1(n_121),
.B2(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_67),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_171),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_133),
.B1(n_168),
.B2(n_157),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_185),
.B1(n_194),
.B2(n_151),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_198),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_140),
.B1(n_155),
.B2(n_158),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_184),
.B1(n_202),
.B2(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_144),
.B(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_190),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_147),
.C(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_136),
.B(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_161),
.B1(n_163),
.B2(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_142),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_202),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_152),
.C(n_165),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_134),
.C(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_216),
.B1(n_219),
.B2(n_228),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_164),
.B(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_226),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_194),
.B1(n_185),
.B2(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_218),
.B1(n_182),
.B2(n_195),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_193),
.B1(n_196),
.B2(n_179),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_192),
.B1(n_173),
.B2(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_203),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_192),
.B(n_190),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_205),
.B1(n_204),
.B2(n_183),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_182),
.B1(n_176),
.B2(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_186),
.Y(n_234)
);

BUFx4f_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_186),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_240),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_242),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_220),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_250),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_207),
.A2(n_195),
.B1(n_215),
.B2(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_221),
.B1(n_222),
.B2(n_230),
.Y(n_261)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_212),
.B1(n_213),
.B2(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_225),
.B(n_206),
.C(n_228),
.D(n_211),
.Y(n_256)
);

XOR2x1_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_249),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_206),
.C(n_208),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_264),
.C(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_231),
.B(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_260),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_244),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_250),
.B1(n_242),
.B2(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

AOI221xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_240),
.B1(n_232),
.B2(n_239),
.C(n_241),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_235),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_243),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_249),
.B(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_275),
.Y(n_281)
);

AOI321xp33_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_235),
.A3(n_236),
.B1(n_265),
.B2(n_259),
.C(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_257),
.C(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_284),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_254),
.B1(n_251),
.B2(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_285),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_264),
.B(n_252),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_270),
.B(n_268),
.C(n_271),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_276),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_277),
.C(n_282),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_269),
.C(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_281),
.C(n_282),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_266),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_284),
.Y(n_293)
);

XOR2x2_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_297),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_294),
.B(n_290),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_298),
.C(n_291),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_287),
.Y(n_306)
);


endmodule