module fake_ibex_1801_n_3998 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_673, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_679, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_672, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_411, n_135, n_520, n_658, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3998);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_673;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_672;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_658;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3998;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_3479;
wire n_711;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3780;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_738;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_1032;
wire n_936;
wire n_3813;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_724;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_2699;
wire n_847;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_721;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_757;
wire n_3948;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_687;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_3929;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_961;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_768;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_3139;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2433;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2494;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3655;
wire n_3543;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2148;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_3945;
wire n_763;
wire n_1882;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_683;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_483),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_88),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_254),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_100),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_437),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_285),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_11),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_20),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_221),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

BUFx10_ASAP7_75t_L g694 ( 
.A(n_635),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_652),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_74),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_589),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_524),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_34),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_525),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_267),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_74),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_423),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_658),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_54),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_229),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_533),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_520),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_215),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_195),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_342),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_493),
.Y(n_713)
);

BUFx2_ASAP7_75t_SL g714 ( 
.A(n_468),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_380),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_197),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_330),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_133),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_612),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_625),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_645),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_466),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_26),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_274),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_520),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_378),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_244),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_159),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_190),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_666),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_163),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_13),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_124),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_527),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_424),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_386),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_660),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_354),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_623),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_616),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_233),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_222),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_171),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_194),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_414),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_430),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_452),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_241),
.Y(n_748)
);

INVx4_ASAP7_75t_R g749 ( 
.A(n_363),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_239),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_460),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_655),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_330),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_27),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_528),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_82),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_559),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_99),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_109),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_229),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_109),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_135),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_495),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_621),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_217),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_441),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_479),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_127),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_639),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_586),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_494),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_82),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_39),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_129),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_554),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_491),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_649),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_593),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_626),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_636),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_501),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_274),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_418),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_318),
.Y(n_784)
);

INVxp33_ASAP7_75t_R g785 ( 
.A(n_250),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_305),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_342),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_122),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_209),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_367),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_191),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_551),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_560),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_199),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_256),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_531),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_281),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_521),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_627),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_662),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_14),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_18),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_493),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_64),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_206),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_266),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_13),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_104),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_17),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_228),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_250),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_680),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_631),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_516),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_650),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_418),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_7),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_599),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_465),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_390),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_343),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_339),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_574),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_154),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_183),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_157),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_405),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_293),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_175),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_254),
.Y(n_830)
);

BUFx10_ASAP7_75t_L g831 ( 
.A(n_578),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_517),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_595),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_173),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_90),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_526),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_64),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_443),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_609),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_678),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_276),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_339),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_509),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_455),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_584),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_359),
.Y(n_846)
);

CKINVDCx16_ASAP7_75t_R g847 ( 
.A(n_94),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_646),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_295),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_69),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_548),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_549),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_500),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_449),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_519),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_507),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_194),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_30),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_106),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_415),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_596),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_67),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_668),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_540),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_349),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_30),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_96),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_204),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_159),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_111),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_585),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_178),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_326),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_197),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_570),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_572),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_143),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_146),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_350),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_325),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_153),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_617),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_477),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_237),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_360),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_333),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_36),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_672),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_372),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_24),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_665),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_653),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_409),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_288),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_436),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_220),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_546),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_486),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_614),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_508),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_192),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_633),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_316),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_656),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_49),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_651),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_490),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_669),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_654),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_566),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_294),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_426),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_131),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_513),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_299),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_634),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_210),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_7),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_519),
.Y(n_919)
);

CKINVDCx14_ASAP7_75t_R g920 ( 
.A(n_187),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_210),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_671),
.Y(n_922)
);

BUFx5_ASAP7_75t_L g923 ( 
.A(n_452),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_316),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_514),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_6),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_467),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_168),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_504),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_663),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_485),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_72),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_407),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_363),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_491),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_353),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_201),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_304),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_103),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_12),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_174),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_73),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_270),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_131),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_528),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_379),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_239),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_199),
.Y(n_948)
);

CKINVDCx14_ASAP7_75t_R g949 ( 
.A(n_409),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_647),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_195),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_269),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_419),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_163),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_331),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_271),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_529),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_471),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_280),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_85),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_644),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_123),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_499),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_667),
.Y(n_964)
);

BUFx5_ASAP7_75t_L g965 ( 
.A(n_365),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_550),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_513),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_187),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_624),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_577),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_290),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_598),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_637),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_127),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_230),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_673),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_59),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_641),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_430),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_35),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_206),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_630),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_216),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_568),
.Y(n_984)
);

BUFx10_ASAP7_75t_L g985 ( 
.A(n_52),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_515),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_437),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_168),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_442),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_516),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_101),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_293),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_31),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_468),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_424),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_590),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_0),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_270),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_245),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_244),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_65),
.Y(n_1001)
);

BUFx8_ASAP7_75t_SL g1002 ( 
.A(n_6),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_303),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_151),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_359),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_438),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_314),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_575),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_192),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_592),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_369),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_332),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_523),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_640),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_364),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_225),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_323),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_427),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_657),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_518),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_314),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_477),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_487),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_436),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_498),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_618),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_46),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_83),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_387),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_529),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_38),
.Y(n_1031)
);

CKINVDCx16_ASAP7_75t_R g1032 ( 
.A(n_642),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_305),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_50),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_530),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_255),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_438),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_68),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_45),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_358),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_361),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_4),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_150),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_341),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_202),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_225),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_20),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_21),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_386),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_16),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_67),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_208),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_606),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_441),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_622),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_165),
.Y(n_1056)
);

BUFx10_ASAP7_75t_L g1057 ( 
.A(n_408),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_620),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_281),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_297),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_558),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_427),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_628),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_26),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_108),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_116),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_541),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_259),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_296),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_414),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_681),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_92),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_260),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_629),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_396),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_632),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_569),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_464),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_619),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_676),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_403),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_267),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_648),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_201),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_167),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_587),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_643),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_321),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_423),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_233),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_364),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_408),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_117),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_594),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_545),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_547),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_522),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_81),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_101),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_428),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_133),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_124),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_600),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_348),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_428),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_193),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_661),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_571),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_306),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_177),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_242),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_79),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_413),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_69),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_392),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_674),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_366),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_10),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_19),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_59),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_328),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_309),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_677),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_313),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_245),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_312),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_562),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_679),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_488),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_148),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_114),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_503),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_434),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_553),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_102),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_664),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_758),
.B(n_1025),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_693),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1028),
.B(n_1),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_923),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_941),
.Y(n_1142)
);

BUFx8_ASAP7_75t_SL g1143 ( 
.A(n_1002),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1067),
.B(n_0),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_693),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_806),
.B(n_2),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_923),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_772),
.B(n_3),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_773),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1067),
.B(n_2),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_693),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_693),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_694),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_699),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_847),
.B(n_3),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_719),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_694),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_689),
.B(n_4),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_920),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1032),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_694),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_941),
.Y(n_1162)
);

BUFx8_ASAP7_75t_SL g1163 ( 
.A(n_1002),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_831),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_737),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1110),
.B(n_8),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_815),
.B(n_8),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_719),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_941),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_719),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_719),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1035),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_699),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_909),
.B(n_9),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_699),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_923),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_727),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_949),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_727),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_885),
.B(n_5),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1019),
.B(n_9),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_885),
.B(n_5),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1035),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_911),
.B(n_11),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_911),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_695),
.B(n_10),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_1035),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_831),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_936),
.B(n_14),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_831),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_936),
.B(n_945),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_705),
.B(n_12),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_735),
.Y(n_1193)
);

BUFx8_ASAP7_75t_SL g1194 ( 
.A(n_746),
.Y(n_1194)
);

INVx5_ASAP7_75t_L g1195 ( 
.A(n_1035),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_802),
.Y(n_1196)
);

BUFx12f_ASAP7_75t_L g1197 ( 
.A(n_735),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_945),
.B(n_15),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_923),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1076),
.B(n_15),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_923),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_923),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_967),
.B(n_17),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_967),
.B(n_16),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_683),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_802),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_923),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_769),
.B(n_18),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_720),
.B(n_670),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1076),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_735),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_865),
.B(n_19),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_965),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1076),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_697),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1076),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_710),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_710),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1059),
.B(n_21),
.Y(n_1219)
);

BUFx8_ASAP7_75t_SL g1220 ( 
.A(n_746),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_780),
.B(n_22),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_710),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_710),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_683),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_765),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_712),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_701),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1059),
.Y(n_1228)
);

AND2x6_ASAP7_75t_L g1229 ( 
.A(n_779),
.B(n_675),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_712),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_739),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_915),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_712),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_958),
.B(n_23),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_965),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_712),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1030),
.B(n_22),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_762),
.Y(n_1238)
);

AND2x6_ASAP7_75t_L g1239 ( 
.A(n_779),
.B(n_682),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_718),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_965),
.Y(n_1241)
);

BUFx8_ASAP7_75t_SL g1242 ( 
.A(n_783),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_874),
.B(n_1119),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_718),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_690),
.B(n_23),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_723),
.Y(n_1246)
);

BUFx8_ASAP7_75t_SL g1247 ( 
.A(n_783),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_723),
.B(n_25),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_965),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_915),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_724),
.B(n_25),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_724),
.B(n_27),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_740),
.Y(n_1253)
);

AND2x6_ASAP7_75t_L g1254 ( 
.A(n_813),
.B(n_659),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_762),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_725),
.B(n_28),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_799),
.B(n_24),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_762),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_965),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_752),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_762),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_935),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_935),
.B(n_28),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1142),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1142),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1205),
.A2(n_726),
.B1(n_729),
.B2(n_725),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1224),
.A2(n_729),
.B1(n_1130),
.B2(n_726),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1173),
.B(n_937),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1138),
.A2(n_1134),
.B1(n_1136),
.B2(n_1130),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1159),
.B(n_765),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1165),
.A2(n_798),
.B1(n_900),
.B2(n_895),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1180),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1149),
.B(n_1134),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1154),
.B(n_714),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1240),
.A2(n_764),
.B1(n_775),
.B2(n_737),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1244),
.A2(n_1136),
.B1(n_775),
.B2(n_812),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1246),
.A2(n_812),
.B1(n_871),
.B2(n_764),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1162),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1160),
.A2(n_910),
.B1(n_1071),
.B2(n_871),
.Y(n_1279)
);

INVx8_ASAP7_75t_L g1280 ( 
.A(n_1197),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1157),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1180),
.A2(n_1182),
.B1(n_1204),
.B2(n_1198),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1182),
.A2(n_1071),
.B1(n_1108),
.B2(n_910),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1169),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1198),
.A2(n_1108),
.B1(n_685),
.B2(n_686),
.Y(n_1285)
);

AO22x2_ASAP7_75t_L g1286 ( 
.A1(n_1146),
.A2(n_785),
.B1(n_1133),
.B2(n_1016),
.Y(n_1286)
);

AO22x2_ASAP7_75t_L g1287 ( 
.A1(n_1155),
.A2(n_1049),
.B1(n_1075),
.B2(n_738),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1204),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1219),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1178),
.B(n_765),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1217),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1157),
.B(n_868),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1161),
.B(n_868),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1161),
.B(n_868),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1234),
.A2(n_1127),
.B1(n_895),
.B2(n_900),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1173),
.B(n_937),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1248),
.A2(n_687),
.B1(n_688),
.B2(n_684),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1263),
.A2(n_698),
.B1(n_700),
.B2(n_691),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1188),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1211),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1263),
.A2(n_1188),
.B1(n_1243),
.B2(n_1237),
.Y(n_1302)
);

AO22x2_ASAP7_75t_L g1303 ( 
.A1(n_1212),
.A2(n_1097),
.B1(n_1118),
.B2(n_1082),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1177),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1175),
.A2(n_704),
.B1(n_706),
.B2(n_703),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1245),
.A2(n_1175),
.B1(n_1225),
.B2(n_1193),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1196),
.B(n_985),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1140),
.A2(n_1127),
.B1(n_903),
.B2(n_918),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1193),
.A2(n_709),
.B1(n_711),
.B2(n_707),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1217),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1194),
.A2(n_903),
.B1(n_918),
.B2(n_798),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1217),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1251),
.A2(n_733),
.B1(n_734),
.B2(n_713),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1225),
.A2(n_741),
.B1(n_742),
.B2(n_736),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1158),
.A2(n_747),
.B1(n_748),
.B2(n_744),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1148),
.A2(n_1166),
.B1(n_1256),
.B2(n_1252),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_R g1317 ( 
.A1(n_1220),
.A2(n_696),
.B1(n_702),
.B2(n_692),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1153),
.B(n_940),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1179),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1222),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1185),
.Y(n_1321)
);

OA22x2_ASAP7_75t_L g1322 ( 
.A1(n_1228),
.A2(n_1206),
.B1(n_1250),
.B2(n_1191),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1167),
.A2(n_751),
.B1(n_753),
.B2(n_750),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1259),
.A2(n_1181),
.B1(n_1174),
.B2(n_1150),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1184),
.A2(n_760),
.B1(n_761),
.B2(n_759),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1139),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1242),
.A2(n_991),
.B1(n_1031),
.B2(n_986),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1189),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1203),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1164),
.A2(n_991),
.B1(n_1031),
.B2(n_986),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1232),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1247),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1190),
.B(n_985),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1215),
.B(n_818),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1139),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1143),
.B(n_849),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_R g1337 ( 
.A1(n_1163),
.A2(n_715),
.B1(n_717),
.B2(n_716),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_R g1339 ( 
.A1(n_1186),
.A2(n_722),
.B1(n_732),
.B2(n_731),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1227),
.B(n_840),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1209),
.A2(n_771),
.B1(n_776),
.B2(n_766),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1262),
.A2(n_1040),
.B1(n_1100),
.B2(n_1034),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1259),
.A2(n_784),
.B1(n_786),
.B2(n_782),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1222),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1192),
.A2(n_1040),
.B1(n_1100),
.B2(n_1034),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1213),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1222),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1213),
.A2(n_791),
.B1(n_794),
.B2(n_789),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1200),
.A2(n_797),
.B1(n_803),
.B2(n_795),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1144),
.A2(n_807),
.B1(n_808),
.B2(n_804),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1226),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1226),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1208),
.A2(n_1114),
.B1(n_1120),
.B2(n_1106),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1226),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1231),
.B(n_728),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1231),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1253),
.B(n_743),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1221),
.A2(n_811),
.B1(n_816),
.B2(n_809),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1257),
.A2(n_1114),
.B1(n_1120),
.B2(n_1106),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1141),
.A2(n_745),
.B1(n_755),
.B2(n_754),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1253),
.B(n_985),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1260),
.B(n_1129),
.Y(n_1362)
);

AO22x2_ASAP7_75t_L g1363 ( 
.A1(n_1147),
.A2(n_1132),
.B1(n_1126),
.B2(n_763),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1230),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1229),
.A2(n_821),
.B1(n_822),
.B2(n_817),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1260),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1176),
.B(n_861),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1199),
.B(n_1057),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1201),
.A2(n_826),
.B1(n_827),
.B2(n_824),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1202),
.B(n_1057),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1207),
.B(n_1057),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1235),
.A2(n_756),
.B1(n_768),
.B2(n_767),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1241),
.A2(n_787),
.B1(n_790),
.B2(n_788),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1249),
.A2(n_829),
.B1(n_832),
.B2(n_828),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1230),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1230),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1233),
.A2(n_837),
.B1(n_838),
.B2(n_835),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1229),
.A2(n_843),
.B1(n_844),
.B2(n_841),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1233),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1233),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1218),
.B(n_872),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1238),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1229),
.A2(n_1254),
.B1(n_1239),
.B2(n_853),
.Y(n_1383)
);

AO22x2_ASAP7_75t_L g1384 ( 
.A1(n_1229),
.A2(n_1121),
.B1(n_1115),
.B2(n_819),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1218),
.B(n_805),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1218),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1238),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1238),
.A2(n_854),
.B1(n_855),
.B2(n_850),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1145),
.B(n_1091),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1239),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1145),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1145),
.B(n_1091),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1152),
.Y(n_1393)
);

AO22x2_ASAP7_75t_L g1394 ( 
.A1(n_1239),
.A2(n_825),
.B1(n_830),
.B2(n_820),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1152),
.A2(n_836),
.B1(n_842),
.B2(n_834),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1152),
.A2(n_856),
.B1(n_859),
.B2(n_858),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1239),
.A2(n_860),
.B1(n_866),
.B2(n_862),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1156),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1156),
.A2(n_877),
.B1(n_879),
.B2(n_846),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1156),
.B(n_1129),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1170),
.A2(n_869),
.B1(n_870),
.B2(n_867),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1223),
.A2(n_878),
.B1(n_880),
.B2(n_873),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1170),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1170),
.A2(n_883),
.B1(n_884),
.B2(n_881),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1254),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1254),
.A2(n_887),
.B1(n_896),
.B2(n_893),
.Y(n_1406)
);

NOR2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1223),
.B(n_956),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1183),
.A2(n_889),
.B1(n_894),
.B2(n_886),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1183),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1183),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1187),
.Y(n_1411)
);

AO22x2_ASAP7_75t_L g1412 ( 
.A1(n_1254),
.A2(n_905),
.B1(n_921),
.B2(n_901),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1187),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1187),
.B(n_1091),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1195),
.A2(n_907),
.B1(n_912),
.B2(n_898),
.Y(n_1415)
);

AND2x2_ASAP7_75t_SL g1416 ( 
.A(n_1223),
.B(n_728),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1195),
.A2(n_931),
.B1(n_933),
.B2(n_929),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1195),
.B(n_1113),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1210),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1236),
.A2(n_914),
.B1(n_917),
.B2(n_913),
.Y(n_1420)
);

AO22x2_ASAP7_75t_L g1421 ( 
.A1(n_1210),
.A2(n_946),
.B1(n_955),
.B2(n_944),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1236),
.A2(n_924),
.B1(n_925),
.B2(n_919),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1210),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1236),
.A2(n_927),
.B1(n_928),
.B2(n_926),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1255),
.B(n_801),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1214),
.A2(n_963),
.B1(n_971),
.B2(n_959),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1255),
.B(n_975),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1214),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1214),
.B(n_1113),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1255),
.A2(n_934),
.B1(n_938),
.B2(n_932),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1258),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1258),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1258),
.B(n_1113),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1261),
.B(n_977),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1261),
.A2(n_942),
.B1(n_943),
.B2(n_939),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1261),
.B(n_1131),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1139),
.B(n_1131),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1151),
.A2(n_989),
.B1(n_992),
.B2(n_988),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1151),
.A2(n_995),
.B1(n_997),
.B2(n_993),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1151),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1168),
.A2(n_948),
.B1(n_952),
.B2(n_947),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1168),
.A2(n_1003),
.B1(n_1011),
.B2(n_1001),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1168),
.B(n_801),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1171),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1171),
.A2(n_954),
.B1(n_957),
.B2(n_953),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1171),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1172),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1172),
.A2(n_960),
.B1(n_968),
.B2(n_962),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1172),
.B(n_956),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1216),
.B(n_1017),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1216),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1216),
.Y(n_1452)
);

AO22x2_ASAP7_75t_L g1453 ( 
.A1(n_1146),
.A2(n_1020),
.B1(n_1022),
.B2(n_1015),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1205),
.A2(n_974),
.B1(n_980),
.B2(n_979),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1159),
.B(n_1017),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1138),
.A2(n_1050),
.B1(n_1060),
.B2(n_1047),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1138),
.A2(n_1065),
.B1(n_1068),
.B2(n_1064),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1159),
.B(n_1018),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1138),
.A2(n_1081),
.B1(n_1088),
.B2(n_1073),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1205),
.A2(n_981),
.B1(n_987),
.B2(n_983),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1138),
.B(n_1093),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1180),
.Y(n_1462)
);

AO22x2_ASAP7_75t_L g1463 ( 
.A1(n_1146),
.A2(n_1111),
.B1(n_1107),
.B2(n_849),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1205),
.A2(n_990),
.B1(n_998),
.B2(n_994),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1159),
.B(n_1018),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1234),
.A2(n_999),
.B1(n_1005),
.B2(n_1000),
.Y(n_1466)
);

XNOR2xp5_ASAP7_75t_L g1467 ( 
.A(n_1165),
.B(n_1006),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1157),
.B(n_720),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1180),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1159),
.B(n_1062),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1234),
.A2(n_1009),
.B1(n_1012),
.B2(n_1007),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1180),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1205),
.A2(n_1013),
.B1(n_1023),
.B2(n_1021),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1157),
.B(n_892),
.Y(n_1474)
);

AO22x2_ASAP7_75t_L g1475 ( 
.A1(n_1146),
.A2(n_857),
.B1(n_872),
.B2(n_814),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1205),
.A2(n_1024),
.B1(n_1029),
.B2(n_1027),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1138),
.A2(n_1125),
.B1(n_1123),
.B2(n_1036),
.Y(n_1477)
);

INVx8_ASAP7_75t_L g1478 ( 
.A(n_1154),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1304),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1319),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1280),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1321),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1275),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1363),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1363),
.Y(n_1486)
);

INVx3_ASAP7_75t_R g1487 ( 
.A(n_1461),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1475),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1475),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1385),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1427),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1436),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1434),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1361),
.B(n_1062),
.Y(n_1494)
);

AOI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1346),
.A2(n_916),
.B(n_908),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1264),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1265),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1279),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_R g1499 ( 
.A(n_1274),
.B(n_1033),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1437),
.Y(n_1500)
);

XNOR2xp5_ASAP7_75t_L g1501 ( 
.A(n_1283),
.B(n_1037),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1278),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1381),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1284),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1268),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1450),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1297),
.Y(n_1507)
);

XOR2xp5_ASAP7_75t_L g1508 ( 
.A(n_1467),
.B(n_1101),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1280),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1272),
.B(n_721),
.Y(n_1510)
);

INVxp33_ASAP7_75t_SL g1511 ( 
.A(n_1276),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1433),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1405),
.B(n_721),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1288),
.Y(n_1514)
);

XOR2x2_ASAP7_75t_L g1515 ( 
.A(n_1311),
.B(n_29),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_SL g1516 ( 
.A(n_1405),
.B(n_1390),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1327),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1355),
.B(n_1085),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1290),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1462),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1469),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1472),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1368),
.B(n_965),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1449),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1331),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1463),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1273),
.B(n_1038),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1463),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1292),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1310),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1307),
.B(n_1039),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1289),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1438),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1281),
.B(n_796),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1301),
.B(n_1112),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1438),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1362),
.B(n_966),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1282),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1478),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1370),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1371),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1360),
.Y(n_1542)
);

INVxp33_ASAP7_75t_L g1543 ( 
.A(n_1271),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1357),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1306),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1306),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1270),
.B(n_1041),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1407),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1291),
.B(n_1042),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1389),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1478),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1392),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1414),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1293),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1418),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1300),
.B(n_833),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1429),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1312),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1453),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1453),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1355),
.B(n_1294),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1381),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1425),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1425),
.Y(n_1564)
);

XOR2xp5_ASAP7_75t_L g1565 ( 
.A(n_1277),
.B(n_1043),
.Y(n_1565)
);

INVxp33_ASAP7_75t_L g1566 ( 
.A(n_1345),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1320),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1295),
.B(n_1044),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1421),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1366),
.B(n_1096),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1416),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1421),
.Y(n_1572)
);

XOR2xp5_ASAP7_75t_L g1573 ( 
.A(n_1332),
.B(n_1045),
.Y(n_1573)
);

INVxp33_ASAP7_75t_L g1574 ( 
.A(n_1266),
.Y(n_1574)
);

AND2x6_ASAP7_75t_L g1575 ( 
.A(n_1383),
.B(n_813),
.Y(n_1575)
);

XOR2xp5_ASAP7_75t_L g1576 ( 
.A(n_1286),
.B(n_1098),
.Y(n_1576)
);

AO21x1_ASAP7_75t_L g1577 ( 
.A1(n_1367),
.A2(n_973),
.B(n_972),
.Y(n_1577)
);

XOR2xp5_ASAP7_75t_L g1578 ( 
.A(n_1286),
.B(n_1102),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1356),
.B(n_1135),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1443),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1443),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1455),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1439),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1442),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1285),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1322),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1458),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1465),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1384),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_R g1590 ( 
.A(n_1274),
.B(n_1048),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1470),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1302),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1468),
.B(n_1338),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1344),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1267),
.B(n_1051),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1384),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1394),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1394),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1336),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1412),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1318),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1412),
.Y(n_1602)
);

XOR2xp5_ASAP7_75t_L g1603 ( 
.A(n_1330),
.B(n_1105),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1372),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1333),
.B(n_1052),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1373),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1382),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1316),
.B(n_757),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1395),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1399),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1408),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_SL g1612 ( 
.A(n_1336),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1365),
.A2(n_1397),
.B(n_1378),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1417),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1426),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1405),
.A2(n_730),
.B(n_708),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1474),
.B(n_770),
.Y(n_1617)
);

XOR2xp5_ASAP7_75t_L g1618 ( 
.A(n_1342),
.B(n_1122),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1406),
.B(n_777),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1347),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1402),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1448),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1420),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1422),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1424),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1324),
.B(n_778),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1318),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1430),
.Y(n_1628)
);

AND2x2_ASAP7_75t_SL g1629 ( 
.A(n_1343),
.B(n_814),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1435),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1391),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1393),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1308),
.B(n_1054),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1419),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1410),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1375),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1441),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1445),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1351),
.Y(n_1639)
);

XNOR2xp5_ASAP7_75t_L g1640 ( 
.A(n_1353),
.B(n_1056),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1352),
.Y(n_1641)
);

XOR2xp5_ASAP7_75t_L g1642 ( 
.A(n_1359),
.B(n_1089),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1354),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1296),
.B(n_1269),
.Y(n_1644)
);

XOR2xp5_ASAP7_75t_L g1645 ( 
.A(n_1287),
.B(n_1303),
.Y(n_1645)
);

XNOR2x2_ASAP7_75t_L g1646 ( 
.A(n_1287),
.B(n_857),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1299),
.B(n_1085),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1432),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1364),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1454),
.B(n_1460),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1376),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1379),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1380),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_SL g1654 ( 
.A(n_1317),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1387),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1398),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1369),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1374),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1464),
.B(n_1069),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1349),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1473),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1400),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1403),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1334),
.A2(n_1026),
.B(n_978),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1350),
.B(n_792),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1340),
.B(n_1055),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1409),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1411),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1476),
.Y(n_1669)
);

XOR2xp5_ASAP7_75t_L g1670 ( 
.A(n_1303),
.B(n_1116),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1413),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1423),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1428),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1323),
.B(n_1070),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1305),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1401),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1309),
.B(n_793),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1314),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1404),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1415),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1326),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1358),
.B(n_890),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1396),
.Y(n_1683)
);

XNOR2x2_ASAP7_75t_L g1684 ( 
.A(n_1339),
.B(n_890),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1377),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1388),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1446),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1431),
.Y(n_1688)
);

XOR2x2_ASAP7_75t_L g1689 ( 
.A(n_1466),
.B(n_29),
.Y(n_1689)
);

INVxp33_ASAP7_75t_L g1690 ( 
.A(n_1348),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1315),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1325),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1298),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1313),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1477),
.B(n_800),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1326),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1444),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1456),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1457),
.A2(n_1063),
.B(n_1058),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1459),
.Y(n_1700)
);

INVxp67_ASAP7_75t_SL g1701 ( 
.A(n_1471),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_R g1702 ( 
.A(n_1341),
.B(n_1072),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1386),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1440),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1335),
.B(n_823),
.Y(n_1705)
);

NAND2x1p5_ASAP7_75t_L g1706 ( 
.A(n_1335),
.B(n_940),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1337),
.B(n_1078),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1447),
.B(n_1084),
.Y(n_1708)
);

XOR2xp5_ASAP7_75t_L g1709 ( 
.A(n_1452),
.B(n_1099),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1451),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1452),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1273),
.B(n_1090),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1361),
.B(n_951),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1436),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1273),
.B(n_1092),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1328),
.B(n_839),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1328),
.B(n_845),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1273),
.B(n_1103),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1304),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1304),
.Y(n_1720)
);

XOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1467),
.B(n_31),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1304),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1328),
.B(n_965),
.Y(n_1723)
);

INVx4_ASAP7_75t_SL g1724 ( 
.A(n_1443),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1316),
.A2(n_730),
.B(n_708),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1304),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1304),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1304),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1280),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1438),
.Y(n_1730)
);

INVxp33_ASAP7_75t_SL g1731 ( 
.A(n_1275),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1436),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1304),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1304),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1273),
.B(n_951),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1273),
.B(n_1004),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1304),
.Y(n_1737)
);

XOR2xp5_ASAP7_75t_L g1738 ( 
.A(n_1467),
.B(n_32),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1304),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1304),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1280),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1273),
.B(n_1004),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1304),
.Y(n_1743)
);

NOR2xp67_ASAP7_75t_L g1744 ( 
.A(n_1282),
.B(n_537),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1304),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1273),
.B(n_1046),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1304),
.Y(n_1747)
);

CKINVDCx11_ASAP7_75t_R g1748 ( 
.A(n_1332),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1304),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1304),
.Y(n_1750)
);

INVxp33_ASAP7_75t_SL g1751 ( 
.A(n_1275),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1304),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1304),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1328),
.B(n_1087),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1289),
.Y(n_1755)
);

NOR2xp67_ASAP7_75t_L g1756 ( 
.A(n_1282),
.B(n_539),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1436),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1275),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_R g1759 ( 
.A(n_1280),
.B(n_848),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1304),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1405),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1281),
.B(n_1046),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1273),
.B(n_781),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1436),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1361),
.B(n_1137),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1304),
.Y(n_1766)
);

XNOR2x2_ASAP7_75t_L g1767 ( 
.A(n_1287),
.B(n_749),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1304),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1304),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1436),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1483),
.B(n_1109),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1538),
.B(n_1124),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1761),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1527),
.B(n_1712),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1607),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1551),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1724),
.B(n_1104),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1540),
.B(n_774),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1715),
.B(n_774),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1539),
.Y(n_1780)
);

AND2x6_ASAP7_75t_L g1781 ( 
.A(n_1533),
.B(n_1137),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1718),
.B(n_774),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1542),
.B(n_1604),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1479),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1480),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1582),
.B(n_1544),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1761),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1541),
.B(n_774),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1582),
.B(n_781),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1631),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1554),
.B(n_781),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1482),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1650),
.A2(n_1592),
.B1(n_1604),
.B2(n_1542),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1554),
.B(n_781),
.Y(n_1794)
);

AND2x2_ASAP7_75t_SL g1795 ( 
.A(n_1730),
.B(n_810),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1724),
.B(n_851),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1730),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1632),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1719),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1634),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1724),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1595),
.B(n_810),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_R g1803 ( 
.A(n_1481),
.B(n_852),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1755),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1720),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1722),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1606),
.B(n_904),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1726),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1727),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1728),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1496),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1531),
.B(n_810),
.Y(n_1812)
);

INVx3_ASAP7_75t_SL g1813 ( 
.A(n_1509),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1514),
.B(n_904),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1497),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1502),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1519),
.B(n_1080),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1633),
.B(n_1735),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1561),
.B(n_810),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1736),
.B(n_1066),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1520),
.B(n_1080),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1690),
.B(n_1698),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1733),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1734),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1700),
.B(n_863),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1648),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1521),
.B(n_864),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1601),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1742),
.B(n_1066),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1737),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1504),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1746),
.B(n_1066),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1589),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1739),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1648),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1547),
.B(n_1066),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1529),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1530),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1740),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1608),
.B(n_875),
.Y(n_1840)
);

AND2x6_ASAP7_75t_L g1841 ( 
.A(n_1536),
.B(n_532),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1522),
.B(n_876),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1743),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1761),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1745),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1549),
.B(n_32),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1659),
.B(n_33),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1747),
.Y(n_1848)
);

AND2x2_ASAP7_75t_SL g1849 ( 
.A(n_1589),
.B(n_33),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1681),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1561),
.B(n_34),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1558),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1749),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1725),
.A2(n_888),
.B(n_882),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1750),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1744),
.B(n_891),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1729),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1640),
.B(n_35),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1752),
.B(n_897),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_SL g1860 ( 
.A(n_1516),
.B(n_899),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1644),
.B(n_36),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1753),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1642),
.B(n_37),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1709),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1487),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1567),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1594),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1759),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1568),
.B(n_37),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1532),
.Y(n_1870)
);

AND2x2_ASAP7_75t_SL g1871 ( 
.A(n_1629),
.B(n_38),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1760),
.B(n_902),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1620),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1618),
.B(n_39),
.Y(n_1874)
);

AND2x6_ASAP7_75t_L g1875 ( 
.A(n_1485),
.B(n_534),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1766),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1641),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1587),
.B(n_40),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1486),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1652),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1768),
.B(n_906),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1769),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1588),
.B(n_1591),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1723),
.B(n_922),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1574),
.B(n_40),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1603),
.B(n_41),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1681),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1525),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1518),
.Y(n_1889)
);

INVxp33_ASAP7_75t_L g1890 ( 
.A(n_1535),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1723),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1512),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1663),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1518),
.Y(n_1894)
);

NAND2x1p5_ASAP7_75t_L g1895 ( 
.A(n_1503),
.B(n_41),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1681),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1754),
.B(n_930),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1763),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1526),
.Y(n_1899)
);

NOR2xp67_ASAP7_75t_L g1900 ( 
.A(n_1741),
.B(n_42),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1559),
.B(n_42),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1490),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1703),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1639),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1643),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1641),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1491),
.Y(n_1907)
);

NOR2xp67_ASAP7_75t_L g1908 ( 
.A(n_1627),
.B(n_43),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1649),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1762),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1641),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1725),
.A2(n_961),
.B(n_950),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1616),
.A2(n_969),
.B(n_964),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1762),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1484),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1651),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1528),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1696),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1653),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1635),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1493),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1754),
.B(n_970),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1748),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1609),
.B(n_976),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1599),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1550),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1758),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1605),
.B(n_43),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1647),
.B(n_44),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1560),
.B(n_44),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1647),
.B(n_45),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1683),
.B(n_982),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1503),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1622),
.B(n_984),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1552),
.Y(n_1935)
);

AND2x2_ASAP7_75t_SL g1936 ( 
.A(n_1707),
.B(n_46),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1623),
.B(n_996),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1656),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1616),
.A2(n_1010),
.B(n_1008),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1488),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1553),
.Y(n_1941)
);

BUFx5_ASAP7_75t_L g1942 ( 
.A(n_1569),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1555),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1557),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1624),
.B(n_1014),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1627),
.B(n_47),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1610),
.B(n_1611),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1495),
.A2(n_1061),
.B(n_1053),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1701),
.A2(n_1077),
.B1(n_1079),
.B2(n_1074),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1660),
.B(n_47),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1676),
.B(n_48),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1682),
.B(n_48),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1492),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1500),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1682),
.B(n_49),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1506),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1586),
.B(n_50),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1655),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1713),
.B(n_1501),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1614),
.B(n_1083),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1714),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1679),
.B(n_51),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1713),
.B(n_51),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1537),
.A2(n_1638),
.B(n_1637),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1566),
.B(n_52),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1489),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1680),
.B(n_1685),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1732),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1494),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1596),
.B(n_53),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1505),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1667),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1668),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1757),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1645),
.B(n_53),
.Y(n_1975)
);

OR2x6_ASAP7_75t_L g1976 ( 
.A(n_1691),
.B(n_54),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1615),
.B(n_1086),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1671),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_R g1979 ( 
.A(n_1499),
.B(n_1094),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1672),
.Y(n_1980)
);

INVxp67_ASAP7_75t_L g1981 ( 
.A(n_1494),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1764),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1699),
.B(n_55),
.Y(n_1983)
);

AND2x6_ASAP7_75t_L g1984 ( 
.A(n_1597),
.B(n_535),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1673),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1583),
.B(n_1095),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1584),
.B(n_1117),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1770),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1537),
.B(n_1128),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1699),
.B(n_55),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1744),
.B(n_56),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1523),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_R g1993 ( 
.A(n_1590),
.B(n_56),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1565),
.B(n_57),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1523),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1625),
.B(n_57),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1670),
.B(n_58),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1524),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1756),
.B(n_58),
.Y(n_1999)
);

NOR2xp67_ASAP7_75t_L g2000 ( 
.A(n_1693),
.B(n_60),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1510),
.Y(n_2001)
);

BUFx24_ASAP7_75t_L g2002 ( 
.A(n_1612),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1498),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1686),
.B(n_1657),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1701),
.B(n_1716),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1668),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1628),
.B(n_60),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1717),
.B(n_61),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1708),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1545),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1756),
.B(n_61),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1694),
.B(n_62),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1706),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1546),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1510),
.Y(n_2015)
);

INVx4_ASAP7_75t_L g2016 ( 
.A(n_1612),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1507),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1706),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1630),
.B(n_62),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1692),
.B(n_63),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1572),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1666),
.B(n_63),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1687),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1598),
.Y(n_2024)
);

AND2x6_ASAP7_75t_L g2025 ( 
.A(n_1600),
.B(n_536),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1658),
.B(n_66),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1666),
.B(n_65),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1687),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1543),
.B(n_66),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1621),
.B(n_68),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1688),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1508),
.B(n_70),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1664),
.B(n_70),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1662),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1664),
.B(n_71),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1548),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1619),
.B(n_72),
.Y(n_2037)
);

INVx4_ASAP7_75t_L g2038 ( 
.A(n_1765),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1562),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1636),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1563),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1564),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1580),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1602),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1516),
.B(n_71),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1593),
.B(n_73),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1577),
.B(n_75),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1613),
.B(n_75),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1697),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1613),
.B(n_76),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1765),
.B(n_1626),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1581),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1646),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1702),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1767),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_1571),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1570),
.B(n_76),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1576),
.B(n_77),
.Y(n_2058)
);

INVxp33_ASAP7_75t_L g2059 ( 
.A(n_1573),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1575),
.Y(n_2060)
);

OAI21xp33_ASAP7_75t_L g2061 ( 
.A1(n_1731),
.A2(n_1751),
.B(n_1511),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1665),
.Y(n_2062)
);

INVx3_ASAP7_75t_SL g2063 ( 
.A(n_1515),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1578),
.B(n_77),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1704),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1684),
.Y(n_2066)
);

INVx3_ASAP7_75t_L g2067 ( 
.A(n_1575),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1695),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1575),
.A2(n_543),
.B(n_542),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1575),
.B(n_78),
.Y(n_2070)
);

INVxp67_ASAP7_75t_L g2071 ( 
.A(n_1674),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1677),
.B(n_78),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1585),
.B(n_79),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1661),
.B(n_80),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1710),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1669),
.B(n_80),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1579),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1617),
.B(n_1556),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1675),
.B(n_81),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_1513),
.A2(n_1711),
.B(n_1705),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1678),
.B(n_83),
.Y(n_2081)
);

AND2x2_ASAP7_75t_SL g2082 ( 
.A(n_1654),
.B(n_84),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1571),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1689),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1534),
.B(n_84),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1654),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1721),
.B(n_85),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1738),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_1517),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1483),
.B(n_86),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1483),
.B(n_86),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1607),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1483),
.B(n_87),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1607),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1551),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1551),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1539),
.Y(n_2097)
);

NAND2x1p5_ASAP7_75t_L g2098 ( 
.A(n_1503),
.B(n_87),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1483),
.B(n_88),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1483),
.B(n_89),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1483),
.B(n_89),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1483),
.B(n_90),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1761),
.Y(n_2103)
);

BUFx4f_ASAP7_75t_L g2104 ( 
.A(n_1539),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1483),
.B(n_91),
.Y(n_2105)
);

AND2x2_ASAP7_75t_SL g2106 ( 
.A(n_1730),
.B(n_91),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1607),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1483),
.B(n_92),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1483),
.B(n_93),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1483),
.B(n_93),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1795),
.B(n_94),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1903),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2034),
.B(n_2015),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1914),
.B(n_95),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1822),
.B(n_95),
.Y(n_2115)
);

INVxp67_ASAP7_75t_SL g2116 ( 
.A(n_1797),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_SL g2117 ( 
.A(n_1850),
.B(n_544),
.Y(n_2117)
);

OR2x6_ASAP7_75t_L g2118 ( 
.A(n_1976),
.B(n_96),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2023),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1784),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1785),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1822),
.B(n_97),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1850),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_SL g2124 ( 
.A(n_1850),
.B(n_552),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_1835),
.Y(n_2125)
);

CKINVDCx14_ASAP7_75t_R g2126 ( 
.A(n_1776),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1792),
.Y(n_2127)
);

OR2x6_ASAP7_75t_L g2128 ( 
.A(n_1976),
.B(n_97),
.Y(n_2128)
);

AO21x2_ASAP7_75t_L g2129 ( 
.A1(n_2053),
.A2(n_556),
.B(n_555),
.Y(n_2129)
);

NAND2x1p5_ASAP7_75t_L g2130 ( 
.A(n_2104),
.B(n_98),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_2002),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1799),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1793),
.B(n_98),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1826),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1805),
.Y(n_2135)
);

OR2x6_ASAP7_75t_L g2136 ( 
.A(n_1976),
.B(n_99),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1818),
.B(n_100),
.Y(n_2137)
);

OR2x6_ASAP7_75t_L g2138 ( 
.A(n_1923),
.B(n_102),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2001),
.B(n_103),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2001),
.B(n_104),
.Y(n_2140)
);

BUFx12f_ASAP7_75t_L g2141 ( 
.A(n_2096),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1887),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2005),
.B(n_105),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1806),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_2061),
.B(n_105),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1808),
.Y(n_2146)
);

AND2x6_ASAP7_75t_L g2147 ( 
.A(n_1901),
.B(n_106),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1786),
.B(n_107),
.Y(n_2148)
);

NAND2x1p5_ASAP7_75t_L g2149 ( 
.A(n_2104),
.B(n_107),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_SL g2150 ( 
.A(n_1887),
.B(n_557),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1902),
.B(n_108),
.Y(n_2151)
);

OR2x6_ASAP7_75t_L g2152 ( 
.A(n_2016),
.B(n_110),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1774),
.B(n_110),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1907),
.B(n_111),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1809),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1921),
.B(n_112),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1936),
.B(n_112),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_1780),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2004),
.B(n_113),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_1826),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2004),
.B(n_113),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1858),
.B(n_114),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1887),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1890),
.B(n_115),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1967),
.B(n_115),
.Y(n_2165)
);

AND2x4_ASAP7_75t_SL g2166 ( 
.A(n_1801),
.B(n_116),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2051),
.B(n_117),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2073),
.B(n_118),
.Y(n_2168)
);

NOR2xp67_ASAP7_75t_L g2169 ( 
.A(n_2060),
.B(n_561),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2074),
.B(n_118),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_2023),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2076),
.B(n_119),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_2028),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_2097),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_1910),
.B(n_1967),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1810),
.Y(n_2176)
);

BUFx2_ASAP7_75t_SL g2177 ( 
.A(n_2016),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2079),
.B(n_119),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1823),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1824),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_2095),
.Y(n_2181)
);

NOR2xp67_ASAP7_75t_L g2182 ( 
.A(n_2060),
.B(n_563),
.Y(n_2182)
);

INVx4_ASAP7_75t_L g2183 ( 
.A(n_1813),
.Y(n_2183)
);

OR2x6_ASAP7_75t_L g2184 ( 
.A(n_1851),
.B(n_120),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1910),
.B(n_120),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1896),
.Y(n_2186)
);

AND2x4_ASAP7_75t_L g2187 ( 
.A(n_1830),
.B(n_121),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1861),
.B(n_121),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_2028),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1783),
.B(n_122),
.Y(n_2190)
);

INVx5_ASAP7_75t_L g2191 ( 
.A(n_1844),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2081),
.B(n_123),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1783),
.B(n_125),
.Y(n_2193)
);

NAND2x1p5_ASAP7_75t_L g2194 ( 
.A(n_1857),
.B(n_125),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1834),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2110),
.B(n_126),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2110),
.B(n_126),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1839),
.B(n_128),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1889),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1843),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_1845),
.B(n_128),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_SL g2202 ( 
.A(n_1896),
.B(n_564),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1896),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1848),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1871),
.B(n_129),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1927),
.B(n_130),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1927),
.B(n_130),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_1889),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1853),
.B(n_132),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1855),
.B(n_132),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1862),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_1813),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1876),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_1915),
.B(n_134),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1959),
.B(n_134),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1844),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1882),
.B(n_135),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1888),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1891),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_1894),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_1865),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1775),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_1801),
.B(n_136),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1863),
.B(n_136),
.Y(n_2224)
);

OR2x6_ASAP7_75t_L g2225 ( 
.A(n_1851),
.B(n_137),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_1870),
.B(n_137),
.Y(n_2226)
);

BUFx4f_ASAP7_75t_L g2227 ( 
.A(n_1951),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1918),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1790),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2003),
.B(n_138),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1833),
.B(n_2009),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1844),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_1894),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_1804),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1918),
.Y(n_2235)
);

AND2x2_ASAP7_75t_SL g2236 ( 
.A(n_2106),
.B(n_138),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1833),
.B(n_139),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1849),
.B(n_1886),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2093),
.B(n_139),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_2051),
.B(n_140),
.Y(n_2240)
);

INVx4_ASAP7_75t_L g2241 ( 
.A(n_1918),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_2080),
.A2(n_573),
.B(n_565),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2093),
.B(n_2109),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2103),
.Y(n_2244)
);

OR2x6_ASAP7_75t_L g2245 ( 
.A(n_1895),
.B(n_140),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1879),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1879),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1798),
.Y(n_2248)
);

INVxp67_ASAP7_75t_L g2249 ( 
.A(n_1951),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2109),
.B(n_141),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_1803),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2014),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_1864),
.B(n_141),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2014),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_2103),
.Y(n_2255)
);

AO21x2_ASAP7_75t_L g2256 ( 
.A1(n_2050),
.A2(n_579),
.B(n_576),
.Y(n_2256)
);

BUFx3_ASAP7_75t_L g2257 ( 
.A(n_1925),
.Y(n_2257)
);

NOR2x1_ASAP7_75t_L g2258 ( 
.A(n_2067),
.B(n_142),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2021),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_2103),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1800),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1975),
.B(n_142),
.Y(n_2262)
);

BUFx12f_ASAP7_75t_L g2263 ( 
.A(n_1920),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1883),
.B(n_143),
.Y(n_2264)
);

NOR2xp67_ASAP7_75t_L g2265 ( 
.A(n_2067),
.B(n_580),
.Y(n_2265)
);

OR2x6_ASAP7_75t_L g2266 ( 
.A(n_1895),
.B(n_144),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2092),
.Y(n_2267)
);

INVx5_ASAP7_75t_L g2268 ( 
.A(n_1875),
.Y(n_2268)
);

INVx2_ASAP7_75t_SL g2269 ( 
.A(n_1865),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2021),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2094),
.Y(n_2271)
);

BUFx3_ASAP7_75t_L g2272 ( 
.A(n_2086),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2107),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_1864),
.B(n_2088),
.Y(n_2274)
);

BUFx4f_ASAP7_75t_L g2275 ( 
.A(n_1962),
.Y(n_2275)
);

BUFx8_ASAP7_75t_L g2276 ( 
.A(n_1962),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2013),
.Y(n_2277)
);

INVx5_ASAP7_75t_L g2278 ( 
.A(n_1875),
.Y(n_2278)
);

BUFx2_ASAP7_75t_L g2279 ( 
.A(n_2038),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1926),
.B(n_144),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1994),
.B(n_1929),
.Y(n_2281)
);

NAND2x1_ASAP7_75t_SL g2282 ( 
.A(n_2089),
.B(n_145),
.Y(n_2282)
);

CKINVDCx8_ASAP7_75t_R g2283 ( 
.A(n_1950),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_2038),
.Y(n_2284)
);

INVx5_ASAP7_75t_L g2285 ( 
.A(n_1875),
.Y(n_2285)
);

OR2x6_ASAP7_75t_L g2286 ( 
.A(n_2098),
.B(n_145),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_1868),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1935),
.B(n_146),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2044),
.Y(n_2289)
);

INVxp67_ASAP7_75t_L g2290 ( 
.A(n_1950),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1941),
.B(n_147),
.Y(n_2291)
);

AND2x2_ASAP7_75t_SL g2292 ( 
.A(n_2082),
.B(n_147),
.Y(n_2292)
);

NAND2x1p5_ASAP7_75t_L g2293 ( 
.A(n_1868),
.B(n_148),
.Y(n_2293)
);

BUFx4f_ASAP7_75t_L g2294 ( 
.A(n_2098),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1816),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2044),
.Y(n_2296)
);

CKINVDCx11_ASAP7_75t_R g2297 ( 
.A(n_2063),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1943),
.B(n_149),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2062),
.B(n_149),
.Y(n_2299)
);

BUFx8_ASAP7_75t_SL g2300 ( 
.A(n_2054),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_1944),
.B(n_150),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1831),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2052),
.B(n_151),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_2013),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1993),
.Y(n_2305)
);

OR2x6_ASAP7_75t_SL g2306 ( 
.A(n_1874),
.B(n_152),
.Y(n_2306)
);

BUFx12f_ASAP7_75t_L g2307 ( 
.A(n_1828),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_2052),
.B(n_152),
.Y(n_2308)
);

INVx4_ASAP7_75t_L g2309 ( 
.A(n_1906),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1979),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1811),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_1931),
.B(n_153),
.Y(n_2312)
);

AND2x2_ASAP7_75t_SL g2313 ( 
.A(n_1901),
.B(n_154),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2010),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_1878),
.B(n_1892),
.Y(n_2315)
);

INVx5_ASAP7_75t_L g2316 ( 
.A(n_1875),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_2013),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1815),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1899),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2077),
.B(n_155),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1847),
.B(n_155),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1899),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1934),
.B(n_156),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2084),
.B(n_156),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1934),
.B(n_157),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_2089),
.Y(n_2326)
);

BUFx5_ASAP7_75t_L g2327 ( 
.A(n_1984),
.Y(n_2327)
);

BUFx8_ASAP7_75t_SL g2328 ( 
.A(n_2032),
.Y(n_2328)
);

OR2x6_ASAP7_75t_L g2329 ( 
.A(n_1970),
.B(n_158),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_SL g2330 ( 
.A(n_1860),
.B(n_581),
.Y(n_2330)
);

BUFx12f_ASAP7_75t_L g2331 ( 
.A(n_1819),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2066),
.B(n_158),
.Y(n_2332)
);

BUFx2_ASAP7_75t_L g2333 ( 
.A(n_1797),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_1846),
.B(n_160),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1937),
.B(n_160),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_1969),
.B(n_161),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_2083),
.Y(n_2337)
);

NAND2x1_ASAP7_75t_L g2338 ( 
.A(n_1984),
.B(n_582),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_2083),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1906),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_1937),
.B(n_161),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_1869),
.B(n_162),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_1952),
.B(n_162),
.Y(n_2343)
);

BUFx8_ASAP7_75t_L g2344 ( 
.A(n_1955),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_1930),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_SL g2346 ( 
.A(n_1860),
.B(n_583),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1945),
.B(n_164),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_1906),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_1911),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2063),
.B(n_164),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1945),
.B(n_2108),
.Y(n_2351)
);

INVxp67_ASAP7_75t_L g2352 ( 
.A(n_1930),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2056),
.Y(n_2353)
);

INVxp67_ASAP7_75t_L g2354 ( 
.A(n_1963),
.Y(n_2354)
);

INVxp67_ASAP7_75t_SL g2355 ( 
.A(n_1911),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_1819),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_1928),
.B(n_165),
.Y(n_2357)
);

INVx1_ASAP7_75t_SL g2358 ( 
.A(n_2056),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1904),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_1911),
.Y(n_2360)
);

NAND2x1p5_ASAP7_75t_L g2361 ( 
.A(n_1938),
.B(n_166),
.Y(n_2361)
);

NAND2x1p5_ASAP7_75t_L g2362 ( 
.A(n_1938),
.B(n_166),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_1773),
.Y(n_2363)
);

NAND2x1p5_ASAP7_75t_L g2364 ( 
.A(n_1971),
.B(n_167),
.Y(n_2364)
);

INVx1_ASAP7_75t_SL g2365 ( 
.A(n_1791),
.Y(n_2365)
);

NAND2x1p5_ASAP7_75t_L g2366 ( 
.A(n_1900),
.B(n_169),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1917),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_1953),
.B(n_169),
.Y(n_2368)
);

BUFx12f_ASAP7_75t_L g2369 ( 
.A(n_1997),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1917),
.Y(n_2370)
);

INVx4_ASAP7_75t_L g2371 ( 
.A(n_1984),
.Y(n_2371)
);

OR2x6_ASAP7_75t_L g2372 ( 
.A(n_1970),
.B(n_170),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_SL g2373 ( 
.A(n_1984),
.B(n_588),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_1954),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2024),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1981),
.B(n_170),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_1981),
.B(n_171),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_1956),
.B(n_172),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_2087),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2024),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2090),
.B(n_172),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_1778),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2091),
.B(n_2102),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2029),
.B(n_173),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_1933),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1772),
.B(n_174),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2055),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_1965),
.B(n_175),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_1961),
.B(n_176),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_1772),
.B(n_176),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1773),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_1968),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_1905),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_SL g2394 ( 
.A(n_2025),
.B(n_591),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_1974),
.B(n_177),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_1982),
.B(n_178),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_1909),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1940),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_2055),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2078),
.B(n_2071),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_1947),
.B(n_179),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2058),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_1988),
.B(n_179),
.Y(n_2403)
);

NAND2x1p5_ASAP7_75t_L g2404 ( 
.A(n_1787),
.B(n_180),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_SL g2405 ( 
.A(n_2025),
.B(n_597),
.Y(n_2405)
);

INVx4_ASAP7_75t_L g2406 ( 
.A(n_2025),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1947),
.B(n_180),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_1787),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2078),
.B(n_181),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1916),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2064),
.B(n_181),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1877),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1940),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2031),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1964),
.B(n_182),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_1964),
.B(n_182),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1825),
.B(n_183),
.Y(n_2417)
);

BUFx2_ASAP7_75t_L g2418 ( 
.A(n_1933),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2040),
.B(n_184),
.Y(n_2419)
);

BUFx3_ASAP7_75t_L g2420 ( 
.A(n_2039),
.Y(n_2420)
);

BUFx12f_ASAP7_75t_L g2421 ( 
.A(n_1778),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_1946),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2085),
.B(n_184),
.Y(n_2423)
);

INVxp67_ASAP7_75t_L g2424 ( 
.A(n_2099),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_1788),
.Y(n_2425)
);

BUFx2_ASAP7_75t_L g2426 ( 
.A(n_1788),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_SL g2427 ( 
.A(n_2025),
.B(n_601),
.Y(n_2427)
);

INVxp67_ASAP7_75t_L g2428 ( 
.A(n_2099),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_1919),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2030),
.B(n_185),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_1958),
.Y(n_2431)
);

INVx3_ASAP7_75t_L g2432 ( 
.A(n_2031),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_1972),
.Y(n_2433)
);

AND2x6_ASAP7_75t_L g2434 ( 
.A(n_1983),
.B(n_185),
.Y(n_2434)
);

AND2x2_ASAP7_75t_SL g2435 ( 
.A(n_1990),
.B(n_186),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_1802),
.B(n_186),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_1825),
.B(n_188),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2041),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_1978),
.Y(n_2439)
);

BUFx5_ASAP7_75t_L g2440 ( 
.A(n_1841),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2072),
.B(n_188),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_1966),
.Y(n_2442)
);

INVx2_ASAP7_75t_SL g2443 ( 
.A(n_1812),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_SL g2444 ( 
.A(n_1841),
.B(n_602),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2072),
.B(n_1771),
.Y(n_2445)
);

AND2x6_ASAP7_75t_L g2446 ( 
.A(n_1992),
.B(n_189),
.Y(n_2446)
);

AND2x4_ASAP7_75t_L g2447 ( 
.A(n_2071),
.B(n_189),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_1840),
.B(n_190),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_1973),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_1885),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1966),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1771),
.B(n_2105),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_1841),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_1877),
.Y(n_2454)
);

AND2x4_ASAP7_75t_L g2455 ( 
.A(n_2042),
.B(n_191),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1995),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2018),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_1980),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2105),
.B(n_193),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2085),
.B(n_196),
.Y(n_2460)
);

OR2x6_ASAP7_75t_L g2461 ( 
.A(n_1908),
.B(n_196),
.Y(n_2461)
);

INVxp67_ASAP7_75t_L g2462 ( 
.A(n_2100),
.Y(n_2462)
);

OR2x6_ASAP7_75t_L g2463 ( 
.A(n_1777),
.B(n_198),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2101),
.B(n_198),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_1841),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1837),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_1840),
.B(n_200),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1985),
.Y(n_2468)
);

BUFx3_ASAP7_75t_L g2469 ( 
.A(n_2043),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_1998),
.B(n_200),
.Y(n_2470)
);

NAND2x1_ASAP7_75t_L g2471 ( 
.A(n_2049),
.B(n_603),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2069),
.B(n_604),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2017),
.Y(n_2473)
);

AND2x4_ASAP7_75t_L g2474 ( 
.A(n_1898),
.B(n_202),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_SL g2475 ( 
.A(n_2069),
.B(n_605),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_1796),
.B(n_203),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_1836),
.B(n_203),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_1924),
.B(n_1960),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_1973),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_1781),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2100),
.B(n_204),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2101),
.B(n_205),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_1779),
.B(n_205),
.Y(n_2483)
);

NOR2x1_ASAP7_75t_L g2484 ( 
.A(n_2050),
.B(n_207),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1838),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_1781),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1852),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_1866),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_1867),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1996),
.B(n_207),
.Y(n_2490)
);

INVx4_ASAP7_75t_L g2491 ( 
.A(n_1781),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1996),
.B(n_208),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_1924),
.B(n_209),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_1960),
.B(n_211),
.Y(n_2494)
);

INVx4_ASAP7_75t_L g2495 ( 
.A(n_1781),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2007),
.B(n_211),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1873),
.Y(n_2497)
);

INVx2_ASAP7_75t_SL g2498 ( 
.A(n_1782),
.Y(n_2498)
);

INVxp67_ASAP7_75t_L g2499 ( 
.A(n_2037),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_1794),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_1880),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2070),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_1893),
.Y(n_2503)
);

BUFx8_ASAP7_75t_L g2504 ( 
.A(n_2012),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2006),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1814),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2007),
.B(n_212),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_1957),
.B(n_212),
.Y(n_2508)
);

INVxp67_ASAP7_75t_L g2509 ( 
.A(n_2037),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_1814),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_1817),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2019),
.B(n_213),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_1942),
.Y(n_2513)
);

BUFx8_ASAP7_75t_L g2514 ( 
.A(n_2020),
.Y(n_2514)
);

BUFx2_ASAP7_75t_L g2515 ( 
.A(n_2070),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2068),
.B(n_213),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_1989),
.B(n_214),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1817),
.Y(n_2518)
);

INVxp67_ASAP7_75t_SL g2519 ( 
.A(n_2022),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2036),
.B(n_214),
.Y(n_2520)
);

BUFx2_ASAP7_75t_SL g2521 ( 
.A(n_2000),
.Y(n_2521)
);

NAND2x1p5_ASAP7_75t_L g2522 ( 
.A(n_1789),
.B(n_215),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1821),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_1989),
.B(n_216),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2008),
.B(n_217),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2019),
.B(n_218),
.Y(n_2526)
);

NAND2x1_ASAP7_75t_L g2527 ( 
.A(n_2065),
.B(n_607),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2075),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_1977),
.B(n_2026),
.Y(n_2529)
);

BUFx4f_ASAP7_75t_L g2530 ( 
.A(n_2057),
.Y(n_2530)
);

INVxp67_ASAP7_75t_L g2531 ( 
.A(n_2026),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_1820),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_1977),
.B(n_218),
.Y(n_2533)
);

NAND2x1p5_ASAP7_75t_L g2534 ( 
.A(n_1829),
.B(n_219),
.Y(n_2534)
);

INVx1_ASAP7_75t_SL g2535 ( 
.A(n_1832),
.Y(n_2535)
);

BUFx2_ASAP7_75t_SL g2536 ( 
.A(n_1942),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_1856),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2046),
.B(n_219),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_1942),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_1991),
.Y(n_2540)
);

INVx4_ASAP7_75t_L g2541 ( 
.A(n_1942),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1942),
.Y(n_2542)
);

AND2x6_ASAP7_75t_L g2543 ( 
.A(n_2033),
.B(n_220),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1821),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1807),
.Y(n_2545)
);

OR2x2_ASAP7_75t_L g2546 ( 
.A(n_2059),
.B(n_221),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_1897),
.B(n_222),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_1807),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_SL g2549 ( 
.A(n_2033),
.B(n_608),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2047),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_2022),
.B(n_223),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_1986),
.B(n_223),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_1897),
.B(n_224),
.Y(n_2553)
);

AND2x4_ASAP7_75t_L g2554 ( 
.A(n_1999),
.B(n_224),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2035),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_2045),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2011),
.B(n_226),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_1986),
.B(n_226),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_1854),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_1987),
.B(n_227),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2035),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_1827),
.B(n_227),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2047),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_1987),
.B(n_228),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2027),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_1922),
.B(n_230),
.Y(n_2566)
);

AND2x6_ASAP7_75t_L g2567 ( 
.A(n_2027),
.B(n_231),
.Y(n_2567)
);

BUFx12f_ASAP7_75t_L g2568 ( 
.A(n_1949),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_1922),
.B(n_231),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2048),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_1827),
.B(n_232),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_1859),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1884),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_1842),
.B(n_232),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_SL g2575 ( 
.A(n_1948),
.B(n_610),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2219),
.Y(n_2576)
);

INVx2_ASAP7_75t_SL g2577 ( 
.A(n_2131),
.Y(n_2577)
);

INVx2_ASAP7_75t_SL g2578 ( 
.A(n_2212),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2125),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2236),
.B(n_1932),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2219),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2435),
.B(n_1932),
.Y(n_2582)
);

INVx5_ASAP7_75t_L g2583 ( 
.A(n_2118),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2158),
.Y(n_2584)
);

AO21x2_ASAP7_75t_L g2585 ( 
.A1(n_2415),
.A2(n_1948),
.B(n_1912),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2123),
.Y(n_2586)
);

INVx3_ASAP7_75t_L g2587 ( 
.A(n_2371),
.Y(n_2587)
);

INVx6_ASAP7_75t_SL g2588 ( 
.A(n_2118),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2294),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2456),
.Y(n_2590)
);

CKINVDCx20_ASAP7_75t_R g2591 ( 
.A(n_2251),
.Y(n_2591)
);

BUFx24_ASAP7_75t_L g2592 ( 
.A(n_2223),
.Y(n_2592)
);

NAND2x1p5_ASAP7_75t_L g2593 ( 
.A(n_2183),
.B(n_1859),
.Y(n_2593)
);

INVx8_ASAP7_75t_L g2594 ( 
.A(n_2128),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2478),
.B(n_1842),
.Y(n_2595)
);

INVxp67_ASAP7_75t_SL g2596 ( 
.A(n_2276),
.Y(n_2596)
);

BUFx12f_ASAP7_75t_L g2597 ( 
.A(n_2141),
.Y(n_2597)
);

NAND2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2183),
.B(n_1872),
.Y(n_2598)
);

INVx2_ASAP7_75t_SL g2599 ( 
.A(n_2294),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2456),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2113),
.Y(n_2601)
);

CKINVDCx20_ASAP7_75t_R g2602 ( 
.A(n_2126),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2113),
.B(n_1872),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2314),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2371),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2123),
.Y(n_2606)
);

BUFx3_ASAP7_75t_L g2607 ( 
.A(n_2257),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2406),
.B(n_1881),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2263),
.Y(n_2609)
);

NAND2x1p5_ASAP7_75t_L g2610 ( 
.A(n_2227),
.B(n_1881),
.Y(n_2610)
);

BUFx2_ASAP7_75t_SL g2611 ( 
.A(n_2268),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2134),
.Y(n_2612)
);

NAND2x1p5_ASAP7_75t_L g2613 ( 
.A(n_2227),
.B(n_1884),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2313),
.A2(n_1912),
.B1(n_1854),
.B2(n_1913),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2297),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2160),
.Y(n_2616)
);

INVxp67_ASAP7_75t_SL g2617 ( 
.A(n_2276),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2353),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2314),
.Y(n_2619)
);

BUFx2_ASAP7_75t_R g2620 ( 
.A(n_2310),
.Y(n_2620)
);

INVx5_ASAP7_75t_L g2621 ( 
.A(n_2128),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2123),
.Y(n_2622)
);

BUFx12f_ASAP7_75t_L g2623 ( 
.A(n_2138),
.Y(n_2623)
);

BUFx4f_ASAP7_75t_SL g2624 ( 
.A(n_2307),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2112),
.Y(n_2625)
);

BUFx12f_ASAP7_75t_L g2626 ( 
.A(n_2138),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2120),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2136),
.Y(n_2628)
);

CKINVDCx16_ASAP7_75t_R g2629 ( 
.A(n_2136),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2181),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2272),
.Y(n_2631)
);

INVx5_ASAP7_75t_SL g2632 ( 
.A(n_2152),
.Y(n_2632)
);

INVx4_ASAP7_75t_L g2633 ( 
.A(n_2245),
.Y(n_2633)
);

INVx5_ASAP7_75t_L g2634 ( 
.A(n_2245),
.Y(n_2634)
);

AND2x4_ASAP7_75t_L g2635 ( 
.A(n_2406),
.B(n_1913),
.Y(n_2635)
);

AOI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2292),
.A2(n_1939),
.B1(n_236),
.B2(n_234),
.Y(n_2636)
);

NAND2x1p5_ASAP7_75t_L g2637 ( 
.A(n_2275),
.B(n_234),
.Y(n_2637)
);

BUFx6f_ASAP7_75t_L g2638 ( 
.A(n_2142),
.Y(n_2638)
);

INVxp67_ASAP7_75t_SL g2639 ( 
.A(n_2275),
.Y(n_2639)
);

BUFx2_ASAP7_75t_L g2640 ( 
.A(n_2331),
.Y(n_2640)
);

INVx8_ASAP7_75t_L g2641 ( 
.A(n_2152),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2135),
.Y(n_2642)
);

BUFx8_ASAP7_75t_L g2643 ( 
.A(n_2221),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_2142),
.Y(n_2644)
);

BUFx3_ASAP7_75t_L g2645 ( 
.A(n_2374),
.Y(n_2645)
);

INVx2_ASAP7_75t_SL g2646 ( 
.A(n_2166),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2453),
.Y(n_2647)
);

INVx4_ASAP7_75t_L g2648 ( 
.A(n_2266),
.Y(n_2648)
);

BUFx3_ASAP7_75t_L g2649 ( 
.A(n_2392),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2120),
.Y(n_2650)
);

INVx2_ASAP7_75t_SL g2651 ( 
.A(n_2266),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2234),
.Y(n_2652)
);

AO21x2_ASAP7_75t_L g2653 ( 
.A1(n_2416),
.A2(n_1939),
.B(n_613),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2121),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2400),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2655)
);

BUFx12f_ASAP7_75t_L g2656 ( 
.A(n_2305),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_2142),
.Y(n_2657)
);

BUFx2_ASAP7_75t_SL g2658 ( 
.A(n_2268),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2121),
.Y(n_2659)
);

INVx1_ASAP7_75t_SL g2660 ( 
.A(n_2353),
.Y(n_2660)
);

INVx2_ASAP7_75t_SL g2661 ( 
.A(n_2286),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2144),
.Y(n_2662)
);

BUFx3_ASAP7_75t_L g2663 ( 
.A(n_2421),
.Y(n_2663)
);

BUFx2_ASAP7_75t_L g2664 ( 
.A(n_2184),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2146),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2127),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2269),
.Y(n_2667)
);

INVx4_ASAP7_75t_L g2668 ( 
.A(n_2286),
.Y(n_2668)
);

BUFx4f_ASAP7_75t_L g2669 ( 
.A(n_2147),
.Y(n_2669)
);

INVx6_ASAP7_75t_SL g2670 ( 
.A(n_2184),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2195),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2281),
.B(n_235),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2163),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2453),
.Y(n_2674)
);

INVx2_ASAP7_75t_SL g2675 ( 
.A(n_2223),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2200),
.Y(n_2676)
);

INVxp67_ASAP7_75t_SL g2677 ( 
.A(n_2139),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2127),
.Y(n_2678)
);

BUFx5_ASAP7_75t_L g2679 ( 
.A(n_2446),
.Y(n_2679)
);

INVx3_ASAP7_75t_SL g2680 ( 
.A(n_2225),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2132),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2328),
.Y(n_2682)
);

BUFx12f_ASAP7_75t_L g2683 ( 
.A(n_2326),
.Y(n_2683)
);

BUFx4f_ASAP7_75t_SL g2684 ( 
.A(n_2369),
.Y(n_2684)
);

BUFx8_ASAP7_75t_L g2685 ( 
.A(n_2157),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2225),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_2686)
);

CKINVDCx20_ASAP7_75t_R g2687 ( 
.A(n_2300),
.Y(n_2687)
);

BUFx3_ASAP7_75t_L g2688 ( 
.A(n_2191),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_SL g2689 ( 
.A(n_2283),
.B(n_238),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2238),
.B(n_240),
.Y(n_2690)
);

INVx1_ASAP7_75t_SL g2691 ( 
.A(n_2358),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2191),
.Y(n_2692)
);

BUFx3_ASAP7_75t_L g2693 ( 
.A(n_2191),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2237),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2531),
.B(n_242),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2177),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2333),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2132),
.Y(n_2698)
);

BUFx2_ASAP7_75t_SL g2699 ( 
.A(n_2268),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2155),
.Y(n_2700)
);

BUFx2_ASAP7_75t_R g2701 ( 
.A(n_2306),
.Y(n_2701)
);

NAND2x1p5_ASAP7_75t_L g2702 ( 
.A(n_2358),
.B(n_243),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2274),
.B(n_243),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2155),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2163),
.Y(n_2705)
);

BUFx6f_ASAP7_75t_L g2706 ( 
.A(n_2163),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2249),
.B(n_246),
.Y(n_2707)
);

BUFx5_ASAP7_75t_L g2708 ( 
.A(n_2446),
.Y(n_2708)
);

BUFx12f_ASAP7_75t_L g2709 ( 
.A(n_2130),
.Y(n_2709)
);

INVx3_ASAP7_75t_SL g2710 ( 
.A(n_2387),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2237),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2211),
.Y(n_2712)
);

INVx2_ASAP7_75t_SL g2713 ( 
.A(n_2231),
.Y(n_2713)
);

BUFx3_ASAP7_75t_L g2714 ( 
.A(n_2241),
.Y(n_2714)
);

INVx8_ASAP7_75t_L g2715 ( 
.A(n_2147),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2445),
.B(n_246),
.Y(n_2716)
);

BUFx8_ASAP7_75t_L g2717 ( 
.A(n_2287),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_2572),
.B(n_2278),
.Y(n_2718)
);

INVx6_ASAP7_75t_SL g2719 ( 
.A(n_2329),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2213),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2176),
.Y(n_2721)
);

INVx4_ASAP7_75t_L g2722 ( 
.A(n_2147),
.Y(n_2722)
);

INVx4_ASAP7_75t_L g2723 ( 
.A(n_2147),
.Y(n_2723)
);

INVx3_ASAP7_75t_SL g2724 ( 
.A(n_2399),
.Y(n_2724)
);

NOR2xp67_ASAP7_75t_L g2725 ( 
.A(n_2174),
.B(n_2568),
.Y(n_2725)
);

NAND2x1p5_ASAP7_75t_L g2726 ( 
.A(n_2491),
.B(n_247),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2243),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2290),
.B(n_248),
.Y(n_2728)
);

CKINVDCx16_ASAP7_75t_R g2729 ( 
.A(n_2329),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2176),
.Y(n_2730)
);

BUFx12f_ASAP7_75t_L g2731 ( 
.A(n_2149),
.Y(n_2731)
);

BUFx2_ASAP7_75t_L g2732 ( 
.A(n_2116),
.Y(n_2732)
);

BUFx12f_ASAP7_75t_L g2733 ( 
.A(n_2194),
.Y(n_2733)
);

BUFx2_ASAP7_75t_SL g2734 ( 
.A(n_2278),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2179),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2222),
.Y(n_2736)
);

INVx8_ASAP7_75t_L g2737 ( 
.A(n_2372),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_2186),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2229),
.Y(n_2739)
);

BUFx5_ASAP7_75t_L g2740 ( 
.A(n_2446),
.Y(n_2740)
);

INVx2_ASAP7_75t_SL g2741 ( 
.A(n_2231),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2179),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2180),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2541),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2241),
.Y(n_2745)
);

BUFx12f_ASAP7_75t_L g2746 ( 
.A(n_2350),
.Y(n_2746)
);

BUFx3_ASAP7_75t_L g2747 ( 
.A(n_2379),
.Y(n_2747)
);

INVx1_ASAP7_75t_SL g2748 ( 
.A(n_2185),
.Y(n_2748)
);

INVx8_ASAP7_75t_L g2749 ( 
.A(n_2372),
.Y(n_2749)
);

BUFx12f_ASAP7_75t_L g2750 ( 
.A(n_2546),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2186),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2262),
.B(n_249),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2248),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2228),
.Y(n_2754)
);

BUFx6f_ASAP7_75t_L g2755 ( 
.A(n_2186),
.Y(n_2755)
);

BUFx5_ASAP7_75t_L g2756 ( 
.A(n_2446),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2450),
.B(n_251),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2137),
.B(n_251),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2203),
.Y(n_2759)
);

INVx4_ASAP7_75t_L g2760 ( 
.A(n_2278),
.Y(n_2760)
);

BUFx2_ASAP7_75t_SL g2761 ( 
.A(n_2285),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2139),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2573),
.B(n_252),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2180),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_SL g2765 ( 
.A(n_2447),
.Y(n_2765)
);

BUFx2_ASAP7_75t_SL g2766 ( 
.A(n_2285),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2228),
.Y(n_2767)
);

INVx1_ASAP7_75t_SL g2768 ( 
.A(n_2185),
.Y(n_2768)
);

INVx5_ASAP7_75t_L g2769 ( 
.A(n_2216),
.Y(n_2769)
);

INVx1_ASAP7_75t_SL g2770 ( 
.A(n_2474),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2204),
.Y(n_2771)
);

BUFx5_ASAP7_75t_L g2772 ( 
.A(n_2289),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2203),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2204),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2175),
.Y(n_2775)
);

BUFx6f_ASAP7_75t_L g2776 ( 
.A(n_2203),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2215),
.A2(n_255),
.B1(n_252),
.B2(n_253),
.Y(n_2777)
);

BUFx12f_ASAP7_75t_L g2778 ( 
.A(n_2253),
.Y(n_2778)
);

INVx2_ASAP7_75t_SL g2779 ( 
.A(n_2364),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2175),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2205),
.B(n_253),
.Y(n_2781)
);

INVx2_ASAP7_75t_SL g2782 ( 
.A(n_2303),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2218),
.Y(n_2783)
);

BUFx2_ASAP7_75t_L g2784 ( 
.A(n_2434),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2216),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2285),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2218),
.Y(n_2787)
);

BUFx2_ASAP7_75t_SL g2788 ( 
.A(n_2316),
.Y(n_2788)
);

INVx2_ASAP7_75t_SL g2789 ( 
.A(n_2303),
.Y(n_2789)
);

BUFx12f_ASAP7_75t_L g2790 ( 
.A(n_2344),
.Y(n_2790)
);

BUFx2_ASAP7_75t_L g2791 ( 
.A(n_2434),
.Y(n_2791)
);

BUFx2_ASAP7_75t_R g2792 ( 
.A(n_2402),
.Y(n_2792)
);

INVx5_ASAP7_75t_L g2793 ( 
.A(n_2216),
.Y(n_2793)
);

INVxp67_ASAP7_75t_SL g2794 ( 
.A(n_2419),
.Y(n_2794)
);

INVx1_ASAP7_75t_SL g2795 ( 
.A(n_2474),
.Y(n_2795)
);

INVx4_ASAP7_75t_L g2796 ( 
.A(n_2316),
.Y(n_2796)
);

INVx8_ASAP7_75t_L g2797 ( 
.A(n_2187),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2261),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_SL g2799 ( 
.A(n_2447),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2232),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2235),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2573),
.B(n_2452),
.Y(n_2802)
);

INVx5_ASAP7_75t_L g2803 ( 
.A(n_2232),
.Y(n_2803)
);

CKINVDCx20_ASAP7_75t_R g2804 ( 
.A(n_2344),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2529),
.B(n_256),
.Y(n_2805)
);

BUFx3_ASAP7_75t_L g2806 ( 
.A(n_2235),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2466),
.Y(n_2807)
);

BUFx12f_ASAP7_75t_L g2808 ( 
.A(n_2214),
.Y(n_2808)
);

BUFx3_ASAP7_75t_L g2809 ( 
.A(n_2279),
.Y(n_2809)
);

BUFx3_ASAP7_75t_L g2810 ( 
.A(n_2284),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2434),
.Y(n_2811)
);

BUFx12f_ASAP7_75t_L g2812 ( 
.A(n_2230),
.Y(n_2812)
);

BUFx10_ASAP7_75t_L g2813 ( 
.A(n_2226),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2316),
.B(n_257),
.Y(n_2814)
);

INVx2_ASAP7_75t_SL g2815 ( 
.A(n_2308),
.Y(n_2815)
);

BUFx3_ASAP7_75t_L g2816 ( 
.A(n_2420),
.Y(n_2816)
);

AND2x2_ASAP7_75t_SL g2817 ( 
.A(n_2373),
.B(n_257),
.Y(n_2817)
);

BUFx12f_ASAP7_75t_L g2818 ( 
.A(n_2361),
.Y(n_2818)
);

BUFx2_ASAP7_75t_SL g2819 ( 
.A(n_2327),
.Y(n_2819)
);

CKINVDCx20_ASAP7_75t_R g2820 ( 
.A(n_2504),
.Y(n_2820)
);

INVx4_ASAP7_75t_L g2821 ( 
.A(n_2434),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2267),
.Y(n_2822)
);

INVx1_ASAP7_75t_SL g2823 ( 
.A(n_2308),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2466),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2487),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2541),
.Y(n_2826)
);

BUFx5_ASAP7_75t_L g2827 ( 
.A(n_2289),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2487),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2491),
.Y(n_2829)
);

INVx2_ASAP7_75t_SL g2830 ( 
.A(n_2114),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2153),
.B(n_258),
.Y(n_2831)
);

CKINVDCx20_ASAP7_75t_R g2832 ( 
.A(n_2504),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2438),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2271),
.Y(n_2834)
);

BUFx2_ASAP7_75t_R g2835 ( 
.A(n_2111),
.Y(n_2835)
);

NAND2x1p5_ASAP7_75t_L g2836 ( 
.A(n_2495),
.B(n_258),
.Y(n_2836)
);

INVx1_ASAP7_75t_SL g2837 ( 
.A(n_2368),
.Y(n_2837)
);

INVx3_ASAP7_75t_L g2838 ( 
.A(n_2495),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2273),
.Y(n_2839)
);

CKINVDCx6p67_ASAP7_75t_R g2840 ( 
.A(n_2461),
.Y(n_2840)
);

INVx4_ASAP7_75t_L g2841 ( 
.A(n_2232),
.Y(n_2841)
);

INVxp67_ASAP7_75t_L g2842 ( 
.A(n_2187),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2345),
.B(n_259),
.Y(n_2843)
);

INVx1_ASAP7_75t_SL g2844 ( 
.A(n_2368),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2295),
.Y(n_2845)
);

INVx3_ASAP7_75t_SL g2846 ( 
.A(n_2198),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2488),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2148),
.B(n_260),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2255),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2469),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2385),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2302),
.Y(n_2852)
);

BUFx12f_ASAP7_75t_L g2853 ( 
.A(n_2362),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2418),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2465),
.Y(n_2855)
);

INVx4_ASAP7_75t_L g2856 ( 
.A(n_2255),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2567),
.Y(n_2857)
);

BUFx8_ASAP7_75t_L g2858 ( 
.A(n_2324),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2224),
.B(n_261),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2311),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2488),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2473),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2351),
.B(n_261),
.Y(n_2863)
);

INVx5_ASAP7_75t_L g2864 ( 
.A(n_2255),
.Y(n_2864)
);

INVx8_ASAP7_75t_L g2865 ( 
.A(n_2198),
.Y(n_2865)
);

INVx6_ASAP7_75t_SL g2866 ( 
.A(n_2463),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_2340),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2465),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2114),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2545),
.Y(n_2870)
);

BUFx3_ASAP7_75t_L g2871 ( 
.A(n_2378),
.Y(n_2871)
);

BUFx4_ASAP7_75t_SL g2872 ( 
.A(n_2463),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2411),
.B(n_262),
.Y(n_2873)
);

CKINVDCx8_ASAP7_75t_R g2874 ( 
.A(n_2521),
.Y(n_2874)
);

INVx1_ASAP7_75t_SL g2875 ( 
.A(n_2378),
.Y(n_2875)
);

INVx5_ASAP7_75t_L g2876 ( 
.A(n_2465),
.Y(n_2876)
);

INVxp67_ASAP7_75t_SL g2877 ( 
.A(n_2419),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2545),
.Y(n_2878)
);

INVx2_ASAP7_75t_SL g2879 ( 
.A(n_2389),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2389),
.Y(n_2880)
);

NAND2x1p5_ASAP7_75t_L g2881 ( 
.A(n_2356),
.B(n_262),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2318),
.Y(n_2882)
);

INVx1_ASAP7_75t_SL g2883 ( 
.A(n_2395),
.Y(n_2883)
);

INVx3_ASAP7_75t_L g2884 ( 
.A(n_2486),
.Y(n_2884)
);

INVx4_ASAP7_75t_L g2885 ( 
.A(n_2486),
.Y(n_2885)
);

INVx2_ASAP7_75t_SL g2886 ( 
.A(n_2395),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2340),
.Y(n_2887)
);

INVx3_ASAP7_75t_L g2888 ( 
.A(n_2486),
.Y(n_2888)
);

BUFx8_ASAP7_75t_L g2889 ( 
.A(n_2206),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2168),
.B(n_263),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2499),
.B(n_263),
.Y(n_2891)
);

INVx4_ASAP7_75t_L g2892 ( 
.A(n_2201),
.Y(n_2892)
);

CKINVDCx16_ASAP7_75t_R g2893 ( 
.A(n_2373),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2170),
.B(n_264),
.Y(n_2894)
);

BUFx3_ASAP7_75t_L g2895 ( 
.A(n_2396),
.Y(n_2895)
);

INVx1_ASAP7_75t_SL g2896 ( 
.A(n_2396),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2309),
.Y(n_2897)
);

BUFx5_ASAP7_75t_L g2898 ( 
.A(n_2296),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2309),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2548),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2403),
.Y(n_2901)
);

INVx3_ASAP7_75t_L g2902 ( 
.A(n_2479),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2201),
.Y(n_2903)
);

INVx3_ASAP7_75t_SL g2904 ( 
.A(n_2301),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2509),
.B(n_264),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2359),
.Y(n_2906)
);

BUFx6f_ASAP7_75t_L g2907 ( 
.A(n_2340),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2348),
.Y(n_2908)
);

INVx8_ASAP7_75t_L g2909 ( 
.A(n_2301),
.Y(n_2909)
);

INVx5_ASAP7_75t_L g2910 ( 
.A(n_2348),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2479),
.Y(n_2911)
);

CKINVDCx20_ASAP7_75t_R g2912 ( 
.A(n_2514),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_2315),
.B(n_265),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2403),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2548),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2226),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2567),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2514),
.Y(n_2918)
);

INVx8_ASAP7_75t_L g2919 ( 
.A(n_2455),
.Y(n_2919)
);

INVx1_ASAP7_75t_SL g2920 ( 
.A(n_2455),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2348),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2461),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2506),
.Y(n_2923)
);

INVx1_ASAP7_75t_SL g2924 ( 
.A(n_2460),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2315),
.B(n_265),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_SL g2926 ( 
.A1(n_2293),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.Y(n_2926)
);

CKINVDCx20_ASAP7_75t_R g2927 ( 
.A(n_2207),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2424),
.B(n_268),
.Y(n_2928)
);

BUFx3_ASAP7_75t_L g2929 ( 
.A(n_2520),
.Y(n_2929)
);

BUFx8_ASAP7_75t_SL g2930 ( 
.A(n_2520),
.Y(n_2930)
);

INVx3_ASAP7_75t_SL g2931 ( 
.A(n_2516),
.Y(n_2931)
);

AND2x4_ASAP7_75t_L g2932 ( 
.A(n_2506),
.B(n_271),
.Y(n_2932)
);

CKINVDCx20_ASAP7_75t_R g2933 ( 
.A(n_2199),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_2567),
.Y(n_2934)
);

BUFx4f_ASAP7_75t_SL g2935 ( 
.A(n_2476),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2510),
.Y(n_2936)
);

BUFx3_ASAP7_75t_L g2937 ( 
.A(n_2337),
.Y(n_2937)
);

BUFx2_ASAP7_75t_L g2938 ( 
.A(n_2567),
.Y(n_2938)
);

INVx4_ASAP7_75t_L g2939 ( 
.A(n_2349),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2339),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2208),
.Y(n_2941)
);

BUFx8_ASAP7_75t_L g2942 ( 
.A(n_2476),
.Y(n_2942)
);

BUFx2_ASAP7_75t_L g2943 ( 
.A(n_2534),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_SL g2944 ( 
.A(n_2516),
.Y(n_2944)
);

INVx3_ASAP7_75t_L g2945 ( 
.A(n_2479),
.Y(n_2945)
);

INVx3_ASAP7_75t_L g2946 ( 
.A(n_2513),
.Y(n_2946)
);

INVxp67_ASAP7_75t_SL g2947 ( 
.A(n_2352),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2510),
.Y(n_2948)
);

NAND2x1p5_ASAP7_75t_L g2949 ( 
.A(n_2480),
.B(n_272),
.Y(n_2949)
);

CKINVDCx11_ASAP7_75t_R g2950 ( 
.A(n_2299),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2404),
.Y(n_2951)
);

BUFx2_ASAP7_75t_L g2952 ( 
.A(n_2477),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2349),
.Y(n_2953)
);

BUFx2_ASAP7_75t_SL g2954 ( 
.A(n_2327),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2511),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2477),
.Y(n_2956)
);

CKINVDCx20_ASAP7_75t_R g2957 ( 
.A(n_2220),
.Y(n_2957)
);

CKINVDCx11_ASAP7_75t_R g2958 ( 
.A(n_2299),
.Y(n_2958)
);

NAND2x1_ASAP7_75t_L g2959 ( 
.A(n_2244),
.B(n_611),
.Y(n_2959)
);

INVx1_ASAP7_75t_SL g2960 ( 
.A(n_2172),
.Y(n_2960)
);

INVx1_ASAP7_75t_SL g2961 ( 
.A(n_2178),
.Y(n_2961)
);

BUFx3_ASAP7_75t_L g2962 ( 
.A(n_2393),
.Y(n_2962)
);

CKINVDCx20_ASAP7_75t_R g2963 ( 
.A(n_2820),
.Y(n_2963)
);

INVxp67_ASAP7_75t_SL g2964 ( 
.A(n_2794),
.Y(n_2964)
);

OAI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2729),
.A2(n_2394),
.B1(n_2427),
.B2(n_2405),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2604),
.Y(n_2966)
);

CKINVDCx11_ASAP7_75t_R g2967 ( 
.A(n_2597),
.Y(n_2967)
);

AOI22xp33_ASAP7_75t_SL g2968 ( 
.A1(n_2935),
.A2(n_2405),
.B1(n_2427),
.B2(n_2394),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2604),
.Y(n_2969)
);

BUFx2_ASAP7_75t_L g2970 ( 
.A(n_2719),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2582),
.A2(n_2648),
.B1(n_2668),
.B2(n_2633),
.Y(n_2971)
);

AOI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_2633),
.A2(n_2448),
.B1(n_2145),
.B2(n_2543),
.Y(n_2972)
);

BUFx12f_ASAP7_75t_L g2973 ( 
.A(n_2790),
.Y(n_2973)
);

BUFx12f_ASAP7_75t_L g2974 ( 
.A(n_2615),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2669),
.A2(n_2519),
.B1(n_2530),
.B2(n_2383),
.Y(n_2975)
);

OAI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2669),
.A2(n_2530),
.B1(n_2525),
.B2(n_2342),
.Y(n_2976)
);

INVx1_ASAP7_75t_SL g2977 ( 
.A(n_2696),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2648),
.A2(n_2543),
.B1(n_2409),
.B2(n_2538),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_L g2979 ( 
.A1(n_2668),
.A2(n_2543),
.B1(n_2538),
.B2(n_2493),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2642),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2662),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2893),
.A2(n_2821),
.B1(n_2634),
.B2(n_2817),
.Y(n_2982)
);

INVx2_ASAP7_75t_SL g2983 ( 
.A(n_2737),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2580),
.A2(n_2543),
.B1(n_2494),
.B2(n_2467),
.Y(n_2984)
);

INVxp67_ASAP7_75t_SL g2985 ( 
.A(n_2877),
.Y(n_2985)
);

AND2x4_ASAP7_75t_L g2986 ( 
.A(n_2821),
.B(n_2246),
.Y(n_2986)
);

BUFx8_ASAP7_75t_SL g2987 ( 
.A(n_2602),
.Y(n_2987)
);

NAND2x1p5_ASAP7_75t_L g2988 ( 
.A(n_2634),
.B(n_2338),
.Y(n_2988)
);

AOI22xp33_ASAP7_75t_L g2989 ( 
.A1(n_2634),
.A2(n_2562),
.B1(n_2574),
.B2(n_2571),
.Y(n_2989)
);

OAI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2893),
.A2(n_2525),
.B1(n_2342),
.B2(n_2357),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2737),
.A2(n_2571),
.B1(n_2574),
.B2(n_2562),
.Y(n_2991)
);

OAI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2629),
.A2(n_2444),
.B1(n_2475),
.B2(n_2472),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2619),
.Y(n_2993)
);

OAI22xp33_ASAP7_75t_L g2994 ( 
.A1(n_2749),
.A2(n_2444),
.B1(n_2475),
.B2(n_2472),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2749),
.A2(n_2357),
.B1(n_2334),
.B2(n_2554),
.Y(n_2995)
);

AOI22xp33_ASAP7_75t_L g2996 ( 
.A1(n_2942),
.A2(n_2334),
.B1(n_2557),
.B2(n_2554),
.Y(n_2996)
);

BUFx12f_ASAP7_75t_L g2997 ( 
.A(n_2918),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2592),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2665),
.Y(n_2999)
);

BUFx2_ASAP7_75t_SL g3000 ( 
.A(n_2832),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2619),
.Y(n_3001)
);

INVx1_ASAP7_75t_SL g3002 ( 
.A(n_2933),
.Y(n_3002)
);

BUFx8_ASAP7_75t_SL g3003 ( 
.A(n_2804),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2942),
.A2(n_2557),
.B1(n_2240),
.B2(n_2167),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2732),
.B(n_2192),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2866),
.A2(n_2561),
.B1(n_2462),
.B2(n_2428),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2866),
.A2(n_2162),
.B1(n_2423),
.B2(n_2325),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2627),
.Y(n_3008)
);

AOI22xp33_ASAP7_75t_L g3009 ( 
.A1(n_2719),
.A2(n_2335),
.B1(n_2341),
.B2(n_2323),
.Y(n_3009)
);

OAI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2722),
.A2(n_2511),
.B1(n_2523),
.B2(n_2518),
.Y(n_3010)
);

HB1xp67_ASAP7_75t_L g3011 ( 
.A(n_2697),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2671),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2676),
.Y(n_3013)
);

CKINVDCx11_ASAP7_75t_R g3014 ( 
.A(n_2912),
.Y(n_3014)
);

INVx4_ASAP7_75t_L g3015 ( 
.A(n_2715),
.Y(n_3015)
);

CKINVDCx11_ASAP7_75t_R g3016 ( 
.A(n_2687),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2712),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2624),
.Y(n_3018)
);

AOI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2594),
.A2(n_2347),
.B1(n_2565),
.B2(n_2164),
.Y(n_3019)
);

OAI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2840),
.A2(n_2904),
.B1(n_2846),
.B2(n_2621),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2594),
.A2(n_2515),
.B1(n_2502),
.B2(n_2559),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2588),
.A2(n_2524),
.B1(n_2517),
.B2(n_2547),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2627),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2720),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_SL g3025 ( 
.A1(n_2715),
.A2(n_2575),
.B1(n_2327),
.B2(n_2440),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2576),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2650),
.Y(n_3027)
);

INVx8_ASAP7_75t_L g3028 ( 
.A(n_2641),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_2872),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2650),
.Y(n_3030)
);

OAI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2722),
.A2(n_2518),
.B1(n_2544),
.B2(n_2523),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2576),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2677),
.A2(n_2549),
.B(n_2346),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2802),
.B(n_2133),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2723),
.A2(n_2544),
.B1(n_2522),
.B2(n_2551),
.Y(n_3035)
);

INVx6_ASAP7_75t_L g3036 ( 
.A(n_2717),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2581),
.Y(n_3037)
);

BUFx4f_ASAP7_75t_SL g3038 ( 
.A(n_2588),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2586),
.Y(n_3039)
);

BUFx2_ASAP7_75t_L g3040 ( 
.A(n_2643),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2723),
.A2(n_2765),
.B1(n_2799),
.B2(n_2614),
.Y(n_3041)
);

INVx8_ASAP7_75t_L g3042 ( 
.A(n_2641),
.Y(n_3042)
);

OAI22xp33_ASAP7_75t_L g3043 ( 
.A1(n_2583),
.A2(n_2575),
.B1(n_2332),
.B2(n_2196),
.Y(n_3043)
);

AOI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_2583),
.A2(n_2553),
.B1(n_2555),
.B2(n_2483),
.Y(n_3044)
);

OAI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_2765),
.A2(n_2365),
.B1(n_2483),
.B2(n_2197),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2799),
.A2(n_2535),
.B1(n_2239),
.B2(n_2250),
.Y(n_3046)
);

CKINVDCx20_ASAP7_75t_R g3047 ( 
.A(n_2591),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2581),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2607),
.Y(n_3049)
);

OAI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2583),
.A2(n_2569),
.B1(n_2366),
.B2(n_2330),
.Y(n_3050)
);

BUFx2_ASAP7_75t_L g3051 ( 
.A(n_2643),
.Y(n_3051)
);

INVx8_ASAP7_75t_L g3052 ( 
.A(n_2623),
.Y(n_3052)
);

CKINVDCx11_ASAP7_75t_R g3053 ( 
.A(n_2656),
.Y(n_3053)
);

INVx6_ASAP7_75t_L g3054 ( 
.A(n_2717),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2621),
.A2(n_2555),
.B1(n_2384),
.B2(n_2388),
.Y(n_3055)
);

INVxp67_ASAP7_75t_L g3056 ( 
.A(n_2930),
.Y(n_3056)
);

OAI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2621),
.A2(n_2330),
.B1(n_2346),
.B2(n_2140),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_2670),
.A2(n_2417),
.B1(n_2437),
.B2(n_2550),
.Y(n_3058)
);

BUFx2_ASAP7_75t_L g3059 ( 
.A(n_2670),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2654),
.Y(n_3060)
);

AOI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_2950),
.A2(n_2563),
.B1(n_2484),
.B2(n_2441),
.Y(n_3061)
);

INVx3_ASAP7_75t_L g3062 ( 
.A(n_2587),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2603),
.A2(n_2354),
.B1(n_2422),
.B2(n_2343),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2958),
.A2(n_2484),
.B1(n_2321),
.B2(n_2122),
.Y(n_3064)
);

INVx6_ASAP7_75t_L g3065 ( 
.A(n_2818),
.Y(n_3065)
);

BUFx2_ASAP7_75t_SL g3066 ( 
.A(n_2609),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2654),
.Y(n_3067)
);

AOI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_2603),
.A2(n_2115),
.B1(n_2390),
.B2(n_2386),
.Y(n_3068)
);

OAI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2689),
.A2(n_2549),
.B1(n_2159),
.B2(n_2165),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2590),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2659),
.Y(n_3071)
);

INVx3_ASAP7_75t_L g3072 ( 
.A(n_2587),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_2636),
.A2(n_2312),
.B1(n_2552),
.B2(n_2533),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2659),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2590),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2666),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2816),
.Y(n_3077)
);

CKINVDCx11_ASAP7_75t_R g3078 ( 
.A(n_2683),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2600),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_2944),
.A2(n_2558),
.B1(n_2564),
.B2(n_2560),
.Y(n_3080)
);

OAI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2892),
.A2(n_2903),
.B1(n_2944),
.B2(n_2931),
.Y(n_3081)
);

OAI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2680),
.A2(n_2161),
.B1(n_2188),
.B2(n_2264),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2666),
.Y(n_3083)
);

INVx6_ASAP7_75t_L g3084 ( 
.A(n_2853),
.Y(n_3084)
);

CKINVDCx5p33_ASAP7_75t_R g3085 ( 
.A(n_2626),
.Y(n_3085)
);

BUFx8_ASAP7_75t_L g3086 ( 
.A(n_2709),
.Y(n_3086)
);

BUFx10_ASAP7_75t_L g3087 ( 
.A(n_2589),
.Y(n_3087)
);

AOI22xp33_ASAP7_75t_L g3088 ( 
.A1(n_2628),
.A2(n_2913),
.B1(n_2664),
.B2(n_2632),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2678),
.Y(n_3089)
);

OAI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_2892),
.A2(n_2903),
.B1(n_2961),
.B2(n_2960),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2797),
.A2(n_2909),
.B1(n_2919),
.B2(n_2865),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_SL g3092 ( 
.A(n_2792),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2913),
.A2(n_2566),
.B1(n_2430),
.B2(n_2498),
.Y(n_3093)
);

BUFx10_ASAP7_75t_L g3094 ( 
.A(n_2599),
.Y(n_3094)
);

OAI22x1_ASAP7_75t_L g3095 ( 
.A1(n_2922),
.A2(n_2651),
.B1(n_2661),
.B2(n_2686),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_2632),
.A2(n_2443),
.B1(n_2492),
.B2(n_2490),
.Y(n_3096)
);

BUFx12f_ASAP7_75t_L g3097 ( 
.A(n_2731),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_2595),
.A2(n_2507),
.B1(n_2512),
.B2(n_2496),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2678),
.Y(n_3099)
);

BUFx10_ASAP7_75t_L g3100 ( 
.A(n_2577),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2681),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2784),
.A2(n_2526),
.B1(n_2508),
.B2(n_2540),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2672),
.B(n_2397),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2681),
.Y(n_3104)
);

INVx2_ASAP7_75t_SL g3105 ( 
.A(n_2645),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2698),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_L g3107 ( 
.A1(n_2791),
.A2(n_2532),
.B1(n_2436),
.B2(n_2143),
.Y(n_3107)
);

INVx6_ASAP7_75t_L g3108 ( 
.A(n_2733),
.Y(n_3108)
);

BUFx3_ASAP7_75t_L g3109 ( 
.A(n_2833),
.Y(n_3109)
);

AOI22xp33_ASAP7_75t_L g3110 ( 
.A1(n_2811),
.A2(n_2440),
.B1(n_2327),
.B2(n_2500),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2698),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2778),
.A2(n_2440),
.B1(n_2327),
.B2(n_2426),
.Y(n_3112)
);

OAI22xp5_ASAP7_75t_L g3113 ( 
.A1(n_2797),
.A2(n_2535),
.B1(n_2425),
.B2(n_2381),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2700),
.Y(n_3114)
);

OAI21xp5_ASAP7_75t_SL g3115 ( 
.A1(n_2637),
.A2(n_2258),
.B(n_2376),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_2932),
.A2(n_2440),
.B1(n_2320),
.B2(n_2377),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2600),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2700),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2682),
.Y(n_3119)
);

BUFx2_ASAP7_75t_L g3120 ( 
.A(n_2850),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2704),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2704),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_SL g3123 ( 
.A1(n_2865),
.A2(n_2440),
.B1(n_2536),
.B2(n_2233),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2625),
.Y(n_3124)
);

OAI22xp5_ASAP7_75t_L g3125 ( 
.A1(n_2909),
.A2(n_2193),
.B1(n_2190),
.B2(n_2382),
.Y(n_3125)
);

BUFx3_ASAP7_75t_L g3126 ( 
.A(n_2862),
.Y(n_3126)
);

CKINVDCx6p67_ASAP7_75t_R g3127 ( 
.A(n_2663),
.Y(n_3127)
);

INVx6_ASAP7_75t_L g3128 ( 
.A(n_2649),
.Y(n_3128)
);

INVx8_ASAP7_75t_L g3129 ( 
.A(n_2919),
.Y(n_3129)
);

AOI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_2927),
.A2(n_2470),
.B1(n_2247),
.B2(n_2252),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_2616),
.B(n_2410),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2932),
.A2(n_2956),
.B1(n_2952),
.B2(n_2690),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2736),
.Y(n_3133)
);

INVx6_ASAP7_75t_L g3134 ( 
.A(n_2631),
.Y(n_3134)
);

BUFx10_ASAP7_75t_L g3135 ( 
.A(n_2814),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_2586),
.Y(n_3136)
);

CKINVDCx6p67_ASAP7_75t_R g3137 ( 
.A(n_2710),
.Y(n_3137)
);

BUFx2_ASAP7_75t_L g3138 ( 
.A(n_2957),
.Y(n_3138)
);

BUFx2_ASAP7_75t_L g3139 ( 
.A(n_2593),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2920),
.A2(n_2464),
.B1(n_2481),
.B2(n_2459),
.Y(n_3140)
);

AOI22xp33_ASAP7_75t_L g3141 ( 
.A1(n_2750),
.A2(n_2482),
.B1(n_2570),
.B2(n_2407),
.Y(n_3141)
);

OAI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2929),
.A2(n_2247),
.B1(n_2252),
.B2(n_2246),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2586),
.Y(n_3143)
);

AOI22xp33_ASAP7_75t_SL g3144 ( 
.A1(n_2916),
.A2(n_2129),
.B1(n_2259),
.B2(n_2254),
.Y(n_3144)
);

BUFx8_ASAP7_75t_SL g3145 ( 
.A(n_2640),
.Y(n_3145)
);

INVx3_ASAP7_75t_L g3146 ( 
.A(n_2605),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2739),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2753),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2721),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_2652),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2721),
.Y(n_3151)
);

BUFx8_ASAP7_75t_L g3152 ( 
.A(n_2747),
.Y(n_3152)
);

BUFx2_ASAP7_75t_L g3153 ( 
.A(n_2598),
.Y(n_3153)
);

BUFx2_ASAP7_75t_L g3154 ( 
.A(n_2809),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2606),
.Y(n_3155)
);

AOI21xp33_ASAP7_75t_L g3156 ( 
.A1(n_2608),
.A2(n_2401),
.B(n_2288),
.Y(n_3156)
);

BUFx8_ASAP7_75t_L g3157 ( 
.A(n_2943),
.Y(n_3157)
);

AOI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_2808),
.A2(n_2259),
.B1(n_2270),
.B2(n_2254),
.Y(n_3158)
);

BUFx3_ASAP7_75t_L g3159 ( 
.A(n_2684),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_2812),
.A2(n_2762),
.B1(n_2608),
.B2(n_2871),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2895),
.A2(n_2781),
.B1(n_2886),
.B2(n_2879),
.Y(n_3161)
);

BUFx3_ASAP7_75t_L g3162 ( 
.A(n_2630),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_SL g3163 ( 
.A1(n_2679),
.A2(n_2129),
.B1(n_2319),
.B2(n_2270),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2730),
.Y(n_3164)
);

CKINVDCx11_ASAP7_75t_R g3165 ( 
.A(n_2874),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_2606),
.Y(n_3166)
);

INVx6_ASAP7_75t_L g3167 ( 
.A(n_2685),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2730),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2735),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_2837),
.A2(n_2322),
.B1(n_2367),
.B2(n_2319),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2578),
.Y(n_3171)
);

BUFx2_ASAP7_75t_L g3172 ( 
.A(n_2810),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2606),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2798),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2735),
.Y(n_3175)
);

INVx6_ASAP7_75t_L g3176 ( 
.A(n_2685),
.Y(n_3176)
);

INVx6_ASAP7_75t_L g3177 ( 
.A(n_2889),
.Y(n_3177)
);

INVx2_ASAP7_75t_SL g3178 ( 
.A(n_2667),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2844),
.A2(n_2880),
.B1(n_2883),
.B2(n_2875),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2742),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_2901),
.A2(n_2694),
.B1(n_2711),
.B2(n_2635),
.Y(n_3181)
);

BUFx2_ASAP7_75t_R g3182 ( 
.A(n_2724),
.Y(n_3182)
);

BUFx12f_ASAP7_75t_L g3183 ( 
.A(n_2646),
.Y(n_3183)
);

CKINVDCx20_ASAP7_75t_R g3184 ( 
.A(n_2889),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_L g3185 ( 
.A1(n_2635),
.A2(n_2322),
.B1(n_2370),
.B2(n_2367),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2822),
.Y(n_3186)
);

INVx6_ASAP7_75t_L g3187 ( 
.A(n_2858),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2834),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2742),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_SL g3190 ( 
.A1(n_2679),
.A2(n_2370),
.B1(n_2380),
.B2(n_2375),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2839),
.Y(n_3191)
);

AOI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_2752),
.A2(n_2375),
.B1(n_2398),
.B2(n_2380),
.Y(n_3192)
);

OAI22xp33_ASAP7_75t_SL g3193 ( 
.A1(n_2702),
.A2(n_2258),
.B1(n_2413),
.B2(n_2398),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2743),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2743),
.Y(n_3195)
);

INVx1_ASAP7_75t_SL g3196 ( 
.A(n_2584),
.Y(n_3196)
);

CKINVDCx20_ASAP7_75t_R g3197 ( 
.A(n_2858),
.Y(n_3197)
);

INVxp67_ASAP7_75t_SL g3198 ( 
.A(n_2675),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2845),
.Y(n_3199)
);

BUFx4_ASAP7_75t_R g3200 ( 
.A(n_2679),
.Y(n_3200)
);

OAI22xp5_ASAP7_75t_L g3201 ( 
.A1(n_2896),
.A2(n_2914),
.B1(n_2795),
.B2(n_2770),
.Y(n_3201)
);

BUFx2_ASAP7_75t_SL g3202 ( 
.A(n_2596),
.Y(n_3202)
);

INVx6_ASAP7_75t_L g3203 ( 
.A(n_2688),
.Y(n_3203)
);

INVx6_ASAP7_75t_L g3204 ( 
.A(n_2692),
.Y(n_3204)
);

CKINVDCx6p67_ASAP7_75t_R g3205 ( 
.A(n_2951),
.Y(n_3205)
);

OAI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_2805),
.A2(n_2154),
.B(n_2151),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2870),
.B(n_2413),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2764),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2852),
.Y(n_3209)
);

OAI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_2823),
.A2(n_2442),
.B1(n_2451),
.B2(n_2156),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2713),
.B(n_2429),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2764),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2771),
.Y(n_3213)
);

NAND2x1p5_ASAP7_75t_L g3214 ( 
.A(n_2693),
.B(n_2244),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2771),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2860),
.Y(n_3216)
);

NAND2x1p5_ASAP7_75t_L g3217 ( 
.A(n_2769),
.B(n_2793),
.Y(n_3217)
);

INVx6_ASAP7_75t_L g3218 ( 
.A(n_2714),
.Y(n_3218)
);

BUFx6f_ASAP7_75t_L g3219 ( 
.A(n_2622),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_L g3220 ( 
.A(n_2622),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_2859),
.A2(n_2451),
.B1(n_2442),
.B2(n_2291),
.Y(n_3221)
);

BUFx3_ASAP7_75t_L g3222 ( 
.A(n_2745),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_2873),
.A2(n_2298),
.B1(n_2280),
.B2(n_2210),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2882),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2620),
.Y(n_3225)
);

NAND2x1p5_ASAP7_75t_L g3226 ( 
.A(n_2769),
.B(n_2260),
.Y(n_3226)
);

BUFx2_ASAP7_75t_L g3227 ( 
.A(n_2639),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2741),
.B(n_2431),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2774),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_SL g3230 ( 
.A1(n_2617),
.A2(n_2537),
.B1(n_2282),
.B2(n_2336),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2774),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_2842),
.A2(n_2217),
.B1(n_2209),
.B2(n_2296),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2783),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2906),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_L g3235 ( 
.A1(n_2890),
.A2(n_2439),
.B1(n_2458),
.B2(n_2433),
.Y(n_3235)
);

INVx6_ASAP7_75t_L g3236 ( 
.A(n_2813),
.Y(n_3236)
);

CKINVDCx11_ASAP7_75t_R g3237 ( 
.A(n_2746),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2783),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2870),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2787),
.Y(n_3240)
);

CKINVDCx6p67_ASAP7_75t_R g3241 ( 
.A(n_2611),
.Y(n_3241)
);

BUFx12f_ASAP7_75t_L g3242 ( 
.A(n_2813),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2787),
.Y(n_3243)
);

INVx4_ASAP7_75t_SL g3244 ( 
.A(n_2814),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_2894),
.A2(n_2468),
.B1(n_2432),
.B2(n_2414),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2878),
.Y(n_3246)
);

AOI22xp33_ASAP7_75t_L g3247 ( 
.A1(n_2926),
.A2(n_2432),
.B1(n_2414),
.B2(n_2489),
.Y(n_3247)
);

INVx1_ASAP7_75t_SL g3248 ( 
.A(n_2618),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_2937),
.Y(n_3249)
);

OAI21xp33_ASAP7_75t_SL g3250 ( 
.A1(n_2878),
.A2(n_2182),
.B(n_2169),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2900),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_2940),
.Y(n_3252)
);

OAI21xp5_ASAP7_75t_SL g3253 ( 
.A1(n_2726),
.A2(n_2539),
.B(n_2513),
.Y(n_3253)
);

INVx6_ASAP7_75t_L g3254 ( 
.A(n_2769),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2830),
.A2(n_2503),
.B1(n_2489),
.B2(n_2556),
.Y(n_3255)
);

BUFx5_ASAP7_75t_L g3256 ( 
.A(n_2807),
.Y(n_3256)
);

OAI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_2782),
.A2(n_2182),
.B1(n_2169),
.B2(n_2503),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_2900),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_SL g3259 ( 
.A1(n_2679),
.A2(n_2256),
.B1(n_2539),
.B2(n_2556),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_2990),
.A2(n_2984),
.B1(n_3082),
.B2(n_3156),
.Y(n_3260)
);

AOI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_2989),
.A2(n_2727),
.B1(n_2740),
.B2(n_2708),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2966),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3005),
.B(n_2915),
.Y(n_3263)
);

OAI22xp5_ASAP7_75t_SL g3264 ( 
.A1(n_2998),
.A2(n_3184),
.B1(n_3197),
.B2(n_3176),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_SL g3265 ( 
.A1(n_3167),
.A2(n_2701),
.B1(n_2779),
.B2(n_2881),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3103),
.B(n_2915),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3073),
.A2(n_2740),
.B1(n_2756),
.B2(n_2708),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_SL g3268 ( 
.A1(n_3167),
.A2(n_2757),
.B1(n_2949),
.B2(n_2836),
.Y(n_3268)
);

OAI21xp5_ASAP7_75t_SL g3269 ( 
.A1(n_2968),
.A2(n_2917),
.B(n_2857),
.Y(n_3269)
);

OAI22xp5_ASAP7_75t_L g3270 ( 
.A1(n_2965),
.A2(n_2938),
.B1(n_2934),
.B2(n_2768),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_SL g3271 ( 
.A1(n_2982),
.A2(n_2740),
.B1(n_2756),
.B2(n_2708),
.Y(n_3271)
);

OAI222xp33_ASAP7_75t_L g3272 ( 
.A1(n_3041),
.A2(n_2748),
.B1(n_2789),
.B2(n_2815),
.C1(n_2777),
.C2(n_2691),
.Y(n_3272)
);

OAI21xp33_ASAP7_75t_L g3273 ( 
.A1(n_3009),
.A2(n_2655),
.B(n_2924),
.Y(n_3273)
);

OAI22xp5_ASAP7_75t_SL g3274 ( 
.A1(n_3176),
.A2(n_2703),
.B1(n_2610),
.B2(n_2869),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_3002),
.B(n_2579),
.Y(n_3275)
);

INVx3_ASAP7_75t_SL g3276 ( 
.A(n_3065),
.Y(n_3276)
);

OAI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2994),
.A2(n_2936),
.B1(n_2948),
.B2(n_2923),
.Y(n_3277)
);

INVx3_ASAP7_75t_L g3278 ( 
.A(n_3217),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_SL g3279 ( 
.A1(n_2976),
.A2(n_2740),
.B1(n_2756),
.B2(n_2708),
.Y(n_3279)
);

INVx6_ASAP7_75t_L g3280 ( 
.A(n_3086),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2996),
.A2(n_2756),
.B1(n_2780),
.B2(n_2775),
.Y(n_3281)
);

OAI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_2991),
.A2(n_2854),
.B1(n_2851),
.B2(n_2835),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2980),
.Y(n_3283)
);

AOI22xp33_ASAP7_75t_L g3284 ( 
.A1(n_3004),
.A2(n_2831),
.B1(n_2758),
.B2(n_2728),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_SL g3285 ( 
.A1(n_3035),
.A2(n_2611),
.B1(n_2699),
.B2(n_2658),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2966),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2981),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_2978),
.A2(n_2843),
.B1(n_2707),
.B2(n_2601),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2995),
.A2(n_2660),
.B1(n_2936),
.B2(n_2923),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2999),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3125),
.A2(n_2585),
.B1(n_2716),
.B2(n_2948),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2993),
.B(n_2955),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_L g3293 ( 
.A1(n_2979),
.A2(n_2955),
.B1(n_2863),
.B2(n_2905),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3012),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3131),
.B(n_2612),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2969),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2969),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3046),
.A2(n_2972),
.B1(n_2975),
.B2(n_3095),
.Y(n_3298)
);

AOI22xp33_ASAP7_75t_L g3299 ( 
.A1(n_3068),
.A2(n_2891),
.B1(n_2925),
.B2(n_2695),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_L g3300 ( 
.A1(n_3064),
.A2(n_2941),
.B1(n_2962),
.B2(n_2848),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_SL g3301 ( 
.A1(n_3090),
.A2(n_2699),
.B1(n_2734),
.B2(n_2658),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3022),
.A2(n_2928),
.B1(n_2725),
.B2(n_2763),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_3241),
.Y(n_3303)
);

NAND3xp33_ASAP7_75t_L g3304 ( 
.A(n_3058),
.B(n_3144),
.C(n_3061),
.Y(n_3304)
);

BUFx4f_ASAP7_75t_SL g3305 ( 
.A(n_3086),
.Y(n_3305)
);

AOI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_3140),
.A2(n_2718),
.B1(n_2947),
.B2(n_2613),
.Y(n_3306)
);

AOI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_3232),
.A2(n_2718),
.B1(n_2824),
.B2(n_2807),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_3015),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3060),
.Y(n_3309)
);

INVx4_ASAP7_75t_L g3310 ( 
.A(n_3129),
.Y(n_3310)
);

AOI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_3247),
.A2(n_2825),
.B1(n_2828),
.B2(n_2824),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3001),
.B(n_2825),
.Y(n_3312)
);

AOI211xp5_ASAP7_75t_L g3313 ( 
.A1(n_3230),
.A2(n_3020),
.B(n_3050),
.C(n_3045),
.Y(n_3313)
);

OAI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_2992),
.A2(n_2847),
.B1(n_2861),
.B2(n_2828),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_3154),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3172),
.B(n_2847),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3060),
.Y(n_3317)
);

NOR2x1_ASAP7_75t_L g3318 ( 
.A(n_3040),
.B(n_2760),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3093),
.A2(n_2861),
.B1(n_2556),
.B2(n_2647),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3013),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_SL g3321 ( 
.A1(n_3135),
.A2(n_2761),
.B1(n_2766),
.B2(n_2734),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3017),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3067),
.Y(n_3323)
);

AOI222xp33_ASAP7_75t_L g3324 ( 
.A1(n_3038),
.A2(n_2674),
.B1(n_2605),
.B2(n_2647),
.C1(n_2786),
.C2(n_2760),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3067),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3071),
.Y(n_3326)
);

INVxp33_ASAP7_75t_L g3327 ( 
.A(n_3003),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3008),
.B(n_2754),
.Y(n_3328)
);

OAI21xp33_ASAP7_75t_L g3329 ( 
.A1(n_3130),
.A2(n_2801),
.B(n_2767),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3098),
.A2(n_2674),
.B1(n_2766),
.B2(n_2761),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3024),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3019),
.A2(n_2788),
.B1(n_2827),
.B2(n_2772),
.Y(n_3332)
);

HB1xp67_ASAP7_75t_L g3333 ( 
.A(n_3011),
.Y(n_3333)
);

OAI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3132),
.A2(n_2788),
.B1(n_2826),
.B2(n_2744),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3055),
.A2(n_2827),
.B1(n_2898),
.B2(n_2772),
.Y(n_3335)
);

BUFx6f_ASAP7_75t_L g3336 ( 
.A(n_3222),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3080),
.A2(n_2827),
.B1(n_2898),
.B2(n_2772),
.Y(n_3337)
);

AOI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_3044),
.A2(n_2827),
.B1(n_2898),
.B2(n_2772),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_SL g3339 ( 
.A1(n_3135),
.A2(n_2954),
.B1(n_2819),
.B2(n_2786),
.Y(n_3339)
);

OAI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3006),
.A2(n_2826),
.B1(n_2744),
.B2(n_2819),
.Y(n_3340)
);

INVx2_ASAP7_75t_SL g3341 ( 
.A(n_3065),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3023),
.B(n_3027),
.Y(n_3342)
);

AOI22xp33_ASAP7_75t_L g3343 ( 
.A1(n_3007),
.A2(n_2898),
.B1(n_2653),
.B2(n_2796),
.Y(n_3343)
);

AOI22xp33_ASAP7_75t_L g3344 ( 
.A1(n_3138),
.A2(n_2796),
.B1(n_2505),
.B2(n_2897),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3010),
.A2(n_2505),
.B1(n_2899),
.B2(n_2897),
.Y(n_3345)
);

BUFx8_ASAP7_75t_SL g3346 ( 
.A(n_2973),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_SL g3347 ( 
.A1(n_3193),
.A2(n_2954),
.B1(n_2829),
.B2(n_2838),
.Y(n_3347)
);

BUFx4f_ASAP7_75t_SL g3348 ( 
.A(n_3097),
.Y(n_3348)
);

OAI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3206),
.A2(n_2242),
.B(n_2265),
.Y(n_3349)
);

BUFx12f_ASAP7_75t_L g3350 ( 
.A(n_2967),
.Y(n_3350)
);

CKINVDCx11_ASAP7_75t_R g3351 ( 
.A(n_3016),
.Y(n_3351)
);

BUFx2_ASAP7_75t_L g3352 ( 
.A(n_3244),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3124),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3030),
.B(n_2806),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_3021),
.A2(n_2838),
.B1(n_2829),
.B2(n_2899),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3244),
.Y(n_3356)
);

OAI211xp5_ASAP7_75t_SL g3357 ( 
.A1(n_3088),
.A2(n_2449),
.B(n_2171),
.C(n_2173),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_3031),
.A2(n_2119),
.B1(n_2173),
.B2(n_2171),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3071),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3113),
.A2(n_2119),
.B1(n_2189),
.B2(n_2946),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3102),
.A2(n_2189),
.B1(n_2946),
.B2(n_2449),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3074),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3074),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3211),
.B(n_272),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3133),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3076),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_3223),
.A2(n_2256),
.B1(n_2497),
.B2(n_2485),
.Y(n_3367)
);

OAI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_3192),
.A2(n_2876),
.B1(n_2803),
.B2(n_2864),
.Y(n_3368)
);

OAI222xp33_ASAP7_75t_L g3369 ( 
.A1(n_3092),
.A2(n_3142),
.B1(n_3190),
.B2(n_3227),
.C1(n_2985),
.C2(n_2964),
.Y(n_3369)
);

OAI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3015),
.A2(n_2876),
.B1(n_2885),
.B2(n_2803),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3083),
.B(n_2902),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3089),
.B(n_2902),
.Y(n_3372)
);

OAI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3025),
.A2(n_2876),
.B1(n_2868),
.B2(n_2855),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3228),
.B(n_273),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_3129),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3076),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3111),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3185),
.A2(n_3033),
.B1(n_3116),
.B2(n_3115),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_3084),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3047),
.B(n_273),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3111),
.Y(n_3381)
);

INVx6_ASAP7_75t_L g3382 ( 
.A(n_3108),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3120),
.B(n_275),
.Y(n_3383)
);

OAI22xp5_ASAP7_75t_SL g3384 ( 
.A1(n_3177),
.A2(n_2959),
.B1(n_2885),
.B2(n_2803),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3233),
.Y(n_3385)
);

AOI222xp33_ASAP7_75t_L g3386 ( 
.A1(n_3051),
.A2(n_2265),
.B1(n_2528),
.B2(n_2501),
.C1(n_2868),
.C2(n_2855),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3233),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3249),
.B(n_275),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_SL g3389 ( 
.A1(n_3177),
.A2(n_2864),
.B1(n_2910),
.B2(n_2793),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3099),
.B(n_2911),
.Y(n_3390)
);

HB1xp67_ASAP7_75t_L g3391 ( 
.A(n_3248),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3101),
.B(n_2911),
.Y(n_3392)
);

BUFx4f_ASAP7_75t_SL g3393 ( 
.A(n_2997),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3238),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3141),
.A2(n_2457),
.B1(n_2945),
.B2(n_2888),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3238),
.Y(n_3396)
);

BUFx12f_ASAP7_75t_L g3397 ( 
.A(n_3014),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3252),
.B(n_276),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3147),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_3034),
.A2(n_2457),
.B1(n_2945),
.B2(n_2888),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_3036),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3240),
.Y(n_3402)
);

CKINVDCx14_ASAP7_75t_R g3403 ( 
.A(n_2963),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3210),
.A2(n_2457),
.B1(n_2884),
.B2(n_2277),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_3254),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_3036),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3240),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3104),
.B(n_2793),
.Y(n_3408)
);

BUFx2_ASAP7_75t_L g3409 ( 
.A(n_3139),
.Y(n_3409)
);

AOI22xp33_ASAP7_75t_L g3410 ( 
.A1(n_2986),
.A2(n_3221),
.B1(n_3107),
.B2(n_3043),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_SL g3411 ( 
.A1(n_3153),
.A2(n_2910),
.B1(n_2864),
.B2(n_2856),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_2971),
.A2(n_2910),
.B1(n_2841),
.B2(n_2856),
.Y(n_3412)
);

AOI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3063),
.A2(n_3170),
.B1(n_3161),
.B2(n_3181),
.Y(n_3413)
);

AND2x4_ASAP7_75t_L g3414 ( 
.A(n_2986),
.B(n_2841),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3106),
.B(n_2939),
.Y(n_3415)
);

INVx3_ASAP7_75t_L g3416 ( 
.A(n_3254),
.Y(n_3416)
);

AND2x2_ASAP7_75t_L g3417 ( 
.A(n_3178),
.B(n_3105),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3243),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3157),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3148),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_SL g3421 ( 
.A1(n_3054),
.A2(n_2939),
.B1(n_2884),
.B2(n_2638),
.Y(n_3421)
);

CKINVDCx20_ASAP7_75t_R g3422 ( 
.A(n_2987),
.Y(n_3422)
);

OAI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3235),
.A2(n_2542),
.B1(n_2277),
.B2(n_2317),
.Y(n_3423)
);

OAI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3158),
.A2(n_2304),
.B1(n_2317),
.B2(n_2260),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3174),
.Y(n_3425)
);

INVx1_ASAP7_75t_SL g3426 ( 
.A(n_3196),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3202),
.A2(n_2304),
.B1(n_2391),
.B2(n_2363),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3186),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3243),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3096),
.A2(n_2391),
.B1(n_2408),
.B2(n_2363),
.Y(n_3430)
);

INVx1_ASAP7_75t_SL g3431 ( 
.A(n_3256),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3054),
.A2(n_2391),
.B1(n_2408),
.B2(n_2363),
.Y(n_3432)
);

AOI22xp33_ASAP7_75t_SL g3433 ( 
.A1(n_3187),
.A2(n_2638),
.B1(n_2644),
.B2(n_2622),
.Y(n_3433)
);

OAI21xp5_ASAP7_75t_SL g3434 ( 
.A1(n_3253),
.A2(n_2644),
.B(n_2638),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3114),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3118),
.B(n_3121),
.Y(n_3436)
);

CKINVDCx20_ASAP7_75t_R g3437 ( 
.A(n_3145),
.Y(n_3437)
);

AOI22xp33_ASAP7_75t_SL g3438 ( 
.A1(n_3187),
.A2(n_2657),
.B1(n_2673),
.B2(n_2644),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3245),
.A2(n_2355),
.B1(n_2673),
.B2(n_2657),
.Y(n_3439)
);

CKINVDCx5p33_ASAP7_75t_R g3440 ( 
.A(n_3029),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3122),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3171),
.B(n_277),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3256),
.A2(n_2408),
.B1(n_2454),
.B2(n_2412),
.Y(n_3443)
);

HB1xp67_ASAP7_75t_L g3444 ( 
.A(n_3188),
.Y(n_3444)
);

INVx5_ASAP7_75t_SL g3445 ( 
.A(n_3127),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3191),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3199),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_SL g3448 ( 
.A1(n_3081),
.A2(n_2673),
.B1(n_2705),
.B2(n_2657),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_3123),
.A2(n_2706),
.B1(n_2738),
.B2(n_2705),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_3256),
.A2(n_3246),
.B1(n_3069),
.B2(n_2970),
.Y(n_3450)
);

OAI22xp33_ASAP7_75t_L g3451 ( 
.A1(n_3028),
.A2(n_2124),
.B1(n_2150),
.B2(n_2117),
.Y(n_3451)
);

BUFx12f_ASAP7_75t_L g3452 ( 
.A(n_3165),
.Y(n_3452)
);

CKINVDCx5p33_ASAP7_75t_R g3453 ( 
.A(n_3078),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3149),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3151),
.B(n_2705),
.Y(n_3455)
);

CKINVDCx20_ASAP7_75t_R g3456 ( 
.A(n_3053),
.Y(n_3456)
);

OAI21xp5_ASAP7_75t_SL g3457 ( 
.A1(n_3091),
.A2(n_3057),
.B(n_2988),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_L g3458 ( 
.A1(n_3256),
.A2(n_2454),
.B1(n_2412),
.B2(n_2706),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_3209),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3216),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3207),
.A2(n_3246),
.B1(n_3251),
.B2(n_3239),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3164),
.Y(n_3462)
);

OR2x2_ASAP7_75t_L g3463 ( 
.A(n_3026),
.B(n_2706),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3256),
.A2(n_2454),
.B1(n_2412),
.B2(n_2738),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3168),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3169),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_SL g3467 ( 
.A1(n_3236),
.A2(n_2751),
.B1(n_2755),
.B2(n_2738),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3175),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3180),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3189),
.B(n_2751),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3077),
.B(n_3109),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3258),
.A2(n_2751),
.B1(n_2759),
.B2(n_2755),
.Y(n_3472)
);

OR2x2_ASAP7_75t_L g3473 ( 
.A(n_3032),
.B(n_2755),
.Y(n_3473)
);

AOI22xp33_ASAP7_75t_SL g3474 ( 
.A1(n_3236),
.A2(n_2773),
.B1(n_2776),
.B2(n_2759),
.Y(n_3474)
);

BUFx4f_ASAP7_75t_L g3475 ( 
.A(n_3028),
.Y(n_3475)
);

INVx3_ASAP7_75t_L g3476 ( 
.A(n_3226),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3126),
.B(n_277),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3194),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3066),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3224),
.Y(n_3480)
);

CKINVDCx11_ASAP7_75t_R g3481 ( 
.A(n_2974),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3195),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3208),
.Y(n_3483)
);

OAI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3042),
.A2(n_2124),
.B1(n_2150),
.B2(n_2117),
.Y(n_3484)
);

OAI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3042),
.A2(n_2202),
.B1(n_2773),
.B2(n_2759),
.Y(n_3485)
);

AOI22xp33_ASAP7_75t_L g3486 ( 
.A1(n_3179),
.A2(n_2776),
.B1(n_2785),
.B2(n_2773),
.Y(n_3486)
);

AOI22xp33_ASAP7_75t_L g3487 ( 
.A1(n_3201),
.A2(n_2785),
.B1(n_2800),
.B2(n_2776),
.Y(n_3487)
);

INVx4_ASAP7_75t_L g3488 ( 
.A(n_3218),
.Y(n_3488)
);

AOI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3059),
.A2(n_3048),
.B1(n_3070),
.B2(n_3037),
.Y(n_3489)
);

CKINVDCx5p33_ASAP7_75t_R g3490 ( 
.A(n_3137),
.Y(n_3490)
);

OAI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3075),
.A2(n_2800),
.B1(n_2849),
.B2(n_2785),
.Y(n_3491)
);

BUFx12f_ASAP7_75t_L g3492 ( 
.A(n_3108),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3079),
.A2(n_2849),
.B1(n_2867),
.B2(n_2800),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3260),
.A2(n_3160),
.B1(n_3112),
.B2(n_3198),
.Y(n_3494)
);

AOI22xp33_ASAP7_75t_L g3495 ( 
.A1(n_3304),
.A2(n_3117),
.B1(n_3072),
.B2(n_3062),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3316),
.B(n_3212),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3410),
.A2(n_3072),
.B1(n_3146),
.B2(n_3062),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3304),
.A2(n_3146),
.B1(n_3152),
.B2(n_3213),
.Y(n_3498)
);

OAI22xp5_ASAP7_75t_L g3499 ( 
.A1(n_3307),
.A2(n_3182),
.B1(n_3110),
.B2(n_3205),
.Y(n_3499)
);

OAI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3313),
.A2(n_2983),
.B1(n_3255),
.B2(n_3084),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3273),
.A2(n_3152),
.B1(n_3229),
.B2(n_3215),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3285),
.A2(n_3218),
.B1(n_3162),
.B2(n_3163),
.Y(n_3502)
);

AOI211xp5_ASAP7_75t_SL g3503 ( 
.A1(n_3265),
.A2(n_3056),
.B(n_3200),
.C(n_3257),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3298),
.A2(n_3231),
.B1(n_3128),
.B2(n_3242),
.Y(n_3504)
);

OAI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3306),
.A2(n_3128),
.B1(n_3150),
.B2(n_3203),
.Y(n_3505)
);

OAI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3413),
.A2(n_3204),
.B1(n_3203),
.B2(n_3259),
.Y(n_3506)
);

OAI21xp5_ASAP7_75t_SL g3507 ( 
.A1(n_3457),
.A2(n_3018),
.B(n_2977),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3263),
.B(n_3234),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3378),
.A2(n_3204),
.B1(n_3134),
.B2(n_3183),
.Y(n_3509)
);

AND2x6_ASAP7_75t_L g3510 ( 
.A(n_3431),
.B(n_3039),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_SL g3511 ( 
.A1(n_3268),
.A2(n_3000),
.B1(n_3052),
.B2(n_3157),
.Y(n_3511)
);

OAI22xp5_ASAP7_75t_L g3512 ( 
.A1(n_3284),
.A2(n_3134),
.B1(n_3049),
.B2(n_3214),
.Y(n_3512)
);

AOI22xp5_ASAP7_75t_L g3513 ( 
.A1(n_3282),
.A2(n_3052),
.B1(n_3085),
.B2(n_3225),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3378),
.A2(n_3302),
.B1(n_3293),
.B2(n_3261),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3435),
.Y(n_3515)
);

AOI221xp5_ASAP7_75t_L g3516 ( 
.A1(n_3299),
.A2(n_3119),
.B1(n_3159),
.B2(n_3250),
.C(n_3039),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3289),
.A2(n_3100),
.B1(n_3237),
.B2(n_3136),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3314),
.A2(n_3100),
.B1(n_3136),
.B2(n_3039),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_SL g3519 ( 
.A1(n_3314),
.A2(n_3094),
.B1(n_3087),
.B2(n_3136),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3444),
.B(n_3143),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3270),
.A2(n_3220),
.B1(n_3155),
.B2(n_3166),
.Y(n_3521)
);

AOI22xp33_ASAP7_75t_L g3522 ( 
.A1(n_3270),
.A2(n_3220),
.B1(n_3155),
.B2(n_3166),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3275),
.A2(n_3220),
.B1(n_3155),
.B2(n_3166),
.Y(n_3523)
);

OAI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3457),
.A2(n_3173),
.B1(n_3219),
.B2(n_3143),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_SL g3525 ( 
.A1(n_3315),
.A2(n_3094),
.B1(n_3087),
.B2(n_3143),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3459),
.B(n_3295),
.Y(n_3526)
);

OA222x2_ASAP7_75t_L g3527 ( 
.A1(n_3303),
.A2(n_3219),
.B1(n_3173),
.B2(n_280),
.C1(n_282),
.C2(n_283),
.Y(n_3527)
);

AOI22xp33_ASAP7_75t_L g3528 ( 
.A1(n_3277),
.A2(n_3219),
.B1(n_3173),
.B2(n_2471),
.Y(n_3528)
);

AOI22xp33_ASAP7_75t_SL g3529 ( 
.A1(n_3315),
.A2(n_3277),
.B1(n_3264),
.B2(n_3280),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3274),
.A2(n_2202),
.B1(n_2527),
.B2(n_2849),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3321),
.A2(n_2887),
.B1(n_2907),
.B2(n_2867),
.Y(n_3531)
);

OAI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_3301),
.A2(n_2887),
.B1(n_2907),
.B2(n_2867),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3311),
.A2(n_2907),
.B1(n_2908),
.B2(n_2887),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3266),
.B(n_3426),
.Y(n_3534)
);

AOI22xp33_ASAP7_75t_L g3535 ( 
.A1(n_3333),
.A2(n_2921),
.B1(n_2953),
.B2(n_2908),
.Y(n_3535)
);

OAI22xp5_ASAP7_75t_L g3536 ( 
.A1(n_3330),
.A2(n_2921),
.B1(n_2908),
.B2(n_2953),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3283),
.Y(n_3537)
);

OR2x2_ASAP7_75t_L g3538 ( 
.A(n_3426),
.B(n_278),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3441),
.B(n_278),
.Y(n_3539)
);

INVxp67_ASAP7_75t_L g3540 ( 
.A(n_3336),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3300),
.A2(n_2953),
.B1(n_2921),
.B2(n_2360),
.Y(n_3541)
);

AOI22xp33_ASAP7_75t_L g3542 ( 
.A1(n_3291),
.A2(n_2360),
.B1(n_2349),
.B2(n_283),
.Y(n_3542)
);

AOI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3288),
.A2(n_2360),
.B1(n_284),
.B2(n_279),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3391),
.A2(n_284),
.B1(n_279),
.B2(n_282),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_L g3545 ( 
.A1(n_3386),
.A2(n_3383),
.B1(n_3374),
.B2(n_3364),
.Y(n_3545)
);

AND2x6_ASAP7_75t_L g3546 ( 
.A(n_3431),
.B(n_615),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3454),
.B(n_285),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3386),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3319),
.A2(n_289),
.B1(n_286),
.B2(n_287),
.Y(n_3549)
);

OAI21xp33_ASAP7_75t_L g3550 ( 
.A1(n_3380),
.A2(n_289),
.B(n_290),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3287),
.Y(n_3551)
);

AOI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3329),
.A2(n_294),
.B1(n_291),
.B2(n_292),
.Y(n_3552)
);

AOI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_3281),
.A2(n_295),
.B1(n_291),
.B2(n_292),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3442),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3401),
.A2(n_3406),
.B1(n_3388),
.B2(n_3398),
.Y(n_3555)
);

AOI21x1_ASAP7_75t_L g3556 ( 
.A1(n_3352),
.A2(n_298),
.B(n_299),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3462),
.B(n_300),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3450),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3489),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3356),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3465),
.B(n_307),
.Y(n_3561)
);

OAI221xp5_ASAP7_75t_L g3562 ( 
.A1(n_3361),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.C(n_311),
.Y(n_3562)
);

AOI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3357),
.A2(n_311),
.B1(n_308),
.B2(n_310),
.Y(n_3563)
);

AOI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3269),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3477),
.A2(n_318),
.B1(n_315),
.B2(n_317),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3466),
.B(n_317),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3468),
.B(n_319),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_3360),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3290),
.Y(n_3569)
);

OAI222xp33_ASAP7_75t_L g3570 ( 
.A1(n_3461),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.C1(n_324),
.C2(n_325),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_3269),
.A2(n_326),
.B1(n_322),
.B2(n_324),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3469),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3479),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3461),
.A2(n_331),
.B1(n_327),
.B2(n_329),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3478),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3294),
.B(n_332),
.Y(n_3576)
);

AOI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_3324),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3409),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3482),
.B(n_334),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3267),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3580)
);

OAI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3404),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_3408),
.A2(n_341),
.B1(n_338),
.B2(n_340),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3320),
.B(n_340),
.Y(n_3583)
);

INVxp67_ASAP7_75t_SL g3584 ( 
.A(n_3463),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3332),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_3585)
);

OAI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3305),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_3586)
);

OAI221xp5_ASAP7_75t_L g3587 ( 
.A1(n_3395),
.A2(n_3344),
.B1(n_3343),
.B2(n_3347),
.C(n_3430),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3483),
.B(n_3262),
.Y(n_3588)
);

AOI221xp5_ASAP7_75t_L g3589 ( 
.A1(n_3369),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.C(n_349),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3286),
.B(n_3296),
.Y(n_3590)
);

AOI22xp33_ASAP7_75t_L g3591 ( 
.A1(n_3324),
.A2(n_351),
.B1(n_347),
.B2(n_350),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3322),
.B(n_351),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3337),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_3593)
);

AOI22xp33_ASAP7_75t_L g3594 ( 
.A1(n_3358),
.A2(n_356),
.B1(n_352),
.B2(n_355),
.Y(n_3594)
);

AOI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3355),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3595)
);

OA21x2_ASAP7_75t_L g3596 ( 
.A1(n_3349),
.A2(n_357),
.B(n_358),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3335),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3597)
);

AOI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3334),
.A2(n_366),
.B1(n_362),
.B2(n_365),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3297),
.B(n_367),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3279),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3419),
.A2(n_3414),
.B1(n_3417),
.B2(n_3488),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3345),
.A2(n_371),
.B1(n_368),
.B2(n_370),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3309),
.B(n_371),
.Y(n_3603)
);

OAI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3339),
.A2(n_3445),
.B1(n_3448),
.B2(n_3308),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3317),
.B(n_372),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3331),
.B(n_3353),
.Y(n_3606)
);

NAND3xp33_ASAP7_75t_L g3607 ( 
.A(n_3367),
.B(n_3318),
.C(n_3400),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3414),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3323),
.B(n_373),
.Y(n_3609)
);

AOI22xp33_ASAP7_75t_L g3610 ( 
.A1(n_3488),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3445),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3611)
);

AOI22xp33_ASAP7_75t_L g3612 ( 
.A1(n_3415),
.A2(n_380),
.B1(n_377),
.B2(n_379),
.Y(n_3612)
);

AOI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3280),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3325),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3445),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3336),
.A2(n_387),
.B1(n_384),
.B2(n_385),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3336),
.A2(n_388),
.B1(n_384),
.B2(n_385),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3326),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_SL g3619 ( 
.A1(n_3449),
.A2(n_392),
.B1(n_389),
.B2(n_391),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3365),
.B(n_391),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3359),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3362),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3399),
.B(n_393),
.Y(n_3623)
);

AOI22xp33_ASAP7_75t_L g3624 ( 
.A1(n_3363),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3366),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3376),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3626)
);

OAI22xp5_ASAP7_75t_L g3627 ( 
.A1(n_3308),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_3627)
);

OAI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_3411),
.A2(n_3433),
.B1(n_3438),
.B2(n_3338),
.Y(n_3628)
);

NOR3xp33_ASAP7_75t_L g3629 ( 
.A(n_3272),
.B(n_400),
.C(n_401),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3377),
.B(n_402),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3381),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3385),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3387),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3394),
.A2(n_406),
.B1(n_410),
.B2(n_411),
.Y(n_3634)
);

NAND3xp33_ASAP7_75t_L g3635 ( 
.A(n_3328),
.B(n_410),
.C(n_411),
.Y(n_3635)
);

OAI21xp5_ASAP7_75t_SL g3636 ( 
.A1(n_3434),
.A2(n_412),
.B(n_413),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3396),
.A2(n_412),
.B1(n_415),
.B2(n_416),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3402),
.B(n_416),
.Y(n_3638)
);

OAI21xp33_ASAP7_75t_SL g3639 ( 
.A1(n_3405),
.A2(n_417),
.B(n_419),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3407),
.B(n_417),
.Y(n_3640)
);

OAI21xp33_ASAP7_75t_L g3641 ( 
.A1(n_3434),
.A2(n_420),
.B(n_421),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_SL g3642 ( 
.A1(n_3340),
.A2(n_3303),
.B1(n_3373),
.B2(n_3403),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3418),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3429),
.A2(n_422),
.B1(n_425),
.B2(n_426),
.Y(n_3644)
);

AOI22xp5_ASAP7_75t_L g3645 ( 
.A1(n_3382),
.A2(n_425),
.B1(n_429),
.B2(n_431),
.Y(n_3645)
);

NAND3xp33_ASAP7_75t_L g3646 ( 
.A(n_3354),
.B(n_429),
.C(n_431),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3496),
.B(n_3342),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3534),
.B(n_3436),
.Y(n_3648)
);

NOR2xp33_ASAP7_75t_L g3649 ( 
.A(n_3513),
.B(n_3327),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3515),
.Y(n_3650)
);

OAI211xp5_ASAP7_75t_L g3651 ( 
.A1(n_3507),
.A2(n_3529),
.B(n_3642),
.C(n_3511),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3606),
.B(n_3420),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3584),
.B(n_3471),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3526),
.B(n_3405),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3572),
.B(n_3425),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3575),
.B(n_3428),
.Y(n_3656)
);

NOR2xp33_ASAP7_75t_L g3657 ( 
.A(n_3540),
.B(n_3341),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3508),
.B(n_3446),
.Y(n_3658)
);

AND2x2_ASAP7_75t_SL g3659 ( 
.A(n_3601),
.B(n_3475),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3529),
.A2(n_3421),
.B1(n_3475),
.B2(n_3271),
.Y(n_3660)
);

NAND3xp33_ASAP7_75t_L g3661 ( 
.A(n_3498),
.B(n_3509),
.C(n_3504),
.Y(n_3661)
);

AOI211xp5_ASAP7_75t_L g3662 ( 
.A1(n_3604),
.A2(n_3276),
.B(n_3389),
.C(n_3384),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3578),
.B(n_3447),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3614),
.B(n_3460),
.Y(n_3664)
);

OAI21xp5_ASAP7_75t_SL g3665 ( 
.A1(n_3636),
.A2(n_3375),
.B(n_3278),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3537),
.B(n_3480),
.Y(n_3666)
);

NOR3xp33_ASAP7_75t_SL g3667 ( 
.A(n_3499),
.B(n_3453),
.C(n_3490),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3551),
.B(n_3473),
.Y(n_3668)
);

NAND3xp33_ASAP7_75t_L g3669 ( 
.A(n_3589),
.B(n_3487),
.C(n_3486),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3569),
.B(n_3455),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3622),
.B(n_3292),
.Y(n_3671)
);

OAI221xp5_ASAP7_75t_L g3672 ( 
.A1(n_3514),
.A2(n_3310),
.B1(n_3278),
.B2(n_3382),
.C(n_3379),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3520),
.B(n_3470),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3631),
.B(n_3312),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3588),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3590),
.B(n_3371),
.Y(n_3676)
);

AOI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_3629),
.A2(n_3373),
.B1(n_3423),
.B2(n_3439),
.Y(n_3677)
);

OAI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3545),
.A2(n_3310),
.B1(n_3427),
.B2(n_3467),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3555),
.B(n_3416),
.Y(n_3679)
);

OAI21xp33_ASAP7_75t_L g3680 ( 
.A1(n_3641),
.A2(n_3474),
.B(n_3390),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3523),
.B(n_3501),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3495),
.B(n_3372),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3576),
.B(n_3392),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3583),
.B(n_3416),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3538),
.B(n_3472),
.Y(n_3685)
);

OAI221xp5_ASAP7_75t_SL g3686 ( 
.A1(n_3550),
.A2(n_3476),
.B1(n_3370),
.B2(n_3485),
.C(n_3432),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3517),
.B(n_3493),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_SL g3688 ( 
.A1(n_3503),
.A2(n_3375),
.B(n_3476),
.Y(n_3688)
);

OAI221xp5_ASAP7_75t_L g3689 ( 
.A1(n_3639),
.A2(n_3375),
.B1(n_3368),
.B2(n_3349),
.C(n_3412),
.Y(n_3689)
);

NOR3xp33_ASAP7_75t_L g3690 ( 
.A(n_3635),
.B(n_3351),
.C(n_3424),
.Y(n_3690)
);

NOR3xp33_ASAP7_75t_L g3691 ( 
.A(n_3646),
.B(n_3481),
.C(n_3451),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3525),
.B(n_3491),
.Y(n_3692)
);

OAI221xp5_ASAP7_75t_L g3693 ( 
.A1(n_3619),
.A2(n_3491),
.B1(n_3464),
.B2(n_3458),
.C(n_3443),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3539),
.Y(n_3694)
);

NOR3xp33_ASAP7_75t_L g3695 ( 
.A(n_3500),
.B(n_3571),
.C(n_3570),
.Y(n_3695)
);

OAI21xp5_ASAP7_75t_SL g3696 ( 
.A1(n_3525),
.A2(n_3484),
.B(n_3348),
.Y(n_3696)
);

AOI21xp33_ASAP7_75t_L g3697 ( 
.A1(n_3502),
.A2(n_3492),
.B(n_3397),
.Y(n_3697)
);

NAND3xp33_ASAP7_75t_L g3698 ( 
.A(n_3619),
.B(n_3440),
.C(n_3422),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3535),
.B(n_432),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3527),
.B(n_432),
.Y(n_3700)
);

NOR3xp33_ASAP7_75t_L g3701 ( 
.A(n_3586),
.B(n_433),
.C(n_434),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3570),
.A2(n_3437),
.B(n_3456),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3592),
.B(n_433),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3620),
.B(n_435),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3623),
.B(n_435),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3547),
.B(n_439),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3518),
.B(n_439),
.Y(n_3707)
);

NAND3xp33_ASAP7_75t_L g3708 ( 
.A(n_3516),
.B(n_440),
.C(n_442),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3521),
.B(n_440),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3557),
.B(n_443),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3506),
.A2(n_3452),
.B1(n_3350),
.B2(n_3393),
.Y(n_3711)
);

NAND3xp33_ASAP7_75t_L g3712 ( 
.A(n_3564),
.B(n_444),
.C(n_445),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3561),
.B(n_444),
.Y(n_3713)
);

NAND3xp33_ASAP7_75t_L g3714 ( 
.A(n_3519),
.B(n_445),
.C(n_446),
.Y(n_3714)
);

OAI21xp5_ASAP7_75t_SL g3715 ( 
.A1(n_3519),
.A2(n_3346),
.B(n_446),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3522),
.B(n_447),
.Y(n_3716)
);

OAI221xp5_ASAP7_75t_SL g3717 ( 
.A1(n_3548),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.C(n_450),
.Y(n_3717)
);

AOI221xp5_ASAP7_75t_L g3718 ( 
.A1(n_3611),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.C(n_453),
.Y(n_3718)
);

NAND3xp33_ASAP7_75t_L g3719 ( 
.A(n_3607),
.B(n_451),
.C(n_453),
.Y(n_3719)
);

OAI21xp5_ASAP7_75t_SL g3720 ( 
.A1(n_3524),
.A2(n_454),
.B(n_455),
.Y(n_3720)
);

OAI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3556),
.A2(n_454),
.B(n_456),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3651),
.B(n_3532),
.Y(n_3722)
);

OR2x2_ASAP7_75t_L g3723 ( 
.A(n_3647),
.B(n_3599),
.Y(n_3723)
);

INVxp67_ASAP7_75t_L g3724 ( 
.A(n_3649),
.Y(n_3724)
);

NOR3xp33_ASAP7_75t_L g3725 ( 
.A(n_3651),
.B(n_3615),
.C(n_3505),
.Y(n_3725)
);

INVxp67_ASAP7_75t_L g3726 ( 
.A(n_3653),
.Y(n_3726)
);

AOI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3695),
.A2(n_3494),
.B1(n_3497),
.B2(n_3512),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3654),
.B(n_3541),
.Y(n_3728)
);

AO21x2_ASAP7_75t_L g3729 ( 
.A1(n_3719),
.A2(n_3721),
.B(n_3691),
.Y(n_3729)
);

AO21x2_ASAP7_75t_L g3730 ( 
.A1(n_3691),
.A2(n_3567),
.B(n_3566),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3675),
.B(n_3596),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3663),
.B(n_3533),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3673),
.B(n_3596),
.Y(n_3733)
);

HB1xp67_ASAP7_75t_L g3734 ( 
.A(n_3652),
.Y(n_3734)
);

OR2x2_ASAP7_75t_L g3735 ( 
.A(n_3648),
.B(n_3603),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3650),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3679),
.B(n_3536),
.Y(n_3737)
);

AOI221xp5_ASAP7_75t_L g3738 ( 
.A1(n_3660),
.A2(n_3573),
.B1(n_3560),
.B2(n_3627),
.C(n_3562),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3671),
.B(n_3605),
.Y(n_3739)
);

AO21x2_ASAP7_75t_L g3740 ( 
.A1(n_3690),
.A2(n_3579),
.B(n_3609),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3674),
.B(n_3630),
.Y(n_3741)
);

NOR3xp33_ASAP7_75t_L g3742 ( 
.A(n_3715),
.B(n_3587),
.C(n_3628),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3666),
.B(n_3638),
.Y(n_3743)
);

NAND4xp75_ASAP7_75t_L g3744 ( 
.A(n_3659),
.B(n_3577),
.C(n_3598),
.D(n_3613),
.Y(n_3744)
);

NOR3xp33_ASAP7_75t_L g3745 ( 
.A(n_3697),
.B(n_3602),
.C(n_3581),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3668),
.B(n_3531),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3655),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3670),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3681),
.B(n_3510),
.Y(n_3749)
);

NAND4xp75_ASAP7_75t_L g3750 ( 
.A(n_3700),
.B(n_3702),
.C(n_3667),
.D(n_3692),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3656),
.Y(n_3751)
);

NAND4xp75_ASAP7_75t_L g3752 ( 
.A(n_3687),
.B(n_3595),
.C(n_3645),
.D(n_3553),
.Y(n_3752)
);

NAND3xp33_ASAP7_75t_L g3753 ( 
.A(n_3711),
.B(n_3720),
.C(n_3665),
.Y(n_3753)
);

OR2x2_ASAP7_75t_L g3754 ( 
.A(n_3658),
.B(n_3640),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3685),
.B(n_3510),
.Y(n_3755)
);

NOR3xp33_ASAP7_75t_L g3756 ( 
.A(n_3708),
.B(n_3549),
.C(n_3530),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3657),
.B(n_3510),
.Y(n_3757)
);

OA211x2_ASAP7_75t_L g3758 ( 
.A1(n_3680),
.A2(n_3552),
.B(n_3591),
.C(n_3528),
.Y(n_3758)
);

NAND3xp33_ASAP7_75t_L g3759 ( 
.A(n_3662),
.B(n_3574),
.C(n_3558),
.Y(n_3759)
);

AOI22xp33_ASAP7_75t_L g3760 ( 
.A1(n_3690),
.A2(n_3661),
.B1(n_3701),
.B2(n_3672),
.Y(n_3760)
);

NAND2x1_ASAP7_75t_L g3761 ( 
.A(n_3698),
.B(n_3546),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3676),
.B(n_3510),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3696),
.A2(n_3546),
.B1(n_3600),
.B2(n_3565),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3664),
.Y(n_3764)
);

NOR3xp33_ASAP7_75t_L g3765 ( 
.A(n_3686),
.B(n_3542),
.C(n_3546),
.Y(n_3765)
);

OR2x2_ASAP7_75t_L g3766 ( 
.A(n_3683),
.B(n_3559),
.Y(n_3766)
);

OA21x2_ASAP7_75t_L g3767 ( 
.A1(n_3688),
.A2(n_3563),
.B(n_3585),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3694),
.B(n_3510),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3714),
.A2(n_3546),
.B(n_3543),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3682),
.B(n_3546),
.Y(n_3770)
);

NOR3xp33_ASAP7_75t_L g3771 ( 
.A(n_3686),
.B(n_3610),
.C(n_3544),
.Y(n_3771)
);

BUFx3_ASAP7_75t_L g3772 ( 
.A(n_3684),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3709),
.B(n_3554),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3716),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_L g3775 ( 
.A(n_3672),
.B(n_3582),
.Y(n_3775)
);

AOI22xp5_ASAP7_75t_L g3776 ( 
.A1(n_3678),
.A2(n_3608),
.B1(n_3612),
.B2(n_3568),
.Y(n_3776)
);

HB1xp67_ASAP7_75t_L g3777 ( 
.A(n_3699),
.Y(n_3777)
);

NAND4xp75_ASAP7_75t_L g3778 ( 
.A(n_3707),
.B(n_3593),
.C(n_3597),
.D(n_3580),
.Y(n_3778)
);

INVx2_ASAP7_75t_SL g3779 ( 
.A(n_3703),
.Y(n_3779)
);

XOR2x2_ASAP7_75t_L g3780 ( 
.A(n_3750),
.B(n_3701),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3736),
.Y(n_3781)
);

INVx2_ASAP7_75t_SL g3782 ( 
.A(n_3757),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3734),
.B(n_3748),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3747),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3751),
.B(n_3704),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3731),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3731),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3764),
.Y(n_3788)
);

XOR2x2_ASAP7_75t_L g3789 ( 
.A(n_3742),
.B(n_3689),
.Y(n_3789)
);

NAND3xp33_ASAP7_75t_SL g3790 ( 
.A(n_3760),
.B(n_3689),
.C(n_3718),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3768),
.Y(n_3791)
);

HB1xp67_ASAP7_75t_L g3792 ( 
.A(n_3733),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3761),
.A2(n_3693),
.B(n_3677),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3768),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3743),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3753),
.B(n_3718),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3737),
.B(n_3669),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3777),
.B(n_3706),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3743),
.Y(n_3799)
);

NAND4xp75_ASAP7_75t_SL g3800 ( 
.A(n_3767),
.B(n_3717),
.C(n_3712),
.D(n_3693),
.Y(n_3800)
);

AOI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3725),
.A2(n_3713),
.B1(n_3710),
.B2(n_3705),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3754),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3728),
.B(n_3594),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3739),
.B(n_3618),
.Y(n_3804)
);

NOR4xp25_ASAP7_75t_L g3805 ( 
.A(n_3722),
.B(n_3717),
.C(n_3616),
.D(n_3617),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3726),
.B(n_3621),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3739),
.B(n_3624),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3749),
.B(n_3625),
.Y(n_3808)
);

BUFx3_ASAP7_75t_L g3809 ( 
.A(n_3772),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3735),
.B(n_3626),
.Y(n_3810)
);

INVx1_ASAP7_75t_SL g3811 ( 
.A(n_3732),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3746),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3741),
.Y(n_3813)
);

OAI31xp33_ASAP7_75t_SL g3814 ( 
.A1(n_3753),
.A2(n_3644),
.A3(n_3643),
.B(n_3637),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3741),
.Y(n_3815)
);

INVx3_ASAP7_75t_L g3816 ( 
.A(n_3755),
.Y(n_3816)
);

NAND4xp75_ASAP7_75t_L g3817 ( 
.A(n_3758),
.B(n_3727),
.C(n_3763),
.D(n_3767),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3762),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3723),
.Y(n_3819)
);

XNOR2x2_ASAP7_75t_L g3820 ( 
.A(n_3759),
.B(n_3632),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3774),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3779),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3770),
.B(n_3633),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3766),
.Y(n_3824)
);

NAND4xp75_ASAP7_75t_SL g3825 ( 
.A(n_3775),
.B(n_456),
.C(n_457),
.D(n_458),
.Y(n_3825)
);

NOR2x1_ASAP7_75t_R g3826 ( 
.A(n_3773),
.B(n_457),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3730),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3730),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3740),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3783),
.Y(n_3830)
);

INVxp67_ASAP7_75t_L g3831 ( 
.A(n_3796),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3802),
.Y(n_3832)
);

XOR2x2_ASAP7_75t_L g3833 ( 
.A(n_3789),
.B(n_3759),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3824),
.B(n_3724),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3783),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3786),
.Y(n_3836)
);

XOR2x2_ASAP7_75t_L g3837 ( 
.A(n_3789),
.B(n_3744),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3802),
.Y(n_3838)
);

XOR2x2_ASAP7_75t_L g3839 ( 
.A(n_3817),
.B(n_3752),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3824),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3784),
.Y(n_3841)
);

OAI22x1_ASAP7_75t_SL g3842 ( 
.A1(n_3780),
.A2(n_3729),
.B1(n_3740),
.B2(n_3765),
.Y(n_3842)
);

XNOR2x2_ASAP7_75t_L g3843 ( 
.A(n_3820),
.B(n_3738),
.Y(n_3843)
);

OA22x2_ASAP7_75t_L g3844 ( 
.A1(n_3796),
.A2(n_3776),
.B1(n_3729),
.B2(n_3771),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3788),
.Y(n_3845)
);

XOR2x2_ASAP7_75t_L g3846 ( 
.A(n_3780),
.B(n_3778),
.Y(n_3846)
);

INVx1_ASAP7_75t_SL g3847 ( 
.A(n_3809),
.Y(n_3847)
);

INVx2_ASAP7_75t_SL g3848 ( 
.A(n_3809),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3781),
.Y(n_3849)
);

INVx2_ASAP7_75t_SL g3850 ( 
.A(n_3782),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3786),
.Y(n_3851)
);

NOR2x1_ASAP7_75t_R g3852 ( 
.A(n_3826),
.B(n_3769),
.Y(n_3852)
);

AND2x4_ASAP7_75t_L g3853 ( 
.A(n_3782),
.B(n_3769),
.Y(n_3853)
);

XOR2x2_ASAP7_75t_L g3854 ( 
.A(n_3800),
.B(n_3745),
.Y(n_3854)
);

INVx1_ASAP7_75t_SL g3855 ( 
.A(n_3822),
.Y(n_3855)
);

XOR2x2_ASAP7_75t_L g3856 ( 
.A(n_3820),
.B(n_3756),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3792),
.B(n_3634),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3791),
.B(n_458),
.Y(n_3858)
);

INVxp67_ASAP7_75t_L g3859 ( 
.A(n_3828),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3787),
.Y(n_3860)
);

OAI22xp5_ASAP7_75t_L g3861 ( 
.A1(n_3847),
.A2(n_3793),
.B1(n_3811),
.B2(n_3797),
.Y(n_3861)
);

OR2x2_ASAP7_75t_L g3862 ( 
.A(n_3840),
.B(n_3787),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3834),
.Y(n_3863)
);

OAI22xp5_ASAP7_75t_L g3864 ( 
.A1(n_3847),
.A2(n_3797),
.B1(n_3792),
.B2(n_3816),
.Y(n_3864)
);

HB1xp67_ASAP7_75t_L g3865 ( 
.A(n_3848),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3830),
.Y(n_3866)
);

OAI22x1_ASAP7_75t_L g3867 ( 
.A1(n_3831),
.A2(n_3829),
.B1(n_3827),
.B2(n_3801),
.Y(n_3867)
);

XNOR2x1_ASAP7_75t_SL g3868 ( 
.A(n_3854),
.B(n_3790),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3841),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3845),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3849),
.Y(n_3871)
);

INVx1_ASAP7_75t_SL g3872 ( 
.A(n_3855),
.Y(n_3872)
);

OA22x2_ASAP7_75t_L g3873 ( 
.A1(n_3831),
.A2(n_3827),
.B1(n_3819),
.B2(n_3815),
.Y(n_3873)
);

OA22x2_ASAP7_75t_L g3874 ( 
.A1(n_3853),
.A2(n_3813),
.B1(n_3798),
.B2(n_3816),
.Y(n_3874)
);

XOR2x2_ASAP7_75t_L g3875 ( 
.A(n_3837),
.B(n_3825),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3832),
.Y(n_3876)
);

AOI22x1_ASAP7_75t_L g3877 ( 
.A1(n_3843),
.A2(n_3806),
.B1(n_3821),
.B2(n_3810),
.Y(n_3877)
);

HB1xp67_ASAP7_75t_L g3878 ( 
.A(n_3855),
.Y(n_3878)
);

XOR2x2_ASAP7_75t_L g3879 ( 
.A(n_3846),
.B(n_3839),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3850),
.Y(n_3880)
);

OAI22xp5_ASAP7_75t_L g3881 ( 
.A1(n_3844),
.A2(n_3816),
.B1(n_3812),
.B2(n_3821),
.Y(n_3881)
);

OA22x2_ASAP7_75t_L g3882 ( 
.A1(n_3853),
.A2(n_3795),
.B1(n_3799),
.B2(n_3812),
.Y(n_3882)
);

BUFx3_ASAP7_75t_L g3883 ( 
.A(n_3858),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3838),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3859),
.Y(n_3885)
);

AO22x1_ASAP7_75t_L g3886 ( 
.A1(n_3858),
.A2(n_3806),
.B1(n_3804),
.B2(n_3807),
.Y(n_3886)
);

XNOR2x1_ASAP7_75t_L g3887 ( 
.A(n_3856),
.B(n_3785),
.Y(n_3887)
);

BUFx3_ASAP7_75t_L g3888 ( 
.A(n_3844),
.Y(n_3888)
);

INVx3_ASAP7_75t_L g3889 ( 
.A(n_3830),
.Y(n_3889)
);

NAND3x1_ASAP7_75t_SL g3890 ( 
.A(n_3852),
.B(n_3803),
.C(n_3805),
.Y(n_3890)
);

AO22x2_ASAP7_75t_L g3891 ( 
.A1(n_3859),
.A2(n_3794),
.B1(n_3818),
.B2(n_3823),
.Y(n_3891)
);

HB1xp67_ASAP7_75t_L g3892 ( 
.A(n_3836),
.Y(n_3892)
);

BUFx2_ASAP7_75t_L g3893 ( 
.A(n_3842),
.Y(n_3893)
);

OA22x2_ASAP7_75t_L g3894 ( 
.A1(n_3833),
.A2(n_3803),
.B1(n_3818),
.B2(n_3808),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3889),
.Y(n_3895)
);

INVx1_ASAP7_75t_SL g3896 ( 
.A(n_3865),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3889),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3878),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3862),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3863),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3885),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3869),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3872),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3870),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3876),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3887),
.B(n_3888),
.Y(n_3906)
);

OAI322xp33_ASAP7_75t_L g3907 ( 
.A1(n_3893),
.A2(n_3857),
.A3(n_3835),
.B1(n_3851),
.B2(n_3836),
.C1(n_3860),
.C2(n_3823),
.Y(n_3907)
);

BUFx2_ASAP7_75t_L g3908 ( 
.A(n_3883),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3871),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3866),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3880),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3884),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3892),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3877),
.Y(n_3914)
);

BUFx2_ASAP7_75t_L g3915 ( 
.A(n_3891),
.Y(n_3915)
);

BUFx2_ASAP7_75t_L g3916 ( 
.A(n_3891),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3877),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3861),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3864),
.Y(n_3919)
);

NAND4xp75_ASAP7_75t_L g3920 ( 
.A(n_3906),
.B(n_3868),
.C(n_3890),
.D(n_3879),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3903),
.Y(n_3921)
);

AOI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3906),
.A2(n_3894),
.B1(n_3893),
.B2(n_3886),
.Y(n_3922)
);

AOI22x1_ASAP7_75t_L g3923 ( 
.A1(n_3914),
.A2(n_3867),
.B1(n_3875),
.B2(n_3886),
.Y(n_3923)
);

AO22x1_ASAP7_75t_L g3924 ( 
.A1(n_3917),
.A2(n_3881),
.B1(n_3882),
.B2(n_3873),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3898),
.Y(n_3925)
);

AOI22x1_ASAP7_75t_L g3926 ( 
.A1(n_3918),
.A2(n_3874),
.B1(n_3835),
.B2(n_3851),
.Y(n_3926)
);

OAI322xp33_ASAP7_75t_L g3927 ( 
.A1(n_3919),
.A2(n_3860),
.A3(n_3814),
.B1(n_461),
.B2(n_462),
.C1(n_463),
.C2(n_464),
.Y(n_3927)
);

OA22x2_ASAP7_75t_L g3928 ( 
.A1(n_3896),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_3928)
);

AOI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3911),
.A2(n_459),
.B1(n_462),
.B2(n_463),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3905),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3905),
.Y(n_3931)
);

BUFx2_ASAP7_75t_L g3932 ( 
.A(n_3908),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3915),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3913),
.Y(n_3934)
);

BUFx4_ASAP7_75t_R g3935 ( 
.A(n_3899),
.Y(n_3935)
);

AOI221xp5_ASAP7_75t_L g3936 ( 
.A1(n_3907),
.A2(n_3916),
.B1(n_3901),
.B2(n_3900),
.C(n_3909),
.Y(n_3936)
);

AOI221xp5_ASAP7_75t_L g3937 ( 
.A1(n_3902),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.C(n_472),
.Y(n_3937)
);

AOI22xp5_ASAP7_75t_L g3938 ( 
.A1(n_3899),
.A2(n_469),
.B1(n_470),
.B2(n_472),
.Y(n_3938)
);

INVxp67_ASAP7_75t_SL g3939 ( 
.A(n_3928),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3932),
.Y(n_3940)
);

AO22x2_ASAP7_75t_L g3941 ( 
.A1(n_3920),
.A2(n_3904),
.B1(n_3912),
.B2(n_3910),
.Y(n_3941)
);

OAI211xp5_ASAP7_75t_L g3942 ( 
.A1(n_3922),
.A2(n_3897),
.B(n_3895),
.C(n_3910),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3921),
.Y(n_3943)
);

A2O1A1Ixp33_ASAP7_75t_L g3944 ( 
.A1(n_3936),
.A2(n_3897),
.B(n_3895),
.C(n_475),
.Y(n_3944)
);

INVxp67_ASAP7_75t_L g3945 ( 
.A(n_3933),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3930),
.Y(n_3946)
);

OAI22x1_ASAP7_75t_L g3947 ( 
.A1(n_3923),
.A2(n_473),
.B1(n_474),
.B2(n_475),
.Y(n_3947)
);

HB1xp67_ASAP7_75t_L g3948 ( 
.A(n_3931),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3925),
.Y(n_3949)
);

OAI22x1_ASAP7_75t_L g3950 ( 
.A1(n_3926),
.A2(n_473),
.B1(n_474),
.B2(n_476),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3935),
.Y(n_3951)
);

O2A1O1Ixp33_ASAP7_75t_L g3952 ( 
.A1(n_3927),
.A2(n_476),
.B(n_478),
.C(n_479),
.Y(n_3952)
);

AO22x2_ASAP7_75t_L g3953 ( 
.A1(n_3934),
.A2(n_478),
.B1(n_480),
.B2(n_481),
.Y(n_3953)
);

OAI22x1_ASAP7_75t_L g3954 ( 
.A1(n_3929),
.A2(n_3938),
.B1(n_3924),
.B2(n_3937),
.Y(n_3954)
);

AOI22x1_ASAP7_75t_SL g3955 ( 
.A1(n_3929),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_3955)
);

AOI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3951),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3947),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3940),
.Y(n_3958)
);

OAI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3939),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3944),
.B(n_489),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3953),
.Y(n_3961)
);

O2A1O1Ixp33_ASAP7_75t_L g3962 ( 
.A1(n_3948),
.A2(n_490),
.B(n_492),
.C(n_494),
.Y(n_3962)
);

AOI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3941),
.A2(n_492),
.B1(n_495),
.B2(n_496),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3945),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3950),
.B(n_497),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3953),
.Y(n_3966)
);

AO22x2_ASAP7_75t_L g3967 ( 
.A1(n_3946),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_3967)
);

AOI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3959),
.A2(n_3941),
.B1(n_3954),
.B2(n_3942),
.Y(n_3968)
);

INVxp67_ASAP7_75t_SL g3969 ( 
.A(n_3965),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3958),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3967),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3961),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3964),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3966),
.Y(n_3974)
);

AO22x2_ASAP7_75t_L g3975 ( 
.A1(n_3960),
.A2(n_3943),
.B1(n_3955),
.B2(n_3949),
.Y(n_3975)
);

AOI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3957),
.A2(n_3952),
.B1(n_503),
.B2(n_504),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3969),
.Y(n_3977)
);

HB1xp67_ASAP7_75t_L g3978 ( 
.A(n_3970),
.Y(n_3978)
);

OAI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3968),
.A2(n_3963),
.B1(n_3956),
.B2(n_3962),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3972),
.Y(n_3980)
);

HB1xp67_ASAP7_75t_L g3981 ( 
.A(n_3974),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3980),
.Y(n_3982)
);

INVx1_ASAP7_75t_SL g3983 ( 
.A(n_3978),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3981),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3977),
.B(n_3976),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3979),
.A2(n_3973),
.B1(n_3975),
.B2(n_3971),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3986),
.A2(n_502),
.B1(n_505),
.B2(n_506),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3982),
.Y(n_3988)
);

BUFx2_ASAP7_75t_L g3989 ( 
.A(n_3984),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3983),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3990),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3988),
.Y(n_3992)
);

AOI221xp5_ASAP7_75t_L g3993 ( 
.A1(n_3992),
.A2(n_3987),
.B1(n_3989),
.B2(n_3985),
.C(n_507),
.Y(n_3993)
);

HB1xp67_ASAP7_75t_L g3994 ( 
.A(n_3993),
.Y(n_3994)
);

AO22x2_ASAP7_75t_L g3995 ( 
.A1(n_3994),
.A2(n_3991),
.B1(n_505),
.B2(n_506),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3995),
.Y(n_3996)
);

AOI221xp5_ASAP7_75t_L g3997 ( 
.A1(n_3996),
.A2(n_502),
.B1(n_508),
.B2(n_509),
.C(n_510),
.Y(n_3997)
);

AOI211xp5_ASAP7_75t_L g3998 ( 
.A1(n_3997),
.A2(n_510),
.B(n_511),
.C(n_512),
.Y(n_3998)
);


endmodule