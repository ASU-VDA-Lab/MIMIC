module real_aes_2177_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_0), .B(n_141), .Y(n_164) );
AOI22xp5_ASAP7_75t_SL g117 ( .A1(n_1), .A2(n_118), .B1(n_121), .B2(n_122), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_1), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_2), .A2(n_135), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_3), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_4), .B(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g140 ( .A(n_5), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_6), .B(n_152), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_7), .B(n_176), .Y(n_561) );
INVx1_ASAP7_75t_L g478 ( .A(n_8), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_9), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_10), .Y(n_494) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_11), .B(n_150), .Y(n_252) );
INVx2_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
AOI221x1_ASAP7_75t_L g134 ( .A1(n_13), .A2(n_25), .B1(n_135), .B2(n_141), .C(n_148), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_15), .B(n_141), .Y(n_248) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_16), .A2(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g569 ( .A(n_17), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_18), .B(n_130), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_19), .B(n_152), .Y(n_234) );
AO21x1_ASAP7_75t_L g174 ( .A1(n_20), .A2(n_141), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g113 ( .A(n_21), .Y(n_113) );
INVx1_ASAP7_75t_L g567 ( .A(n_22), .Y(n_567) );
INVx1_ASAP7_75t_SL g532 ( .A(n_23), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_24), .B(n_142), .Y(n_553) );
NAND2x1_ASAP7_75t_L g162 ( .A(n_26), .B(n_152), .Y(n_162) );
AOI33xp33_ASAP7_75t_L g506 ( .A1(n_27), .A2(n_54), .A3(n_460), .B1(n_465), .B2(n_507), .B3(n_508), .Y(n_506) );
NAND2x1_ASAP7_75t_L g208 ( .A(n_28), .B(n_150), .Y(n_208) );
INVx1_ASAP7_75t_L g487 ( .A(n_29), .Y(n_487) );
OR2x2_ASAP7_75t_L g133 ( .A(n_30), .B(n_89), .Y(n_133) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_30), .A2(n_89), .B(n_132), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_31), .B(n_468), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_32), .B(n_150), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_33), .A2(n_94), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_33), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_34), .B(n_152), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_35), .B(n_150), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_36), .A2(n_135), .B(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g136 ( .A(n_37), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g147 ( .A(n_37), .B(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g459 ( .A(n_37), .Y(n_459) );
OR2x6_ASAP7_75t_L g111 ( .A(n_38), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_39), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_40), .A2(n_51), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_40), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_41), .B(n_141), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_42), .B(n_468), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_43), .A2(n_167), .B1(n_176), .B2(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_44), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_45), .B(n_142), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_46), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_47), .B(n_150), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_48), .B(n_246), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_49), .B(n_142), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_50), .A2(n_135), .B(n_207), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_51), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_52), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_53), .B(n_150), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_55), .B(n_142), .Y(n_518) );
INVx1_ASAP7_75t_L g139 ( .A(n_56), .Y(n_139) );
INVx1_ASAP7_75t_L g144 ( .A(n_56), .Y(n_144) );
AND2x2_ASAP7_75t_L g519 ( .A(n_57), .B(n_130), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_58), .A2(n_76), .B1(n_457), .B2(n_468), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_59), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_60), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_61), .B(n_167), .Y(n_496) );
AOI21xp5_ASAP7_75t_SL g456 ( .A1(n_62), .A2(n_457), .B(n_462), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_63), .A2(n_135), .B(n_161), .Y(n_160) );
XNOR2xp5_ASAP7_75t_L g440 ( .A(n_64), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g564 ( .A(n_65), .Y(n_564) );
AO21x1_ASAP7_75t_L g177 ( .A1(n_66), .A2(n_135), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_67), .B(n_141), .Y(n_198) );
INVx1_ASAP7_75t_L g517 ( .A(n_68), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_69), .B(n_141), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_70), .A2(n_457), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g191 ( .A(n_71), .B(n_131), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_72), .A2(n_440), .B1(n_445), .B2(n_772), .Y(n_439) );
INVx1_ASAP7_75t_L g137 ( .A(n_73), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
AND2x2_ASAP7_75t_L g212 ( .A(n_74), .B(n_166), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_75), .B(n_468), .Y(n_509) );
AND2x2_ASAP7_75t_L g534 ( .A(n_77), .B(n_166), .Y(n_534) );
INVx1_ASAP7_75t_L g565 ( .A(n_78), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_79), .A2(n_457), .B(n_531), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_80), .A2(n_457), .B(n_501), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_81), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
AND2x2_ASAP7_75t_L g196 ( .A(n_83), .B(n_166), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_84), .B(n_141), .Y(n_236) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_85), .B(n_166), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_86), .A2(n_457), .B1(n_504), .B2(n_505), .Y(n_503) );
XNOR2xp5_ASAP7_75t_L g441 ( .A(n_87), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g175 ( .A(n_88), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g169 ( .A(n_90), .B(n_166), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_91), .B(n_150), .Y(n_235) );
INVx1_ASAP7_75t_L g463 ( .A(n_92), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_93), .B(n_152), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_94), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_95), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_96), .A2(n_135), .B(n_233), .Y(n_232) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_97), .A2(n_104), .B1(n_433), .B2(n_438), .C1(n_782), .C2(n_787), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g115 ( .A(n_97), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g510 ( .A(n_97), .B(n_166), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_98), .B(n_152), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_99), .A2(n_485), .B(n_486), .C(n_489), .Y(n_484) );
BUFx2_ASAP7_75t_L g437 ( .A(n_100), .Y(n_437) );
BUFx2_ASAP7_75t_SL g791 ( .A(n_100), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_101), .A2(n_135), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_102), .B(n_142), .Y(n_466) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_115), .B(n_430), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g432 ( .A(n_108), .Y(n_432) );
BUFx2_ASAP7_75t_L g793 ( .A(n_108), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OR2x6_ASAP7_75t_SL g767 ( .A(n_109), .B(n_110), .Y(n_767) );
AND2x6_ASAP7_75t_SL g771 ( .A(n_109), .B(n_111), .Y(n_771) );
OR2x2_ASAP7_75t_L g774 ( .A(n_109), .B(n_111), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
XNOR2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVx1_ASAP7_75t_L g121 ( .A(n_118), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_123), .A2(n_446), .B1(n_765), .B2(n_768), .Y(n_445) );
INVx3_ASAP7_75t_L g779 ( .A(n_123), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g123 ( .A(n_124), .B(n_340), .C(n_380), .D(n_409), .Y(n_123) );
NOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_302), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_259), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_192), .B(n_213), .Y(n_126) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_128), .B(n_155), .Y(n_127) );
AND2x4_ASAP7_75t_L g258 ( .A(n_128), .B(n_218), .Y(n_258) );
INVx1_ASAP7_75t_SL g311 ( .A(n_128), .Y(n_311) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_128), .A2(n_347), .B(n_350), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_SL g350 ( .A1(n_128), .A2(n_351), .B(n_352), .C(n_353), .Y(n_350) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_128), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_128), .B(n_352), .Y(n_413) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_129), .Y(n_290) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_130), .A2(n_198), .B(n_199), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_130), .Y(n_211) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_300) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x4_ASAP7_75t_L g176 ( .A(n_132), .B(n_133), .Y(n_176) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
BUFx3_ASAP7_75t_L g471 ( .A(n_136), .Y(n_471) );
AND2x6_ASAP7_75t_L g150 ( .A(n_137), .B(n_143), .Y(n_150) );
INVx2_ASAP7_75t_L g461 ( .A(n_137), .Y(n_461) );
AND2x4_ASAP7_75t_L g457 ( .A(n_138), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g152 ( .A(n_139), .B(n_145), .Y(n_152) );
INVx2_ASAP7_75t_L g465 ( .A(n_139), .Y(n_465) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_140), .Y(n_470) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
INVx1_ASAP7_75t_L g488 ( .A(n_142), .Y(n_488) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx5_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_147), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_153), .Y(n_148) );
INVxp67_ASAP7_75t_L g568 ( .A(n_150), .Y(n_568) );
INVxp67_ASAP7_75t_L g570 ( .A(n_152), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_153), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_153), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_153), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_153), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_153), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_153), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_153), .A2(n_251), .B(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_153), .A2(n_463), .B(n_464), .C(n_466), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_153), .A2(n_464), .B(n_478), .C(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g504 ( .A(n_153), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_153), .A2(n_464), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_153), .A2(n_464), .B(n_532), .C(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_153), .A2(n_553), .B(n_554), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_153), .B(n_176), .Y(n_571) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_170), .Y(n_155) );
AND2x2_ASAP7_75t_L g282 ( .A(n_156), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g363 ( .A(n_156), .B(n_218), .Y(n_363) );
INVx1_ASAP7_75t_L g423 ( .A(n_156), .Y(n_423) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g267 ( .A(n_157), .B(n_183), .Y(n_267) );
AND2x2_ASAP7_75t_L g392 ( .A(n_157), .B(n_184), .Y(n_392) );
AND2x2_ASAP7_75t_L g397 ( .A(n_157), .B(n_357), .Y(n_397) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVxp67_ASAP7_75t_L g273 ( .A(n_158), .Y(n_273) );
BUFx3_ASAP7_75t_L g306 ( .A(n_158), .Y(n_306) );
AND2x2_ASAP7_75t_L g352 ( .A(n_158), .B(n_184), .Y(n_352) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_165), .B(n_169), .Y(n_158) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_159), .A2(n_165), .B(n_169), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B(n_191), .Y(n_184) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_165), .A2(n_185), .B(n_191), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_165), .A2(n_166), .B1(n_484), .B2(n_490), .Y(n_483) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_165), .A2(n_513), .B(n_519), .Y(n_512) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_165), .A2(n_513), .B(n_519), .Y(n_577) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_167), .B(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
AND2x2_ASAP7_75t_L g337 ( .A(n_170), .B(n_215), .Y(n_337) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
AND2x4_ASAP7_75t_L g218 ( .A(n_171), .B(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g329 ( .A(n_171), .B(n_313), .Y(n_329) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_171), .B(n_300), .Y(n_372) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx2_ASAP7_75t_L g308 ( .A(n_172), .Y(n_308) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g269 ( .A(n_173), .Y(n_269) );
OAI21x1_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_177), .B(n_181), .Y(n_173) );
INVx1_ASAP7_75t_L g182 ( .A(n_175), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_176), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g230 ( .A(n_176), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_176), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_176), .A2(n_456), .B(n_467), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_183), .B(n_269), .Y(n_272) );
AND2x2_ASAP7_75t_L g357 ( .A(n_183), .B(n_300), .Y(n_357) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g354 ( .A(n_184), .B(n_216), .Y(n_354) );
AND2x2_ASAP7_75t_L g374 ( .A(n_184), .B(n_300), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_186), .B(n_190), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_192), .B(n_263), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_192), .A2(n_386), .B1(n_387), .B2(n_388), .C(n_390), .Y(n_385) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OAI332xp33_ASAP7_75t_L g419 ( .A1(n_193), .A2(n_279), .A3(n_286), .B1(n_345), .B2(n_420), .B3(n_421), .C1(n_422), .C2(n_424), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
AND2x2_ASAP7_75t_L g224 ( .A(n_194), .B(n_204), .Y(n_224) );
AND2x2_ASAP7_75t_L g241 ( .A(n_194), .B(n_242), .Y(n_241) );
INVx4_ASAP7_75t_L g254 ( .A(n_194), .Y(n_254) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_194), .B(n_255), .Y(n_314) );
INVx5_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_SL g276 ( .A(n_195), .B(n_242), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_195), .B(n_203), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_195), .B(n_204), .Y(n_287) );
BUFx2_ASAP7_75t_L g322 ( .A(n_195), .Y(n_322) );
AND2x2_ASAP7_75t_L g377 ( .A(n_195), .B(n_245), .Y(n_377) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
OR2x2_ASAP7_75t_L g244 ( .A(n_203), .B(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g255 ( .A(n_203), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g295 ( .A(n_203), .Y(n_295) );
AND2x2_ASAP7_75t_L g365 ( .A(n_203), .B(n_264), .Y(n_365) );
AND2x2_ASAP7_75t_L g378 ( .A(n_203), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_203), .B(n_379), .Y(n_396) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_204), .Y(n_262) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_211), .A2(n_528), .B(n_534), .Y(n_527) );
OAI32xp33_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .A3(n_225), .B1(n_239), .B2(n_257), .Y(n_213) );
INVx2_ASAP7_75t_L g323 ( .A(n_214), .Y(n_323) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
INVx1_ASAP7_75t_L g334 ( .A(n_215), .Y(n_334) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x4_ASAP7_75t_L g268 ( .A(n_216), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g401 ( .A(n_216), .B(n_306), .Y(n_401) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g313 ( .A(n_219), .Y(n_313) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
INVx2_ASAP7_75t_L g301 ( .A(n_222), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_222), .B(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_223), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g389 ( .A(n_223), .Y(n_389) );
AND2x2_ASAP7_75t_L g407 ( .A(n_223), .B(n_269), .Y(n_407) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp67_ASAP7_75t_SL g351 ( .A(n_226), .B(n_280), .Y(n_351) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_227), .B(n_262), .Y(n_349) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g425 ( .A(n_228), .B(n_295), .Y(n_425) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
INVx2_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_237), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_230), .B(n_238), .Y(n_237) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_230), .A2(n_231), .B(n_237), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_236), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_253), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_240), .B(n_299), .Y(n_384) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
AND3x2_ASAP7_75t_L g339 ( .A(n_241), .B(n_286), .C(n_295), .Y(n_339) );
AND2x2_ASAP7_75t_L g263 ( .A(n_242), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_242), .B(n_245), .Y(n_320) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g274 ( .A(n_244), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
INVx1_ASAP7_75t_L g279 ( .A(n_245), .Y(n_279) );
BUFx3_ASAP7_75t_L g286 ( .A(n_245), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_245), .B(n_297), .Y(n_296) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_246), .A2(n_476), .B(n_480), .Y(n_475) );
INVx2_ASAP7_75t_SL g501 ( .A(n_246), .Y(n_501) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x4_ASAP7_75t_L g305 ( .A(n_254), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_254), .B(n_264), .Y(n_348) );
AND2x2_ASAP7_75t_L g304 ( .A(n_255), .B(n_279), .Y(n_304) );
INVx2_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AOI211xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_265), .B(n_270), .C(n_291), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_260), .A2(n_387), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_263), .B(n_322), .Y(n_321) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_263), .A2(n_342), .B(n_346), .C(n_355), .Y(n_341) );
AND2x2_ASAP7_75t_L g327 ( .A(n_264), .B(n_287), .Y(n_327) );
OR2x2_ASAP7_75t_L g330 ( .A(n_264), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_267), .B(n_372), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_268), .B(n_313), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_268), .A2(n_294), .B1(n_374), .B2(n_377), .C(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g345 ( .A(n_269), .B(n_300), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_274), .B1(n_277), .B2(n_281), .C(n_284), .Y(n_270) );
AND2x2_ASAP7_75t_L g416 ( .A(n_271), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g283 ( .A(n_272), .Y(n_283) );
INVx1_ASAP7_75t_L g369 ( .A(n_273), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_274), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g288 ( .A(n_276), .B(n_279), .Y(n_288) );
AND2x2_ASAP7_75t_L g364 ( .A(n_276), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g289 ( .A(n_283), .B(n_290), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_289), .Y(n_284) );
INVx1_ASAP7_75t_L g408 ( .A(n_285), .Y(n_408) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g387 ( .A(n_286), .B(n_314), .Y(n_387) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_287), .B(n_296), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_298), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_326), .B1(n_329), .B2(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g398 ( .A(n_292), .Y(n_398) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
INVx1_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_299), .B(n_369), .Y(n_420) );
AND2x2_ASAP7_75t_L g388 ( .A(n_300), .B(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_301), .A2(n_382), .B(n_385), .C(n_393), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_324), .Y(n_302) );
AOI322xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .A3(n_307), .B1(n_309), .B2(n_314), .C1(n_315), .C2(n_323), .Y(n_303) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_305), .Y(n_421) );
AND2x2_ASAP7_75t_L g371 ( .A(n_306), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g405 ( .A(n_306), .Y(n_405) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_SL g356 ( .A(n_308), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_308), .B(n_354), .Y(n_362) );
AND2x2_ASAP7_75t_L g386 ( .A(n_308), .B(n_352), .Y(n_386) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g358 ( .A(n_312), .Y(n_358) );
NAND2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_321), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_SL g361 ( .A1(n_317), .A2(n_362), .B1(n_363), .B2(n_364), .C(n_366), .Y(n_361) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g428 ( .A(n_320), .Y(n_428) );
AOI211xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B(n_328), .C(n_332), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g403 ( .A(n_327), .Y(n_403) );
INVx1_ASAP7_75t_L g335 ( .A(n_329), .Y(n_335) );
OR2x2_ASAP7_75t_L g422 ( .A(n_329), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g418 ( .A(n_330), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .B(n_338), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_334), .B(n_352), .Y(n_429) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_361), .Y(n_340) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_344), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g395 ( .A(n_348), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI21xp33_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_359), .Y(n_355) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AOI31xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .A3(n_373), .B(n_375), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_372), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B1(n_398), .B2(n_399), .C(n_402), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_406), .B2(n_408), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_419), .C(n_426), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g783 ( .A(n_432), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_SL g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx2_ASAP7_75t_L g786 ( .A(n_435), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_435), .A2(n_789), .B(n_792), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_437), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_439), .B(n_775), .Y(n_438) );
INVx1_ASAP7_75t_L g776 ( .A(n_440), .Y(n_776) );
INVx2_ASAP7_75t_L g781 ( .A(n_446), .Y(n_781) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_655), .C(n_720), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_609), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_556), .B(n_582), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_520), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_472), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g656 ( .A1(n_452), .A2(n_657), .B(n_668), .Y(n_656) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_452), .B(n_598), .Y(n_691) );
AND2x2_ASAP7_75t_L g706 ( .A(n_452), .B(n_707), .Y(n_706) );
OR2x6_ASAP7_75t_L g716 ( .A(n_452), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g718 ( .A(n_452), .B(n_708), .Y(n_718) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g592 ( .A(n_453), .Y(n_592) );
AND2x2_ASAP7_75t_L g605 ( .A(n_453), .B(n_606), .Y(n_605) );
INVx4_ASAP7_75t_L g624 ( .A(n_453), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_453), .B(n_545), .Y(n_627) );
NOR2x1_ASAP7_75t_SL g630 ( .A(n_453), .B(n_560), .Y(n_630) );
AND2x4_ASAP7_75t_L g642 ( .A(n_453), .B(n_640), .Y(n_642) );
OR2x2_ASAP7_75t_L g652 ( .A(n_453), .B(n_527), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_453), .B(n_664), .Y(n_669) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVxp67_ASAP7_75t_L g495 ( .A(n_457), .Y(n_495) );
NOR2x1p5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x6_ASAP7_75t_L g464 ( .A(n_461), .B(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g485 ( .A(n_464), .Y(n_485) );
INVx2_ASAP7_75t_L g555 ( .A(n_464), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_464), .A2(n_488), .B1(n_564), .B2(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g469 ( .A(n_465), .B(n_470), .Y(n_469) );
INVxp33_ASAP7_75t_L g507 ( .A(n_465), .Y(n_507) );
INVx1_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_471), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_472), .A2(n_598), .B1(n_693), .B2(n_694), .Y(n_692) );
INVx1_ASAP7_75t_SL g736 ( .A(n_472), .Y(n_736) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_498), .Y(n_472) );
INVx2_ASAP7_75t_L g667 ( .A(n_473), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_473), .B(n_613), .Y(n_739) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_481), .Y(n_473) );
BUFx3_ASAP7_75t_L g585 ( .A(n_474), .Y(n_585) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g578 ( .A(n_475), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_475), .B(n_500), .Y(n_600) );
AND2x4_ASAP7_75t_L g617 ( .A(n_475), .B(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g633 ( .A(n_475), .Y(n_633) );
INVx2_ASAP7_75t_L g690 ( .A(n_475), .Y(n_690) );
AND2x2_ASAP7_75t_L g608 ( .A(n_481), .B(n_574), .Y(n_608) );
NOR2xp67_ASAP7_75t_L g654 ( .A(n_481), .B(n_577), .Y(n_654) );
AND2x2_ASAP7_75t_L g673 ( .A(n_481), .B(n_577), .Y(n_673) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
INVx1_ASAP7_75t_L g616 ( .A(n_482), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_482), .B(n_512), .Y(n_635) );
AND2x4_ASAP7_75t_L g689 ( .A(n_482), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_491), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g648 ( .A(n_498), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_498), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .Y(n_498) );
AND2x2_ASAP7_75t_L g632 ( .A(n_499), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g672 ( .A(n_499), .Y(n_672) );
AND2x2_ASAP7_75t_L g677 ( .A(n_499), .B(n_577), .Y(n_677) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_500), .B(n_512), .Y(n_539) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_510), .Y(n_500) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_501), .A2(n_502), .B(n_510), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_509), .Y(n_502) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g613 ( .A(n_511), .Y(n_613) );
NAND2x1p5_ASAP7_75t_L g731 ( .A(n_511), .B(n_585), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_511), .B(n_537), .Y(n_752) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_512), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI21xp33_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_535), .B(n_540), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_523), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g604 ( .A(n_524), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g638 ( .A(n_524), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g704 ( .A(n_524), .B(n_622), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_524), .B(n_751), .C(n_752), .Y(n_750) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_525), .Y(n_581) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g597 ( .A(n_527), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_527), .B(n_560), .Y(n_603) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_527), .Y(n_614) );
AND2x2_ASAP7_75t_L g659 ( .A(n_527), .B(n_559), .Y(n_659) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_527), .Y(n_682) );
INVx1_ASAP7_75t_L g699 ( .A(n_527), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g741 ( .A(n_535), .Y(n_741) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_536), .B(n_612), .Y(n_713) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g575 ( .A(n_537), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI211x1_ASAP7_75t_L g609 ( .A1(n_541), .A2(n_610), .B(n_619), .C(n_636), .Y(n_609) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_542), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g662 ( .A(n_542), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_559), .Y(n_598) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g558 ( .A(n_545), .B(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
INVx1_ASAP7_75t_L g640 ( .A(n_545), .Y(n_640) );
AND2x2_ASAP7_75t_L g708 ( .A(n_545), .B(n_560), .Y(n_708) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .C(n_550), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_572), .B(n_579), .Y(n_556) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_557), .B(n_624), .Y(n_727) );
INVx2_ASAP7_75t_L g759 ( .A(n_557), .Y(n_759) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g591 ( .A(n_558), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g606 ( .A(n_560), .Y(n_606) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B(n_571), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
OR2x2_ASAP7_75t_L g666 ( .A(n_573), .B(n_667), .Y(n_666) );
NAND2x1_ASAP7_75t_SL g688 ( .A(n_573), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g588 ( .A(n_574), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g618 ( .A(n_574), .Y(n_618) );
INVx1_ASAP7_75t_L g742 ( .A(n_575), .Y(n_742) );
AND2x2_ASAP7_75t_L g607 ( .A(n_576), .B(n_608), .Y(n_607) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g589 ( .A(n_577), .Y(n_589) );
INVxp33_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g646 ( .A(n_581), .B(n_639), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B(n_593), .C(n_601), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g670 ( .A(n_584), .B(n_671), .Y(n_670) );
NOR2xp67_ASAP7_75t_SL g675 ( .A(n_584), .B(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_585), .B(n_672), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
AND2x2_ASAP7_75t_L g719 ( .A(n_588), .B(n_689), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g737 ( .A1(n_591), .A2(n_738), .B1(n_740), .B2(n_743), .C1(n_744), .C2(n_747), .Y(n_737) );
INVx1_ASAP7_75t_L g701 ( .A(n_592), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_599), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_597), .Y(n_628) );
AND2x4_ASAP7_75t_SL g663 ( .A(n_597), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g717 ( .A(n_598), .Y(n_717) );
AND2x2_ASAP7_75t_L g762 ( .A(n_598), .B(n_614), .Y(n_762) );
AND2x2_ASAP7_75t_L g643 ( .A(n_599), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g756 ( .A(n_600), .B(n_635), .Y(n_756) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_604), .B(n_607), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_602), .A2(n_622), .B(n_663), .Y(n_723) );
AND2x2_ASAP7_75t_L g747 ( .A(n_603), .B(n_624), .Y(n_747) );
NOR2xp33_ASAP7_75t_SL g757 ( .A(n_603), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g695 ( .A(n_606), .Y(n_695) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_606), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g730 ( .A(n_608), .Y(n_730) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g733 ( .A(n_613), .B(n_617), .Y(n_733) );
BUFx2_ASAP7_75t_L g621 ( .A(n_614), .Y(n_621) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g644 ( .A(n_616), .Y(n_644) );
INVx2_ASAP7_75t_L g650 ( .A(n_616), .Y(n_650) );
AND2x2_ASAP7_75t_L g686 ( .A(n_616), .B(n_677), .Y(n_686) );
AND2x4_ASAP7_75t_L g653 ( .A(n_617), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g693 ( .A(n_617), .B(n_650), .Y(n_693) );
AND2x2_ASAP7_75t_L g744 ( .A(n_617), .B(n_745), .Y(n_744) );
AOI31xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_625), .A3(n_629), .B(n_631), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g641 ( .A(n_621), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_SL g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x4_ASAP7_75t_L g639 ( .A(n_624), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_627), .A2(n_679), .B1(n_710), .B2(n_713), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_627), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g764 ( .A(n_627), .B(n_680), .Y(n_764) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g679 ( .A(n_630), .B(n_680), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
AND2x2_ASAP7_75t_L g702 ( .A(n_632), .B(n_673), .Y(n_702) );
INVx1_ASAP7_75t_L g712 ( .A(n_634), .Y(n_712) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_645), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g735 ( .A(n_638), .Y(n_735) );
AND2x2_ASAP7_75t_L g743 ( .A(n_639), .B(n_695), .Y(n_743) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_639), .Y(n_749) );
AND2x2_ASAP7_75t_L g694 ( .A(n_642), .B(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B1(n_651), .B2(n_653), .Y(n_645) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_648), .A2(n_667), .B1(n_761), .B2(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g660 ( .A(n_653), .Y(n_660) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_683), .Y(n_655) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_659), .A2(n_662), .B(n_665), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_662), .A2(n_686), .B1(n_687), .B2(n_691), .Y(n_685) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_674), .B2(n_678), .Y(n_668) );
INVx1_ASAP7_75t_L g703 ( .A(n_671), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_684), .B(n_696), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_692), .Y(n_684) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
NAND2xp33_ASAP7_75t_SL g738 ( .A(n_688), .B(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g711 ( .A(n_689), .Y(n_711) );
INVx3_ASAP7_75t_L g725 ( .A(n_693), .Y(n_725) );
INVxp67_ASAP7_75t_L g754 ( .A(n_694), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_697), .B(n_705), .C(n_709), .D(n_714), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g707 ( .A(n_699), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g755 ( .A(n_703), .Y(n_755) );
NAND2xp33_ASAP7_75t_SL g710 ( .A(n_711), .B(n_712), .Y(n_710) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_719), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND3x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_737), .C(n_748), .Y(n_720) );
AOI221x1_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_726), .B2(n_728), .C(n_734), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp33_ASAP7_75t_SL g728 ( .A(n_729), .B(n_732), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_753), .C(n_760), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_753) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_766), .Y(n_780) );
CKINVDCx11_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
CKINVDCx6p67_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g778 ( .A(n_769), .Y(n_778) );
INVx3_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
OAI22x1_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_777) );
BUFx4f_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVxp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
CKINVDCx8_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
endmodule