module fake_jpeg_298_n_64 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_18;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_5),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_0),
.C(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_3),
.C(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_6),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_12),
.B1(n_15),
.B2(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_12),
.B1(n_27),
.B2(n_19),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_26),
.B(n_28),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_31),
.B(n_38),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_13),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_44),
.B1(n_33),
.B2(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_38),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_14),
.B1(n_11),
.B2(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_43),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_39),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_48),
.C(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_44),
.B1(n_41),
.B2(n_35),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_45),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_58),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_57),
.B(n_53),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_14),
.B(n_20),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.A3(n_51),
.B1(n_52),
.B2(n_20),
.C1(n_9),
.C2(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_54),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_59),
.B(n_10),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_9),
.B1(n_18),
.B2(n_20),
.C(n_43),
.Y(n_64)
);


endmodule