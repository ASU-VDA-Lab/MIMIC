module fake_jpeg_1345_n_482 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_482);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_482;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_45),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_55),
.Y(n_125)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_73),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_17),
.Y(n_77)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_89),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_13),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_92),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_22),
.B1(n_21),
.B2(n_41),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_25),
.B1(n_42),
.B2(n_19),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_22),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_103),
.B(n_135),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_20),
.B1(n_38),
.B2(n_21),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_104),
.A2(n_150),
.B1(n_23),
.B2(n_30),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_21),
.B(n_22),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_151),
.B1(n_31),
.B2(n_18),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_27),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_88),
.B(n_18),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_87),
.A2(n_20),
.B1(n_38),
.B2(n_41),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_75),
.A2(n_29),
.B1(n_42),
.B2(n_19),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_156),
.A2(n_159),
.B1(n_162),
.B2(n_167),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_74),
.C(n_71),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_129),
.C(n_97),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_104),
.B1(n_49),
.B2(n_51),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_115),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_160),
.B(n_164),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_166),
.B(n_175),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_123),
.B1(n_148),
.B2(n_136),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_25),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_29),
.A3(n_42),
.B1(n_18),
.B2(n_31),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_19),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_152),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_180),
.A2(n_188),
.B1(n_193),
.B2(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_137),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_185),
.Y(n_201)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_105),
.A2(n_20),
.B1(n_38),
.B2(n_36),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_122),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_36),
.B1(n_26),
.B2(n_23),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_199),
.B(n_31),
.Y(n_215)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_144),
.B(n_134),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_197),
.B(n_157),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_224),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_141),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g251 ( 
.A1(n_211),
.A2(n_205),
.B(n_202),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_161),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_129),
.B1(n_107),
.B2(n_117),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_222),
.B1(n_161),
.B2(n_179),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_117),
.B1(n_107),
.B2(n_30),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_142),
.C(n_98),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_181),
.B1(n_174),
.B2(n_156),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_244),
.B1(n_252),
.B2(n_256),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_164),
.B1(n_162),
.B2(n_185),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_213),
.B(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_159),
.B1(n_175),
.B2(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_249),
.B1(n_253),
.B2(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_167),
.B1(n_121),
.B2(n_132),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_168),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_250),
.Y(n_282)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_258),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_194),
.B1(n_183),
.B2(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_255),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_121),
.B1(n_132),
.B2(n_108),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_211),
.A2(n_191),
.B1(n_198),
.B2(n_193),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_260),
.B(n_216),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_169),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_108),
.B1(n_98),
.B2(n_106),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_201),
.A2(n_111),
.B1(n_106),
.B2(n_112),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_262),
.B1(n_245),
.B2(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_112),
.B1(n_111),
.B2(n_142),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_201),
.B1(n_228),
.B2(n_212),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_267),
.B1(n_274),
.B2(n_283),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_268),
.B(n_269),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_221),
.B1(n_209),
.B2(n_208),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_221),
.B(n_209),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_216),
.B(n_195),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_280),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_208),
.B1(n_210),
.B2(n_227),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_210),
.B1(n_233),
.B2(n_234),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_249),
.B1(n_261),
.B2(n_260),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_219),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_288),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_204),
.B(n_30),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_247),
.C(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_259),
.C(n_239),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_237),
.A2(n_227),
.B1(n_48),
.B2(n_54),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_236),
.A2(n_226),
.B1(n_170),
.B2(n_177),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_287),
.B1(n_257),
.B2(n_244),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_235),
.A2(n_58),
.B1(n_59),
.B2(n_226),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_236),
.B(n_219),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_292),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_242),
.B1(n_256),
.B2(n_245),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_293),
.A2(n_278),
.B1(n_269),
.B2(n_276),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_297),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_288),
.C(n_285),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_277),
.B(n_262),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_258),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_253),
.B(n_252),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_SL g332 ( 
.A(n_301),
.B(n_278),
.C(n_284),
.Y(n_332)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_307),
.B1(n_316),
.B2(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_305),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_308),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_277),
.A2(n_248),
.B1(n_240),
.B2(n_226),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_268),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_311),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_289),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

XOR2x2_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_281),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_319),
.B(n_325),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_336),
.C(n_346),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_322),
.A2(n_334),
.B1(n_323),
.B2(n_339),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_291),
.B1(n_299),
.B2(n_301),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_334),
.B1(n_339),
.B2(n_340),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_281),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_338),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_288),
.C(n_273),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g358 ( 
.A1(n_332),
.A2(n_303),
.B(n_304),
.C(n_315),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_265),
.B1(n_284),
.B2(n_271),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_279),
.C(n_282),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_337),
.A2(n_342),
.B1(n_295),
.B2(n_290),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_282),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_280),
.B1(n_279),
.B2(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_283),
.B1(n_204),
.B2(n_234),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_294),
.A2(n_232),
.B1(n_203),
.B2(n_207),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_203),
.C(n_207),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_348),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_345),
.A2(n_317),
.B(n_292),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_350),
.A2(n_352),
.B(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_343),
.Y(n_351)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_317),
.B(n_300),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_293),
.B(n_297),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_328),
.B(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_354),
.B(n_361),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_337),
.A2(n_293),
.B1(n_313),
.B2(n_306),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_355),
.A2(n_26),
.B1(n_44),
.B2(n_2),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_356),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_302),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_44),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_371),
.B(n_322),
.Y(n_378)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_363),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_368),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_232),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_365),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_214),
.C(n_316),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_370),
.C(n_332),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_367),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_214),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_316),
.C(n_184),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_331),
.A2(n_163),
.B(n_36),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_327),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_338),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_353),
.B(n_358),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_333),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_379),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_362),
.A2(n_329),
.B1(n_318),
.B2(n_340),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_392),
.B1(n_348),
.B2(n_347),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_325),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_326),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

OAI211xp5_ASAP7_75t_L g385 ( 
.A1(n_366),
.A2(n_331),
.B(n_344),
.C(n_342),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_390),
.B1(n_393),
.B2(n_371),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_355),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_344),
.C(n_26),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_388),
.B(n_396),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_369),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_0),
.C(n_1),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_357),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_401),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_370),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_350),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_415),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_391),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_406),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_369),
.C(n_352),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_356),
.C(n_347),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_377),
.B(n_395),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_389),
.B(n_390),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_383),
.A2(n_362),
.B1(n_364),
.B2(n_358),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_358),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_375),
.B(n_12),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_416),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_376),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_413),
.A2(n_379),
.B1(n_389),
.B2(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_420),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_400),
.C(n_410),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_407),
.A2(n_375),
.B(n_386),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_423),
.A2(n_9),
.B(n_1),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_433),
.Y(n_442)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_396),
.C(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_432),
.B(n_435),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_392),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_397),
.C(n_384),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_425),
.A2(n_398),
.B(n_402),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_447),
.B(n_428),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_415),
.C(n_399),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_440),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_431),
.B(n_376),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_441),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_434),
.B(n_409),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_424),
.B(n_404),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_398),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_445),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_422),
.B(n_384),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_416),
.C(n_393),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_449),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_432),
.B(n_9),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_421),
.B(n_428),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_450),
.A2(n_461),
.B(n_419),
.Y(n_463)
);

AOI21xp33_ASAP7_75t_L g469 ( 
.A1(n_452),
.A2(n_453),
.B(n_458),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_443),
.A2(n_418),
.B(n_421),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_454),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_433),
.C(n_419),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_459),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_448),
.B(n_442),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_429),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_429),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_0),
.B(n_3),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_458),
.A2(n_427),
.B(n_1),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_464),
.A2(n_465),
.B(n_467),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_7),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_7),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_451),
.A2(n_0),
.B(n_2),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_468),
.A2(n_0),
.B(n_2),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_466),
.A2(n_461),
.B(n_457),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_SL g477 ( 
.A(n_471),
.B(n_469),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g475 ( 
.A1(n_472),
.A2(n_473),
.B(n_474),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_462),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_470),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_476),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_478)
);

OAI321xp33_ASAP7_75t_L g479 ( 
.A1(n_477),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_475),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_478),
.B(n_479),
.C(n_5),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_480),
.A2(n_5),
.B(n_6),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_6),
.Y(n_482)
);


endmodule