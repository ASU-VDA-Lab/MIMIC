module fake_jpeg_32175_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_53),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_54),
.C(n_55),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_24),
.B1(n_50),
.B2(n_49),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_67),
.B1(n_57),
.B2(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_89),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_116),
.Y(n_132)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_66),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.C(n_71),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_56),
.B1(n_66),
.B2(n_72),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_30),
.B(n_46),
.C(n_44),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_74),
.C(n_59),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_117),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_22),
.B1(n_48),
.B2(n_47),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_56),
.B1(n_94),
.B2(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_126),
.Y(n_146)
);

NOR2x1p5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_84),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_23),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_135),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_137),
.B1(n_7),
.B2(n_9),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_4),
.C(n_5),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_139),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_7),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_25),
.B(n_42),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_123),
.C(n_122),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_148),
.C(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_20),
.C(n_40),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_151),
.B2(n_154),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_10),
.B(n_14),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_163),
.B1(n_152),
.B2(n_146),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_130),
.A3(n_138),
.B1(n_126),
.B2(n_34),
.C1(n_36),
.C2(n_37),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_162),
.A3(n_158),
.B1(n_155),
.B2(n_159),
.C1(n_148),
.C2(n_51),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

OAI31xp33_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_152),
.A3(n_151),
.B(n_153),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_167),
.B(n_159),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_118),
.B1(n_145),
.B2(n_32),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_169),
.C(n_160),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_167),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_15),
.CI(n_16),
.CON(n_173),
.SN(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_38),
.B(n_39),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);


endmodule