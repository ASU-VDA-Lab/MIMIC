module fake_netlist_5_120_n_1924 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1924);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1924;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_92),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_82),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_42),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_41),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_89),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_34),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_58),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_85),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_106),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_55),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_31),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_46),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_59),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_133),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_62),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_102),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_10),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_30),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_75),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_83),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_27),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_56),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_86),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_158),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_119),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_141),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_95),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_72),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_3),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_96),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_19),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_107),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_108),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_17),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_90),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_70),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_25),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_49),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_123),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_127),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_11),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_28),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_64),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_94),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_111),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_121),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_9),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_67),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_30),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_87),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_37),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_113),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_165),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_16),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_56),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_52),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_33),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_63),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_18),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_164),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_57),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_99),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_171),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_29),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_132),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_61),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_118),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_112),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_17),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_16),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_2),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_169),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_59),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_130),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_131),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_148),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_33),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_23),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_74),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_28),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_138),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_4),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_26),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_156),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_7),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_26),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_122),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_32),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_15),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_53),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_88),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_6),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_12),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_97),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_58),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_93),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_21),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_155),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_5),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_172),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_178),
.B(n_190),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_272),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_174),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_175),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_198),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_245),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_183),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_221),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_245),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_189),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_193),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_245),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_197),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_264),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_285),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_199),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_304),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_219),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_221),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_201),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_318),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_320),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_281),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_237),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_178),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_208),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_215),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_190),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_191),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_216),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_191),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_228),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_194),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_232),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_238),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_216),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_239),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_194),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_240),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_195),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_173),
.B(n_0),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_241),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_242),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_249),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_251),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_252),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_227),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_195),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_213),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_277),
.B(n_1),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_213),
.B(n_1),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_256),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_257),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_309),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_281),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_217),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_188),
.B(n_8),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_217),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_223),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_186),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_182),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_223),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_227),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_225),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_225),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_173),
.B(n_8),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_258),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_234),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_342),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_346),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_348),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_347),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_350),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_181),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_388),
.Y(n_434)
);

CKINVDCx8_ASAP7_75t_R g435 ( 
.A(n_369),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_344),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_186),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_357),
.B(n_181),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_351),
.B(n_177),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_359),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_349),
.B(n_352),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_362),
.B(n_274),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_329),
.B(n_274),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_366),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_374),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_381),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_412),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_390),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_363),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_397),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_358),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_184),
.B(n_182),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_360),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_402),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_412),
.A2(n_207),
.B1(n_327),
.B2(n_218),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_364),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_403),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_367),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_370),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_371),
.B(n_231),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_370),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_410),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_394),
.B(n_179),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_405),
.B(n_179),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_425),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_345),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_365),
.Y(n_484)
);

NAND2x1_ASAP7_75t_L g485 ( 
.A(n_419),
.B(n_186),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_368),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_375),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_384),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_375),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_355),
.Y(n_492)
);

BUFx8_ASAP7_75t_L g493 ( 
.A(n_356),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_385),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_376),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_356),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_377),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_444),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_427),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_444),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_434),
.B(n_378),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_388),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_421),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_262),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_273),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_487),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_478),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_463),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_482),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_361),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_489),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_395),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_474),
.B(n_260),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_441),
.B(n_401),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_L g533 ( 
.A1(n_479),
.A2(n_372),
.B1(n_415),
.B2(n_361),
.Y(n_533)
);

AND2x2_ASAP7_75t_SL g534 ( 
.A(n_479),
.B(n_329),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_479),
.B(n_343),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_501),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_436),
.Y(n_538)
);

CKINVDCx8_ASAP7_75t_R g539 ( 
.A(n_455),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_479),
.B(n_186),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_463),
.B(n_184),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_440),
.A2(n_409),
.B1(n_226),
.B2(n_295),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_478),
.B(n_185),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_440),
.B(n_263),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_447),
.B(n_185),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_502),
.B(n_488),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_440),
.B(n_266),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_454),
.B(n_205),
.C(n_187),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_471),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_428),
.B(n_186),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_431),
.B(n_214),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_447),
.B(n_187),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_404),
.Y(n_564)
);

NOR2x1p5_ASAP7_75t_L g565 ( 
.A(n_443),
.B(n_226),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_455),
.A2(n_408),
.B1(n_222),
.B2(n_265),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_463),
.B(n_205),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_440),
.B(n_270),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_450),
.B(n_211),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_440),
.B(n_282),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_429),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_490),
.Y(n_577)
);

INVx4_ASAP7_75t_SL g578 ( 
.A(n_440),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_451),
.B(n_382),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_446),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_440),
.A2(n_299),
.B1(n_295),
.B2(n_235),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_493),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_446),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_457),
.B(n_343),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_472),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_461),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_458),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_440),
.B(n_284),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

OAI221xp5_ASAP7_75t_L g597 ( 
.A1(n_502),
.A2(n_426),
.B1(n_408),
.B2(n_255),
.C(n_331),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_446),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_462),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_465),
.B(n_306),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_502),
.B(n_211),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_502),
.B(n_380),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_452),
.B(n_214),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_453),
.B(n_413),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_462),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_435),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_462),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_484),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_456),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_462),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_488),
.B(n_379),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_176),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_460),
.B(n_214),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_469),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_497),
.A2(n_299),
.B1(n_341),
.B2(n_236),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_473),
.B(n_307),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_488),
.B(n_379),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_497),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_473),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_475),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_468),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_491),
.B(n_386),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_497),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_480),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_486),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_480),
.B(n_312),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_468),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_466),
.B(n_387),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_485),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_470),
.A2(n_321),
.B1(n_333),
.B2(n_338),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_491),
.B(n_387),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_389),
.Y(n_638)
);

NAND3x1_ASAP7_75t_L g639 ( 
.A(n_493),
.B(n_259),
.C(n_255),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_476),
.B(n_180),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_468),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_497),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_485),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_494),
.B(n_212),
.Y(n_645)
);

INVx6_ASAP7_75t_L g646 ( 
.A(n_468),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_468),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_483),
.B(n_300),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_481),
.B(n_192),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_483),
.B(n_212),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_483),
.B(n_220),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_483),
.B(n_220),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_483),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_435),
.B(n_200),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_520),
.A2(n_248),
.B1(n_276),
.B2(n_254),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_516),
.B(n_520),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_516),
.B(n_498),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_520),
.A2(n_340),
.B1(n_336),
.B2(n_314),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_L g659 ( 
.A1(n_549),
.A2(n_323),
.B(n_314),
.C(n_315),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_551),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_498),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_534),
.A2(n_276),
.B1(n_340),
.B2(n_336),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_606),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_518),
.B(n_496),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_517),
.B(n_498),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_515),
.B(n_498),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_507),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_634),
.B(n_493),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_500),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_508),
.B(n_513),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_534),
.A2(n_280),
.B1(n_254),
.B2(n_246),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_535),
.A2(n_243),
.B1(n_317),
.B2(n_246),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_631),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_546),
.A2(n_317),
.B1(n_296),
.B2(n_297),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_498),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_574),
.B(n_498),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_551),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_574),
.B(n_483),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_549),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_546),
.A2(n_297),
.B1(n_243),
.B2(n_280),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_535),
.B(n_494),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_519),
.B(n_296),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_546),
.A2(n_315),
.B1(n_316),
.B2(n_323),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_524),
.B(n_316),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_616),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_527),
.B(n_326),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_528),
.B(n_326),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_616),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_634),
.B(n_188),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_532),
.B(n_494),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_SL g694 ( 
.A1(n_567),
.A2(n_531),
.B1(n_577),
.B2(n_564),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_606),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_537),
.B(n_514),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_514),
.B(n_430),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_560),
.B(n_214),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_546),
.A2(n_214),
.B1(n_302),
.B2(n_229),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_630),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_514),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

CKINVDCx8_ASAP7_75t_R g703 ( 
.A(n_577),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_546),
.A2(n_302),
.B1(n_230),
.B2(n_286),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_535),
.B(n_389),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_609),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_533),
.B(n_188),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_530),
.B(n_430),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_535),
.A2(n_302),
.B1(n_303),
.B2(n_233),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_560),
.A2(n_259),
.B(n_293),
.C(n_292),
.Y(n_710)
);

AO221x1_ASAP7_75t_L g711 ( 
.A1(n_635),
.A2(n_566),
.B1(n_341),
.B2(n_334),
.C(n_331),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_631),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_630),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_560),
.Y(n_714)
);

INVx8_ASAP7_75t_L g715 ( 
.A(n_546),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_538),
.A2(n_541),
.B(n_561),
.C(n_550),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_563),
.B(n_430),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_506),
.B(n_302),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_622),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_635),
.A2(n_605),
.B1(n_645),
.B2(n_572),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_509),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_525),
.B(n_391),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_SL g723 ( 
.A1(n_567),
.A2(n_209),
.B1(n_224),
.B2(n_210),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_506),
.B(n_302),
.Y(n_724)
);

AND3x1_ASAP7_75t_L g725 ( 
.A(n_654),
.B(n_289),
.C(n_293),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_628),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_569),
.B(n_571),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_439),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_617),
.B(n_188),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_590),
.B(n_439),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_510),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_542),
.B(n_202),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_628),
.Y(n_734)
);

NAND2x1_ASAP7_75t_L g735 ( 
.A(n_601),
.B(n_439),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_640),
.B(n_204),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_591),
.B(n_391),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_509),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_649),
.B(n_247),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_512),
.B(n_206),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_593),
.B(n_396),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_586),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_583),
.A2(n_310),
.B1(n_337),
.B2(n_289),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_396),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_522),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_SL g747 ( 
.A(n_512),
.B(n_308),
.C(n_253),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_608),
.B(n_398),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_R g749 ( 
.A(n_539),
.B(n_523),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_636),
.B(n_247),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_544),
.A2(n_511),
.B1(n_594),
.B2(n_575),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_635),
.A2(n_244),
.B1(n_261),
.B2(n_267),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_635),
.A2(n_311),
.B1(n_268),
.B2(n_269),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_605),
.B(n_398),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_619),
.B(n_624),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_605),
.B(n_406),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_557),
.B(n_247),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_525),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_522),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_542),
.A2(n_310),
.B1(n_337),
.B2(n_292),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_625),
.B(n_406),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_637),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_557),
.B(n_247),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_559),
.B(n_250),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_505),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_407),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_637),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_542),
.A2(n_334),
.B1(n_335),
.B2(n_339),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_510),
.B(n_602),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_638),
.B(n_407),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_526),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_621),
.B(n_414),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_559),
.B(n_250),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_565),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_644),
.B(n_68),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_579),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_638),
.B(n_645),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_645),
.B(n_414),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_SL g779 ( 
.A(n_539),
.B(n_319),
.C(n_278),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_536),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_607),
.B(n_250),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_632),
.B(n_416),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_607),
.B(n_250),
.Y(n_783)
);

BUFx12f_ASAP7_75t_L g784 ( 
.A(n_523),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_568),
.A2(n_335),
.B1(n_339),
.B2(n_309),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_568),
.A2(n_309),
.B1(n_271),
.B2(n_301),
.Y(n_786)
);

AND2x6_ASAP7_75t_SL g787 ( 
.A(n_576),
.B(n_416),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_618),
.B(n_417),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_644),
.B(n_417),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_618),
.B(n_275),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_568),
.A2(n_309),
.B1(n_279),
.B2(n_305),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_540),
.B(n_423),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_540),
.B(n_423),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_599),
.B(n_422),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_614),
.B(n_298),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_555),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_572),
.A2(n_322),
.B1(n_288),
.B2(n_330),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_578),
.B(n_422),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_526),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_578),
.B(n_420),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_SL g801 ( 
.A(n_597),
.B(n_325),
.C(n_324),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_582),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_582),
.B(n_603),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_588),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_543),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_543),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_614),
.B(n_523),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_562),
.B(n_584),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_614),
.B(n_294),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_572),
.A2(n_291),
.B1(n_290),
.B2(n_287),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_548),
.A2(n_420),
.B(n_170),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_582),
.B(n_163),
.Y(n_812)
);

BUFx12f_ASAP7_75t_L g813 ( 
.A(n_562),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_592),
.B(n_12),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_545),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_545),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_553),
.A2(n_152),
.B(n_151),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_570),
.B(n_13),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_556),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_611),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_572),
.A2(n_620),
.B1(n_652),
.B2(n_651),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_536),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_556),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_584),
.B(n_578),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_603),
.B(n_136),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_SL g827 ( 
.A(n_747),
.B(n_639),
.C(n_650),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_780),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_673),
.B(n_578),
.Y(n_829)
);

AND3x1_ASAP7_75t_SL g830 ( 
.A(n_787),
.B(n_723),
.C(n_694),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_777),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_SL g832 ( 
.A(n_703),
.B(n_784),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_681),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_SL g834 ( 
.A(n_779),
.B(n_639),
.C(n_613),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_705),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_765),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_660),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_660),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_715),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_687),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_663),
.B(n_572),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_777),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_679),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_687),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_726),
.B(n_595),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_SL g846 ( 
.A(n_707),
.B(n_814),
.C(n_692),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_663),
.B(n_572),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_749),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_679),
.Y(n_849)
);

BUFx4f_ASAP7_75t_L g850 ( 
.A(n_715),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_SL g851 ( 
.A(n_669),
.B(n_653),
.C(n_647),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_726),
.B(n_595),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_633),
.Y(n_854)
);

BUFx8_ASAP7_75t_L g855 ( 
.A(n_813),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_656),
.A2(n_623),
.B1(n_643),
.B2(n_629),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_695),
.B(n_603),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_703),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_700),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_673),
.B(n_596),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_695),
.B(n_734),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_681),
.A2(n_596),
.B1(n_643),
.B2(n_623),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_758),
.B(n_629),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_734),
.B(n_610),
.Y(n_864)
);

CKINVDCx11_ASAP7_75t_R g865 ( 
.A(n_784),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_788),
.B(n_573),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_700),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_690),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_713),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_722),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_762),
.B(n_610),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_762),
.B(n_642),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_713),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_665),
.A2(n_642),
.B1(n_627),
.B2(n_601),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_767),
.B(n_736),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_670),
.B(n_503),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_767),
.B(n_642),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_798),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_681),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_690),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_813),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_780),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_702),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_731),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_702),
.B(n_627),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_SL g886 ( 
.A(n_655),
.B(n_589),
.C(n_573),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_675),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_722),
.B(n_587),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_664),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_719),
.B(n_627),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_691),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_731),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_820),
.B(n_585),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_675),
.B(n_80),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_788),
.B(n_587),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_L g896 ( 
.A(n_673),
.B(n_536),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_691),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_712),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_672),
.A2(n_589),
.B(n_547),
.C(n_552),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_719),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_668),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_547),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_772),
.B(n_782),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_671),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_662),
.A2(n_552),
.B1(n_554),
.B2(n_580),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_720),
.B(n_580),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_672),
.A2(n_683),
.B1(n_769),
.B2(n_701),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_737),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_691),
.B(n_503),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_770),
.B(n_552),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_743),
.Y(n_912)
);

INVx6_ASAP7_75t_L g913 ( 
.A(n_754),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_754),
.B(n_610),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_721),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_721),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_712),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_799),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_743),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_677),
.A2(n_585),
.B(n_598),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_799),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_683),
.A2(n_646),
.B1(n_601),
.B2(n_554),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_770),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_715),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_SL g925 ( 
.A(n_750),
.B(n_14),
.C(n_18),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_739),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_780),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_819),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_795),
.B(n_14),
.C(n_19),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_696),
.A2(n_646),
.B1(n_601),
.B2(n_554),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_798),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_756),
.B(n_580),
.Y(n_932)
);

AND3x1_ASAP7_75t_SL g933 ( 
.A(n_725),
.B(n_20),
.C(n_22),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_655),
.A2(n_558),
.B(n_536),
.C(n_641),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_739),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_809),
.B(n_20),
.C(n_22),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_801),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_819),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_811),
.B(n_714),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_536),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_796),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_714),
.B(n_558),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_714),
.B(n_558),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_796),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_729),
.B(n_23),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_778),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_780),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_808),
.B(n_104),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_740),
.B(n_612),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_778),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_823),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_774),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_823),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_746),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_746),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_780),
.Y(n_956)
);

INVx6_ASAP7_75t_L g957 ( 
.A(n_800),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_807),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_822),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_790),
.B(n_612),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_774),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_757),
.B(n_24),
.C(n_25),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_759),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_759),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_822),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_716),
.B(n_610),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_789),
.B(n_558),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_727),
.B(n_558),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_771),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_822),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_805),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_733),
.B(n_100),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_805),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_733),
.A2(n_751),
.B1(n_800),
.B2(n_657),
.Y(n_974)
);

OR2x2_ASAP7_75t_SL g975 ( 
.A(n_755),
.B(n_24),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_806),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_709),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_806),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_710),
.Y(n_979)
);

CKINVDCx8_ASAP7_75t_R g980 ( 
.A(n_698),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_794),
.B(n_612),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_815),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_815),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_738),
.B(n_29),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_822),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_666),
.B(n_604),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_816),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_816),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_760),
.B(n_604),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_720),
.B(n_604),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_752),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_768),
.B(n_598),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_661),
.B(n_641),
.Y(n_993)
);

CKINVDCx14_ASAP7_75t_R g994 ( 
.A(n_752),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_821),
.B(n_641),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_693),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_824),
.B(n_646),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_697),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_822),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_775),
.B(n_674),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_658),
.B(n_641),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_753),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_753),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_SL g1004 ( 
.A(n_775),
.B(n_641),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_711),
.A2(n_646),
.B1(n_588),
.B2(n_615),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_797),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_678),
.B(n_588),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_742),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_SL g1009 ( 
.A(n_786),
.B(n_32),
.C(n_35),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_680),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_735),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_763),
.B(n_588),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_735),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_SL g1014 ( 
.A(n_791),
.B(n_588),
.Y(n_1014)
);

OA22x2_ASAP7_75t_L g1015 ( 
.A1(n_1006),
.A2(n_711),
.B1(n_797),
.B2(n_810),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_939),
.A2(n_821),
.B(n_667),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_836),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_875),
.A2(n_685),
.B1(n_676),
.B2(n_682),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_870),
.B(n_793),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_903),
.B(n_748),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_901),
.B(n_764),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_SL g1022 ( 
.A1(n_841),
.A2(n_847),
.B(n_959),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_904),
.A2(n_1006),
.B(n_934),
.C(n_1000),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_990),
.B(n_708),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_915),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_SL g1026 ( 
.A(n_887),
.B(n_792),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_908),
.A2(n_785),
.B1(n_699),
.B2(n_804),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_828),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_828),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_862),
.A2(n_825),
.B(n_812),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_828),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_896),
.A2(n_802),
.B(n_803),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_1002),
.A2(n_761),
.B1(n_745),
.B2(n_766),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_934),
.A2(n_688),
.A3(n_684),
.B(n_686),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_828),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_839),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_848),
.B(n_773),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_SL g1038 ( 
.A(n_839),
.B(n_818),
.Y(n_1038)
);

CKINVDCx11_ASAP7_75t_R g1039 ( 
.A(n_865),
.Y(n_1039)
);

O2A1O1Ixp5_ASAP7_75t_L g1040 ( 
.A1(n_876),
.A2(n_783),
.B(n_781),
.C(n_659),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1008),
.B(n_689),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_915),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_858),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_899),
.A2(n_817),
.A3(n_717),
.B(n_728),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_920),
.A2(n_1007),
.B(n_993),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_858),
.B(n_730),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_993),
.A2(n_724),
.B(n_718),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_837),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_939),
.A2(n_724),
.B(n_718),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_835),
.B(n_810),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_864),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_957),
.B(n_698),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_837),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_881),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_990),
.B(n_704),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_925),
.B(n_744),
.C(n_615),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_974),
.A2(n_698),
.B(n_615),
.Y(n_1057)
);

AOI211x1_ASAP7_75t_L g1058 ( 
.A1(n_831),
.A2(n_35),
.B(n_36),
.C(n_38),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_860),
.A2(n_698),
.B(n_615),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_923),
.B(n_698),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_1010),
.A2(n_698),
.B(n_615),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_853),
.B(n_38),
.Y(n_1062)
);

OA21x2_ASAP7_75t_L g1063 ( 
.A1(n_899),
.A2(n_128),
.B(n_126),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_950),
.B(n_39),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_905),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_888),
.B(n_40),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_913),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_995),
.A2(n_117),
.B(n_115),
.Y(n_1069)
);

CKINVDCx9p33_ASAP7_75t_R g1070 ( 
.A(n_937),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_995),
.A2(n_105),
.B(n_98),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_990),
.A2(n_91),
.B1(n_84),
.B2(n_77),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_946),
.B(n_40),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_838),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_979),
.A2(n_41),
.A3(n_46),
.B(n_47),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_996),
.B(n_47),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1004),
.A2(n_69),
.B(n_50),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_842),
.B(n_48),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_967),
.A2(n_50),
.B(n_51),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1009),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_986),
.A2(n_54),
.B(n_60),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_839),
.B(n_60),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_910),
.A2(n_63),
.B(n_64),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_910),
.A2(n_65),
.B(n_66),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_942),
.A2(n_65),
.B(n_66),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_878),
.B(n_931),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_838),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_942),
.A2(n_943),
.B(n_911),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_985),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_985),
.A2(n_960),
.B(n_981),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_882),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_859),
.A2(n_873),
.B(n_869),
.C(n_867),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_872),
.A2(n_877),
.B(n_885),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_913),
.B(n_863),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_855),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_SL g1097 ( 
.A1(n_966),
.A2(n_984),
.B(n_1001),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_861),
.B(n_854),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_998),
.A2(n_991),
.A3(n_1003),
.B(n_1012),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_889),
.B(n_909),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_932),
.A2(n_998),
.B(n_989),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_848),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_890),
.A2(n_968),
.B(n_928),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_843),
.B(n_849),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_977),
.A2(n_846),
.B(n_900),
.C(n_880),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_943),
.A2(n_829),
.B(n_926),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_985),
.A2(n_839),
.B(n_940),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_895),
.B(n_866),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_916),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_866),
.A2(n_895),
.B(n_856),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_926),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_913),
.B(n_977),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_886),
.A2(n_972),
.B(n_930),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_840),
.B(n_844),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_949),
.A2(n_951),
.A3(n_953),
.B(n_918),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_957),
.A2(n_931),
.B1(n_878),
.B2(n_924),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_840),
.B(n_844),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_829),
.A2(n_935),
.B(n_955),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_868),
.A2(n_883),
.B(n_880),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_833),
.B(n_879),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_887),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_868),
.B(n_883),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_874),
.A2(n_852),
.B(n_845),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_963),
.A2(n_982),
.B(n_964),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_845),
.A2(n_852),
.B(n_922),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_957),
.A2(n_826),
.B1(n_850),
.B2(n_924),
.Y(n_1126)
);

AOI211x1_ASAP7_75t_L g1127 ( 
.A1(n_921),
.A2(n_938),
.B(n_857),
.C(n_973),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_985),
.A2(n_826),
.B(n_850),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_963),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_902),
.B(n_893),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_864),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_845),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_826),
.A2(n_850),
.B1(n_891),
.B2(n_897),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_976),
.A2(n_983),
.B(n_982),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_833),
.B(n_897),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_898),
.B(n_917),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_976),
.A2(n_988),
.A3(n_987),
.B(n_971),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_994),
.A2(n_945),
.B(n_1002),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_914),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_959),
.A2(n_965),
.B(n_1014),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_987),
.A2(n_988),
.B(n_970),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_914),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_833),
.A2(n_879),
.B(n_897),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_941),
.B(n_944),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_954),
.A2(n_969),
.A3(n_978),
.B(n_959),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_956),
.A2(n_970),
.B(n_1005),
.Y(n_1146)
);

NAND2x1_ASAP7_75t_L g1147 ( 
.A(n_965),
.B(n_927),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_879),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_956),
.A2(n_970),
.B(n_891),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_994),
.B(n_892),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_891),
.A2(n_1014),
.B(n_907),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_929),
.A2(n_936),
.B(n_962),
.C(n_827),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_907),
.A2(n_906),
.B(n_914),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_907),
.A2(n_1013),
.B(n_966),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_965),
.A2(n_927),
.B(n_947),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_956),
.A2(n_1013),
.B(n_907),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_834),
.B(n_851),
.C(n_912),
.Y(n_1157)
);

OA21x2_ASAP7_75t_L g1158 ( 
.A1(n_966),
.A2(n_864),
.B(n_871),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_882),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_871),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_972),
.A2(n_948),
.B(n_871),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_884),
.B(n_892),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_952),
.B(n_961),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_907),
.A2(n_997),
.B(n_980),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1011),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_907),
.A2(n_997),
.B(n_980),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_919),
.B(n_997),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_898),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_882),
.B(n_947),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_882),
.A2(n_947),
.B(n_999),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1023),
.A2(n_948),
.B(n_997),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1151),
.A2(n_933),
.B(n_975),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1026),
.A2(n_832),
.B1(n_958),
.B2(n_917),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1020),
.B(n_919),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1137),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1090),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1017),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1023),
.A2(n_830),
.A3(n_947),
.B(n_999),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1097),
.A2(n_999),
.B(n_927),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1141),
.A2(n_999),
.B(n_927),
.Y(n_1180)
);

CKINVDCx6p67_ASAP7_75t_R g1181 ( 
.A(n_1102),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1039),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1141),
.A2(n_1011),
.B(n_952),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1105),
.A2(n_1011),
.A3(n_958),
.B(n_961),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1156),
.A2(n_1011),
.B(n_855),
.Y(n_1185)
);

AOI22x1_ASAP7_75t_L g1186 ( 
.A1(n_1032),
.A2(n_894),
.B1(n_855),
.B2(n_865),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1156),
.A2(n_894),
.B(n_1140),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_1091),
.B(n_1108),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1098),
.B(n_1024),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1112),
.B(n_1138),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1137),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1054),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1137),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1137),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_1045),
.B(n_1030),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1167),
.B(n_1164),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1090),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1066),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1152),
.B(n_1021),
.C(n_1157),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1121),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1162),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1114),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1022),
.A2(n_1045),
.B(n_1123),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1079),
.A2(n_1030),
.B(n_1101),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1117),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1095),
.B(n_1041),
.Y(n_1206)
);

BUFx2_ASAP7_75t_R g1207 ( 
.A(n_1121),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1024),
.B(n_1050),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1122),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1160),
.B(n_1051),
.Y(n_1210)
);

CKINVDCx6p67_ASAP7_75t_R g1211 ( 
.A(n_1102),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1021),
.A2(n_1040),
.B(n_1110),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1124),
.A2(n_1134),
.B(n_1061),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1160),
.B(n_1051),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1124),
.A2(n_1134),
.B(n_1061),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1036),
.B(n_1164),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1051),
.B(n_1131),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1025),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1025),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1036),
.A2(n_1090),
.B(n_1128),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1036),
.A2(n_1055),
.B(n_1107),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1048),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1086),
.A2(n_1069),
.B(n_1049),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1027),
.A2(n_1018),
.B(n_1125),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1105),
.A2(n_1033),
.B(n_1153),
.C(n_1154),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1103),
.A2(n_1049),
.B(n_1094),
.Y(n_1227)
);

AND2x6_ASAP7_75t_L g1228 ( 
.A(n_1165),
.B(n_1148),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1149),
.A2(n_1089),
.B(n_1146),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1152),
.A2(n_1076),
.B(n_1055),
.C(n_1077),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1039),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1080),
.A2(n_1067),
.B(n_1062),
.C(n_1093),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1149),
.A2(n_1089),
.B(n_1146),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1042),
.Y(n_1234)
);

CKINVDCx16_ASAP7_75t_R g1235 ( 
.A(n_1043),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1113),
.A2(n_1143),
.B(n_1016),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1096),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1166),
.A2(n_1059),
.B(n_1106),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1112),
.A2(n_1046),
.B1(n_1150),
.B2(n_1168),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1166),
.B(n_1158),
.Y(n_1240)
);

INVx8_ASAP7_75t_L g1241 ( 
.A(n_1052),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1080),
.A2(n_1093),
.B(n_1062),
.C(n_1037),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1042),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1086),
.A2(n_1069),
.B(n_1084),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1126),
.A2(n_1161),
.B(n_1133),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1158),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1038),
.A2(n_1116),
.A3(n_1034),
.B(n_1072),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1015),
.A2(n_1073),
.B1(n_1064),
.B2(n_1078),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1158),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1084),
.A2(n_1085),
.B(n_1047),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1063),
.B(n_1120),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1113),
.A2(n_1016),
.B(n_1119),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1150),
.Y(n_1255)
);

CKINVDCx14_ASAP7_75t_R g1256 ( 
.A(n_1043),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1015),
.A2(n_1060),
.B(n_1087),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1104),
.B(n_1163),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1059),
.A2(n_1106),
.B(n_1118),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1083),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1083),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1087),
.A2(n_1056),
.B1(n_1167),
.B2(n_1161),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1100),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1118),
.A2(n_1047),
.B(n_1085),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1109),
.Y(n_1265)
);

CKINVDCx9p33_ASAP7_75t_R g1266 ( 
.A(n_1070),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1109),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1019),
.B(n_1068),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1170),
.A2(n_1155),
.B(n_1063),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1144),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1052),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1167),
.A2(n_1068),
.B1(n_1131),
.B2(n_1074),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1063),
.A2(n_1094),
.B(n_1103),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1120),
.A2(n_1135),
.B(n_1088),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1081),
.A2(n_1053),
.B(n_1129),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1094),
.A2(n_1103),
.B(n_1135),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1277)
);

AO21x1_ASAP7_75t_L g1278 ( 
.A1(n_1082),
.A2(n_1058),
.B(n_1034),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1111),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1136),
.B(n_1065),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1054),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1071),
.A2(n_1169),
.B(n_1147),
.Y(n_1282)
);

INVx4_ASAP7_75t_SL g1283 ( 
.A(n_1028),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1071),
.A2(n_1111),
.B(n_1129),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1034),
.A2(n_1148),
.B(n_1044),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_SL g1286 ( 
.A(n_1071),
.B(n_1028),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1169),
.A2(n_1082),
.B(n_1165),
.Y(n_1287)
);

AO32x2_ASAP7_75t_L g1288 ( 
.A1(n_1034),
.A2(n_1115),
.A3(n_1099),
.B1(n_1044),
.B2(n_1075),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1052),
.A2(n_1065),
.B1(n_1096),
.B2(n_1031),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1145),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1044),
.A2(n_1145),
.A3(n_1075),
.B(n_1029),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_SL g1295 ( 
.A(n_1028),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1145),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1044),
.A2(n_1145),
.B(n_1031),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1052),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1028),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1031),
.B(n_1035),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1031),
.A2(n_1035),
.B(n_1092),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1035),
.A2(n_1092),
.B(n_1159),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1035),
.B(n_1092),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1159),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1159),
.A2(n_1075),
.B1(n_1006),
.B2(n_1002),
.Y(n_1306)
);

OAI222xp33_ASAP7_75t_L g1307 ( 
.A1(n_1159),
.A2(n_1006),
.B1(n_1002),
.B2(n_707),
.C1(n_977),
.C2(n_655),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1137),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1097),
.A2(n_1141),
.B(n_1156),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1039),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1020),
.B(n_1098),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1020),
.B(n_923),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1112),
.B(n_614),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1023),
.A2(n_1105),
.B(n_934),
.C(n_1080),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1138),
.A2(n_1006),
.B1(n_1002),
.B2(n_1003),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1020),
.B(n_1098),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1036),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1137),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1137),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1023),
.A2(n_1079),
.B(n_1045),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1130),
.A2(n_875),
.B(n_1021),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1130),
.A2(n_875),
.B(n_1021),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1039),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1138),
.A2(n_1006),
.B1(n_1002),
.B2(n_1003),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1137),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_1121),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1137),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1023),
.A2(n_934),
.A3(n_899),
.B(n_1105),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1138),
.A2(n_1006),
.B1(n_1002),
.B2(n_1003),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1311),
.B(n_1316),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1223),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1244),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1312),
.B(n_1206),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1312),
.B(n_1190),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_1182),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1199),
.A2(n_1225),
.B1(n_1172),
.B2(n_1323),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1244),
.Y(n_1338)
);

INVx8_ASAP7_75t_L g1339 ( 
.A(n_1241),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1267),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1241),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1172),
.A2(n_1322),
.B1(n_1212),
.B2(n_1330),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1182),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1258),
.B(n_1174),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1315),
.A2(n_1325),
.B1(n_1208),
.B2(n_1249),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1263),
.B(n_1270),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1239),
.A2(n_1313),
.B1(n_1173),
.B2(n_1235),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1262),
.A2(n_1208),
.B1(n_1226),
.B2(n_1271),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1270),
.B(n_1201),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1189),
.B(n_1201),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1268),
.B(n_1202),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1267),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1218),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1177),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_SL g1356 ( 
.A(n_1232),
.B(n_1243),
.C(n_1230),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1171),
.A2(n_1278),
.B1(n_1306),
.B2(n_1186),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1202),
.B(n_1205),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1218),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1310),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1171),
.A2(n_1278),
.B1(n_1186),
.B2(n_1307),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1280),
.B(n_1192),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1171),
.A2(n_1257),
.B1(n_1188),
.B2(n_1256),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1177),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1219),
.Y(n_1365)
);

CKINVDCx8_ASAP7_75t_R g1366 ( 
.A(n_1200),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1219),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1271),
.A2(n_1272),
.B1(n_1289),
.B2(n_1198),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1205),
.B(n_1209),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1241),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1234),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1291),
.A2(n_1296),
.A3(n_1328),
.B(n_1326),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1209),
.B(n_1222),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1234),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1255),
.B(n_1222),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1260),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1255),
.B(n_1277),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1188),
.A2(n_1255),
.B1(n_1290),
.B2(n_1251),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1261),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1261),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1188),
.A2(n_1290),
.B1(n_1251),
.B2(n_1298),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1271),
.A2(n_1200),
.B1(n_1298),
.B2(n_1211),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1295),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1178),
.B(n_1277),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1175),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1310),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1265),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1217),
.B(n_1242),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1265),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1271),
.A2(n_1241),
.B1(n_1324),
.B2(n_1327),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1221),
.A2(n_1246),
.B(n_1220),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1246),
.A2(n_1187),
.B(n_1271),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1217),
.B(n_1242),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1279),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1242),
.B(n_1321),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1187),
.A2(n_1314),
.B(n_1216),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1194),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1251),
.A2(n_1293),
.B1(n_1292),
.B2(n_1196),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1191),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1291),
.A2(n_1296),
.A3(n_1328),
.B(n_1326),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_R g1403 ( 
.A(n_1285),
.B(n_1320),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1192),
.B(n_1281),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1181),
.A2(n_1211),
.B1(n_1237),
.B2(n_1251),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1191),
.Y(n_1406)
);

AOI222xp33_ASAP7_75t_L g1407 ( 
.A1(n_1324),
.A2(n_1231),
.B1(n_1327),
.B2(n_1281),
.C1(n_1274),
.C2(n_1321),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1321),
.B(n_1178),
.Y(n_1408)
);

NAND2x1_ASAP7_75t_L g1409 ( 
.A(n_1228),
.B(n_1176),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1327),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1196),
.B(n_1283),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1196),
.B(n_1283),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1231),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_R g1415 ( 
.A(n_1285),
.B(n_1320),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_SL g1416 ( 
.A(n_1266),
.B(n_1216),
.C(n_1240),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1181),
.A2(n_1237),
.B1(n_1196),
.B2(n_1228),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1216),
.A2(n_1183),
.B(n_1254),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1317),
.A2(n_1304),
.B1(n_1207),
.B2(n_1236),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1178),
.B(n_1184),
.Y(n_1420)
);

CKINVDCx8_ASAP7_75t_R g1421 ( 
.A(n_1283),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1240),
.A2(n_1253),
.B1(n_1317),
.B2(n_1247),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1299),
.B(n_1305),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1178),
.B(n_1184),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1300),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1301),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1228),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1303),
.Y(n_1428)
);

OR2x6_ASAP7_75t_SL g1429 ( 
.A(n_1299),
.B(n_1305),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1240),
.A2(n_1253),
.B1(n_1250),
.B2(n_1247),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1301),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1193),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1178),
.B(n_1184),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1308),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1176),
.B(n_1197),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1308),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1184),
.B(n_1304),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1247),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1318),
.A2(n_1319),
.B1(n_1250),
.B2(n_1253),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1275),
.A2(n_1320),
.B1(n_1286),
.B2(n_1245),
.C(n_1197),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1236),
.A2(n_1285),
.B1(n_1254),
.B2(n_1203),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1250),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1176),
.A2(n_1197),
.B1(n_1320),
.B2(n_1284),
.Y(n_1443)
);

AOI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1185),
.A2(n_1286),
.B(n_1287),
.C(n_1297),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1302),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1228),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1184),
.B(n_1329),
.Y(n_1447)
);

CKINVDCx14_ASAP7_75t_R g1448 ( 
.A(n_1228),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1183),
.A2(n_1254),
.B(n_1203),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1236),
.A2(n_1285),
.B1(n_1203),
.B2(n_1275),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1309),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1329),
.B(n_1228),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_SL g1454 ( 
.A(n_1248),
.B(n_1329),
.C(n_1185),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1287),
.B(n_1302),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1227),
.B(n_1284),
.Y(n_1456)
);

BUFx2_ASAP7_75t_SL g1457 ( 
.A(n_1275),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1180),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1294),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1329),
.B(n_1294),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1329),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1269),
.A2(n_1213),
.B(n_1215),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1294),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1294),
.B(n_1288),
.Y(n_1465)
);

CKINVDCx14_ASAP7_75t_R g1466 ( 
.A(n_1288),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1245),
.A2(n_1252),
.B1(n_1224),
.B2(n_1204),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1288),
.B(n_1248),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1179),
.Y(n_1469)
);

INVx6_ASAP7_75t_L g1470 ( 
.A(n_1179),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1282),
.B(n_1238),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1393),
.B(n_1238),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1356),
.A2(n_1245),
.B1(n_1204),
.B2(n_1224),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1353),
.B(n_1288),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1337),
.A2(n_1224),
.B1(n_1252),
.B2(n_1276),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1337),
.A2(n_1342),
.B1(n_1347),
.B2(n_1345),
.C(n_1331),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1342),
.A2(n_1252),
.B1(n_1282),
.B2(n_1195),
.Y(n_1477)
);

OAI211xp5_ASAP7_75t_L g1478 ( 
.A1(n_1345),
.A2(n_1195),
.B(n_1227),
.C(n_1252),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1335),
.B(n_1276),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1344),
.A2(n_1273),
.B(n_1229),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1334),
.A2(n_1195),
.B1(n_1248),
.B2(n_1288),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1348),
.A2(n_1195),
.B1(n_1229),
.B2(n_1233),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1407),
.A2(n_1264),
.B1(n_1259),
.B2(n_1248),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1361),
.B(n_1248),
.C(n_1259),
.Y(n_1484)
);

AOI211xp5_ASAP7_75t_L g1485 ( 
.A1(n_1405),
.A2(n_1368),
.B(n_1383),
.C(n_1392),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1361),
.A2(n_1391),
.B1(n_1357),
.B2(n_1351),
.C(n_1363),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1366),
.Y(n_1487)
);

OAI211xp5_ASAP7_75t_L g1488 ( 
.A1(n_1363),
.A2(n_1357),
.B(n_1350),
.C(n_1346),
.Y(n_1488)
);

AO22x1_ASAP7_75t_L g1489 ( 
.A1(n_1362),
.A2(n_1413),
.B1(n_1343),
.B2(n_1387),
.Y(n_1489)
);

OAI211xp5_ASAP7_75t_L g1490 ( 
.A1(n_1391),
.A2(n_1410),
.B(n_1358),
.C(n_1370),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1332),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1374),
.B(n_1349),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1404),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1360),
.B1(n_1378),
.B2(n_1364),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1414),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1355),
.A2(n_1376),
.B1(n_1362),
.B2(n_1419),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1419),
.A2(n_1405),
.B1(n_1462),
.B2(n_1447),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1462),
.A2(n_1425),
.B1(n_1428),
.B2(n_1395),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_L g1499 ( 
.A1(n_1397),
.A2(n_1389),
.B(n_1453),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1336),
.A2(n_1417),
.B1(n_1421),
.B2(n_1371),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1448),
.A2(n_1429),
.B1(n_1400),
.B2(n_1379),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1341),
.A2(n_1371),
.B1(n_1339),
.B2(n_1384),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1448),
.A2(n_1400),
.B1(n_1379),
.B2(n_1382),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1466),
.A2(n_1339),
.B1(n_1404),
.B2(n_1333),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1466),
.A2(n_1339),
.B1(n_1420),
.B2(n_1411),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1454),
.A2(n_1398),
.B1(n_1382),
.B2(n_1439),
.C(n_1433),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1338),
.A2(n_1340),
.B1(n_1352),
.B2(n_1341),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1416),
.A2(n_1384),
.B1(n_1411),
.B2(n_1412),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1412),
.A2(n_1414),
.B1(n_1437),
.B2(n_1427),
.Y(n_1509)
);

AO31x2_ASAP7_75t_L g1510 ( 
.A1(n_1443),
.A2(n_1449),
.A3(n_1451),
.B(n_1452),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1385),
.B(n_1408),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1439),
.A2(n_1424),
.B1(n_1461),
.B2(n_1464),
.C(n_1459),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1414),
.A2(n_1469),
.B1(n_1446),
.B2(n_1427),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1446),
.A2(n_1460),
.B1(n_1409),
.B2(n_1435),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1435),
.A2(n_1354),
.B1(n_1359),
.B2(n_1365),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1367),
.A2(n_1372),
.B1(n_1390),
.B2(n_1375),
.Y(n_1516)
);

AOI222xp33_ASAP7_75t_L g1517 ( 
.A1(n_1377),
.A2(n_1380),
.B1(n_1381),
.B2(n_1388),
.C1(n_1468),
.C2(n_1423),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1394),
.A2(n_1396),
.B1(n_1438),
.B2(n_1442),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1426),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1456),
.A2(n_1418),
.B(n_1440),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1438),
.A2(n_1442),
.B1(n_1406),
.B2(n_1401),
.Y(n_1521)
);

BUFx4f_ASAP7_75t_SL g1522 ( 
.A(n_1431),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1436),
.A2(n_1434),
.B1(n_1386),
.B2(n_1432),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1470),
.B2(n_1455),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1444),
.A2(n_1441),
.B(n_1450),
.C(n_1455),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1450),
.A2(n_1441),
.B(n_1467),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1470),
.A2(n_1426),
.B1(n_1386),
.B2(n_1432),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1465),
.B(n_1434),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1470),
.A2(n_1457),
.B1(n_1426),
.B2(n_1445),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1436),
.B(n_1373),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1373),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1458),
.A2(n_1403),
.B1(n_1415),
.B2(n_1373),
.C1(n_1402),
.C2(n_1471),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1463),
.A2(n_1471),
.B1(n_1403),
.B2(n_1415),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1402),
.Y(n_1534)
);

AOI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1463),
.A2(n_1286),
.B(n_1284),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1402),
.B(n_1344),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1402),
.A2(n_1002),
.B1(n_1356),
.B2(n_1199),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_SL g1538 ( 
.A(n_1360),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1356),
.A2(n_1002),
.B1(n_1199),
.B2(n_994),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1540)
);

AOI33xp33_ASAP7_75t_L g1541 ( 
.A1(n_1337),
.A2(n_533),
.A3(n_1325),
.B1(n_1330),
.B2(n_1315),
.B3(n_566),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1335),
.B(n_1307),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1331),
.A2(n_1126),
.B(n_1311),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1546)
);

OAI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1337),
.A2(n_707),
.B(n_655),
.C(n_1342),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1404),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1347),
.A2(n_670),
.B1(n_776),
.B2(n_564),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1399),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1348),
.A2(n_994),
.B1(n_1002),
.B2(n_1190),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1552)
);

NAND4xp25_ASAP7_75t_L g1553 ( 
.A(n_1335),
.B(n_1199),
.C(n_814),
.D(n_670),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1344),
.B(n_1334),
.Y(n_1554)
);

OAI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1337),
.A2(n_1342),
.B1(n_1002),
.B2(n_1006),
.C1(n_994),
.C2(n_1345),
.Y(n_1555)
);

OAI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1337),
.A2(n_670),
.B1(n_665),
.B2(n_531),
.C(n_529),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1407),
.A2(n_776),
.B(n_1325),
.C(n_1315),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1356),
.A2(n_1002),
.B1(n_1199),
.B2(n_994),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1407),
.A2(n_776),
.B(n_1325),
.C(n_1315),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1563)
);

AOI222xp33_ASAP7_75t_L g1564 ( 
.A1(n_1356),
.A2(n_1307),
.B1(n_707),
.B2(n_533),
.C1(n_467),
.C2(n_1009),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1356),
.A2(n_1002),
.B1(n_1199),
.B2(n_994),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1346),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1356),
.A2(n_533),
.B1(n_1307),
.B2(n_725),
.C(n_1337),
.Y(n_1567)
);

BUFx8_ASAP7_75t_SL g1568 ( 
.A(n_1343),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1337),
.A2(n_1315),
.B1(n_1330),
.B2(n_1325),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1347),
.A2(n_1006),
.B1(n_1002),
.B2(n_977),
.Y(n_1570)
);

AOI222xp33_ASAP7_75t_L g1571 ( 
.A1(n_1356),
.A2(n_1307),
.B1(n_707),
.B2(n_533),
.C1(n_467),
.C2(n_1009),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1531),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1534),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1479),
.B(n_1520),
.Y(n_1575)
);

OAI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1556),
.A2(n_1567),
.B(n_1564),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1540),
.A2(n_1542),
.B1(n_1569),
.B2(n_1546),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1544),
.A2(n_1563),
.B1(n_1571),
.B2(n_1476),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1479),
.B(n_1474),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1508),
.Y(n_1581)
);

NOR2xp67_ASAP7_75t_L g1582 ( 
.A(n_1484),
.B(n_1519),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1533),
.B(n_1532),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1533),
.B(n_1473),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1475),
.B(n_1510),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1543),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1545),
.B(n_1490),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1524),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1520),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1543),
.B(n_1555),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1566),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1568),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1510),
.B(n_1525),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1472),
.Y(n_1596)
);

OAI222xp33_ASAP7_75t_L g1597 ( 
.A1(n_1537),
.A2(n_1551),
.B1(n_1560),
.B2(n_1565),
.C1(n_1539),
.C2(n_1486),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1526),
.B(n_1477),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1472),
.B(n_1506),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1536),
.B(n_1481),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1550),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1519),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1539),
.A2(n_1565),
.B1(n_1560),
.B2(n_1559),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1483),
.B(n_1482),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1549),
.B(n_1485),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1535),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1491),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1480),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1512),
.B(n_1497),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1504),
.B(n_1503),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1541),
.B(n_1547),
.C(n_1537),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1504),
.B(n_1499),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1561),
.A2(n_1570),
.B1(n_1554),
.B2(n_1498),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1527),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1478),
.B(n_1523),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1517),
.B(n_1492),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1488),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1529),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1507),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1596),
.Y(n_1621)
);

AO21x1_ASAP7_75t_SL g1622 ( 
.A1(n_1616),
.A2(n_1496),
.B(n_1498),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1573),
.Y(n_1623)
);

NAND2x1_ASAP7_75t_SL g1624 ( 
.A(n_1595),
.B(n_1562),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1501),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1586),
.B(n_1493),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1595),
.B(n_1521),
.Y(n_1628)
);

OAI31xp33_ASAP7_75t_L g1629 ( 
.A1(n_1576),
.A2(n_1500),
.A3(n_1496),
.B(n_1513),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1591),
.B(n_1507),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1576),
.A2(n_1494),
.B1(n_1509),
.B2(n_1538),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1576),
.A2(n_1494),
.B1(n_1548),
.B2(n_1502),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1557),
.B1(n_1552),
.B2(n_1558),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1514),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1518),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1605),
.A2(n_1515),
.B1(n_1487),
.B2(n_1495),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1612),
.A2(n_1577),
.B1(n_1578),
.B2(n_1590),
.Y(n_1637)
);

OAI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1578),
.A2(n_1495),
.B1(n_1518),
.B2(n_1489),
.C(n_1516),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1601),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1607),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1592),
.Y(n_1641)
);

AND2x6_ASAP7_75t_SL g1642 ( 
.A(n_1586),
.B(n_1590),
.Y(n_1642)
);

AO21x2_ASAP7_75t_L g1643 ( 
.A1(n_1606),
.A2(n_1582),
.B(n_1598),
.Y(n_1643)
);

AOI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1597),
.A2(n_1612),
.B(n_1609),
.C(n_1598),
.Y(n_1644)
);

O2A1O1Ixp5_ASAP7_75t_L g1645 ( 
.A1(n_1597),
.A2(n_1609),
.B(n_1598),
.C(n_1604),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1577),
.A2(n_1609),
.B1(n_1603),
.B2(n_1588),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1585),
.B(n_1579),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1592),
.B(n_1617),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1609),
.A2(n_1603),
.B1(n_1588),
.B2(n_1610),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1574),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1574),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1607),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1575),
.B(n_1579),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_SL g1656 ( 
.A1(n_1610),
.A2(n_1588),
.B1(n_1611),
.B2(n_1583),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_R g1657 ( 
.A(n_1593),
.B(n_1583),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1572),
.Y(n_1658)
);

CKINVDCx12_ASAP7_75t_R g1659 ( 
.A(n_1593),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1585),
.B(n_1579),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1585),
.B(n_1579),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1614),
.B(n_1587),
.C(n_1598),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1591),
.B(n_1594),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1623),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1644),
.A2(n_1610),
.B1(n_1614),
.B2(n_1611),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1658),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1648),
.B(n_1596),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1647),
.B(n_1594),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1660),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1647),
.B(n_1594),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1658),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1655),
.B(n_1575),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

INVx3_ASAP7_75t_SL g1676 ( 
.A(n_1618),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1660),
.B(n_1661),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1663),
.B(n_1591),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1661),
.B(n_1585),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1661),
.B(n_1599),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1654),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1663),
.B(n_1599),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1655),
.B(n_1575),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_R g1685 ( 
.A(n_1649),
.B(n_1583),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1654),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1620),
.B(n_1575),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1652),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1599),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1662),
.A2(n_1588),
.B1(n_1587),
.B2(n_1610),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1643),
.B(n_1599),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1620),
.B(n_1608),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1584),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1648),
.B(n_1584),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.B(n_1589),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1630),
.B(n_1580),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1630),
.B(n_1580),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1665),
.A2(n_1644),
.B(n_1645),
.Y(n_1705)
);

NAND2x1p5_ASAP7_75t_L g1706 ( 
.A(n_1673),
.B(n_1596),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1665),
.A2(n_1645),
.B(n_1636),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1703),
.B(n_1704),
.Y(n_1709)
);

AND2x4_ASAP7_75t_SL g1710 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1671),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1703),
.B(n_1634),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1681),
.B(n_1619),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1619),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1704),
.B(n_1634),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1692),
.B(n_1641),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1680),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1682),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1637),
.C(n_1662),
.Y(n_1722)
);

AOI32xp33_ASAP7_75t_L g1723 ( 
.A1(n_1693),
.A2(n_1656),
.A3(n_1636),
.B1(n_1650),
.B2(n_1646),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1692),
.B(n_1641),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1686),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1667),
.B(n_1651),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1676),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1687),
.B(n_1639),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1687),
.B(n_1625),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1683),
.B(n_1618),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1686),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1681),
.B(n_1635),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1683),
.B(n_1625),
.Y(n_1736)
);

INVx3_ASAP7_75t_SL g1737 ( 
.A(n_1676),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1683),
.B(n_1628),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1666),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1699),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1688),
.Y(n_1742)
);

INVx5_ASAP7_75t_L g1743 ( 
.A(n_1673),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1742),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1742),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1713),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1737),
.B(n_1669),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1731),
.B(n_1674),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1715),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1722),
.B(n_1642),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_SL g1751 ( 
.A(n_1737),
.B(n_1685),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1710),
.B(n_1669),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1734),
.B(n_1705),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1731),
.B(n_1674),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1738),
.B(n_1684),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1738),
.B(n_1684),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1710),
.B(n_1669),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1705),
.A2(n_1629),
.B(n_1587),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1717),
.Y(n_1759)
);

OR2x6_ASAP7_75t_L g1760 ( 
.A(n_1707),
.B(n_1667),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1711),
.B(n_1693),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1735),
.B(n_1694),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1734),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1720),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1721),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1723),
.B(n_1656),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1724),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1728),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1743),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1732),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1725),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1707),
.B(n_1673),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1739),
.A2(n_1694),
.B1(n_1691),
.B2(n_1689),
.C(n_1627),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1743),
.B(n_1702),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_1657),
.C(n_1629),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1727),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1729),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1733),
.B(n_1677),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1727),
.B(n_1668),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1741),
.B(n_1730),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1750),
.A2(n_1706),
.B(n_1689),
.Y(n_1787)
);

AND2x4_ASAP7_75t_SL g1788 ( 
.A(n_1782),
.B(n_1740),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1771),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1712),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1746),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1706),
.B(n_1689),
.Y(n_1792)
);

AOI211xp5_ASAP7_75t_L g1793 ( 
.A1(n_1753),
.A2(n_1691),
.B(n_1694),
.C(n_1638),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1775),
.A2(n_1583),
.B1(n_1691),
.B2(n_1604),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1779),
.B(n_1718),
.Y(n_1795)
);

O2A1O1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1767),
.A2(n_1631),
.B(n_1638),
.C(n_1699),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1770),
.B(n_1695),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1773),
.B(n_1695),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1746),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1773),
.B(n_1709),
.Y(n_1800)
);

OAI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1781),
.A2(n_1633),
.B(n_1632),
.C(n_1743),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1781),
.B(n_1702),
.Y(n_1802)
);

XNOR2xp5_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1633),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1749),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

AOI222xp33_ASAP7_75t_L g1806 ( 
.A1(n_1777),
.A2(n_1611),
.B1(n_1604),
.B2(n_1613),
.C1(n_1628),
.C2(n_1635),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1759),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1773),
.B(n_1729),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1759),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1765),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1752),
.B(n_1668),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1744),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1760),
.A2(n_1604),
.B(n_1611),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1760),
.A2(n_1581),
.B1(n_1678),
.B2(n_1658),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1765),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1744),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1771),
.B(n_1572),
.Y(n_1817)
);

AOI21xp33_ASAP7_75t_L g1818 ( 
.A1(n_1760),
.A2(n_1617),
.B(n_1666),
.Y(n_1818)
);

AOI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1760),
.A2(n_1697),
.B(n_1701),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1747),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1752),
.B(n_1668),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1744),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

AOI32xp33_ASAP7_75t_L g1824 ( 
.A1(n_1793),
.A2(n_1747),
.A3(n_1780),
.B1(n_1757),
.B2(n_1761),
.Y(n_1824)
);

OAI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1801),
.A2(n_1780),
.A3(n_1782),
.B(n_1774),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1822),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1802),
.A2(n_1760),
.B1(n_1780),
.B2(n_1757),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1788),
.B(n_1782),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1788),
.B(n_1782),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1812),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

OAI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1794),
.A2(n_1802),
.B1(n_1813),
.B2(n_1818),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1803),
.A2(n_1774),
.B1(n_1780),
.B2(n_1779),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1812),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1820),
.Y(n_1835)
);

OAI21xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1792),
.A2(n_1785),
.B(n_1778),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1817),
.A2(n_1774),
.B(n_1783),
.Y(n_1837)
);

AOI211xp5_ASAP7_75t_L g1838 ( 
.A1(n_1796),
.A2(n_1762),
.B(n_1761),
.C(n_1783),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1800),
.B(n_1795),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1789),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1789),
.B(n_1817),
.Y(n_1841)
);

OAI321xp33_ASAP7_75t_L g1842 ( 
.A1(n_1787),
.A2(n_1762),
.A3(n_1779),
.B1(n_1786),
.B2(n_1763),
.C(n_1745),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1817),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1816),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1797),
.A2(n_1785),
.B1(n_1678),
.B2(n_1756),
.Y(n_1845)
);

NAND4xp75_ASAP7_75t_L g1846 ( 
.A(n_1816),
.B(n_1745),
.C(n_1763),
.D(n_1786),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1791),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1799),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1831),
.B(n_1789),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1839),
.B(n_1835),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1851)
);

XNOR2xp5_ASAP7_75t_L g1852 ( 
.A(n_1833),
.B(n_1790),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1840),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1831),
.B(n_1806),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1841),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1840),
.B(n_1804),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1832),
.B(n_1659),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1823),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1832),
.B(n_1795),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1825),
.A2(n_1842),
.B(n_1837),
.C(n_1843),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1828),
.B(n_1811),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1824),
.A2(n_1798),
.B(n_1808),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1826),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1830),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1841),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_R g1867 ( 
.A(n_1847),
.B(n_1572),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1838),
.B(n_1805),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1853),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1849),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1851),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1855),
.B(n_1866),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1861),
.B(n_1828),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1850),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1855),
.B(n_1848),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1864),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1851),
.B(n_1829),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1866),
.B(n_1846),
.Y(n_1878)
);

NOR3x1_ASAP7_75t_L g1879 ( 
.A(n_1854),
.B(n_1814),
.C(n_1834),
.Y(n_1879)
);

AND3x1_ASAP7_75t_L g1880 ( 
.A(n_1857),
.B(n_1827),
.C(n_1829),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1874),
.A2(n_1859),
.B1(n_1857),
.B2(n_1852),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1880),
.A2(n_1860),
.B1(n_1859),
.B2(n_1868),
.C(n_1862),
.Y(n_1882)
);

OAI211xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1878),
.A2(n_1856),
.B(n_1863),
.C(n_1858),
.Y(n_1883)
);

NAND3xp33_ASAP7_75t_L g1884 ( 
.A(n_1870),
.B(n_1865),
.C(n_1844),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1876),
.A2(n_1867),
.B1(n_1845),
.B2(n_1836),
.C(n_1810),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1869),
.A2(n_1815),
.B(n_1807),
.C(n_1809),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1871),
.B(n_1867),
.Y(n_1887)
);

OAI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1871),
.A2(n_1819),
.B1(n_1745),
.B2(n_1754),
.C(n_1748),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1869),
.A2(n_1766),
.B1(n_1768),
.B2(n_1772),
.C(n_1821),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1872),
.A2(n_1748),
.B1(n_1754),
.B2(n_1756),
.C(n_1755),
.Y(n_1890)
);

AOI322xp5_ASAP7_75t_L g1891 ( 
.A1(n_1875),
.A2(n_1821),
.A3(n_1778),
.B1(n_1776),
.B2(n_1679),
.C1(n_1784),
.C2(n_1672),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1882),
.A2(n_1873),
.B1(n_1877),
.B2(n_1879),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1884),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1887),
.Y(n_1894)
);

INVx5_ASAP7_75t_SL g1895 ( 
.A(n_1883),
.Y(n_1895)
);

AND2x2_ASAP7_75t_SL g1896 ( 
.A(n_1881),
.B(n_1877),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1885),
.B(n_1873),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1888),
.A2(n_1769),
.B(n_1768),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1892),
.A2(n_1886),
.B(n_1889),
.C(n_1891),
.Y(n_1899)
);

OA22x2_ASAP7_75t_L g1900 ( 
.A1(n_1893),
.A2(n_1897),
.B1(n_1894),
.B2(n_1895),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1896),
.A2(n_1890),
.B1(n_1772),
.B2(n_1766),
.Y(n_1901)
);

NOR2x1p5_ASAP7_75t_L g1902 ( 
.A(n_1895),
.B(n_1572),
.Y(n_1902)
);

CKINVDCx16_ASAP7_75t_R g1903 ( 
.A(n_1898),
.Y(n_1903)
);

BUFx12f_ASAP7_75t_L g1904 ( 
.A(n_1896),
.Y(n_1904)
);

AND2x2_ASAP7_75t_SL g1905 ( 
.A(n_1896),
.B(n_1755),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1769),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1904),
.A2(n_1899),
.B1(n_1900),
.B2(n_1902),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1903),
.A2(n_1769),
.B1(n_1666),
.B2(n_1702),
.Y(n_1908)
);

AND3x4_ASAP7_75t_L g1909 ( 
.A(n_1901),
.B(n_1581),
.C(n_1702),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_SL g1910 ( 
.A(n_1901),
.B(n_1776),
.C(n_1784),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1906),
.Y(n_1911)
);

AND2x2_ASAP7_75t_SL g1912 ( 
.A(n_1907),
.B(n_1702),
.Y(n_1912)
);

OR3x2_ASAP7_75t_L g1913 ( 
.A(n_1909),
.B(n_1616),
.C(n_1622),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1911),
.B(n_1908),
.Y(n_1914)
);

AOI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1912),
.B1(n_1913),
.B2(n_1910),
.Y(n_1915)
);

OAI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1581),
.B1(n_1621),
.B2(n_1624),
.C(n_1698),
.Y(n_1916)
);

XNOR2xp5_ASAP7_75t_L g1917 ( 
.A(n_1915),
.B(n_1581),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1698),
.B(n_1695),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1916),
.Y(n_1919)
);

AO221x1_ASAP7_75t_L g1920 ( 
.A1(n_1919),
.A2(n_1602),
.B1(n_1621),
.B2(n_1664),
.C(n_1675),
.Y(n_1920)
);

AO221x1_ASAP7_75t_L g1921 ( 
.A1(n_1918),
.A2(n_1602),
.B1(n_1675),
.B2(n_1664),
.C(n_1701),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1920),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1921),
.B1(n_1698),
.B2(n_1700),
.C(n_1679),
.Y(n_1923)
);

AOI211xp5_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1700),
.B(n_1615),
.C(n_1582),
.Y(n_1924)
);


endmodule