module fake_jpeg_22993_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

O2A1O1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_16),
.A2(n_24),
.B(n_13),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_9),
.B1(n_8),
.B2(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_9),
.B1(n_24),
.B2(n_7),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_21),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_30),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_31),
.C(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_33),
.B1(n_27),
.B2(n_15),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_31),
.C(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_20),
.B1(n_29),
.B2(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_40),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_6),
.C(n_5),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_5),
.C(n_15),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.C(n_46),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_45),
.Y(n_52)
);


endmodule