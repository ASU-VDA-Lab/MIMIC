module fake_aes_11541_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
OAI221xp5_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_3), .Y(n_5) );
CKINVDCx20_ASAP7_75t_R g6 ( .A(n_4), .Y(n_6) );
AOI221xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_6), .Y(n_7) );
AOI22xp33_ASAP7_75t_SL g8 ( .A1(n_7), .A2(n_5), .B1(n_1), .B2(n_2), .Y(n_8) );
NAND3xp33_ASAP7_75t_SL g9 ( .A(n_8), .B(n_0), .C(n_1), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_9), .Y(n_10) );
OAI222xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .B1(n_2), .B2(n_6), .C1(n_8), .C2(n_5), .Y(n_11) );
endmodule