module fake_ariane_3213_n_994 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_994);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_994;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_726;
wire n_479;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_731;
wire n_665;
wire n_336;
wire n_779;
wire n_754;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_705;
wire n_630;
wire n_616;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_69),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_35),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_25),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_1),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_46),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_60),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_1),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_49),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_72),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_98),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_24),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_157),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_102),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_11),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_154),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_168),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_134),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_176),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_40),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_172),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_188),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_148),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_109),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_13),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_160),
.Y(n_253)
);

INVxp33_ASAP7_75t_R g254 ( 
.A(n_67),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_115),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_7),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_144),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_123),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_79),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_151),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_146),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_185),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_177),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_87),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_0),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_224),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_205),
.B(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_203),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_198),
.B(n_2),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

XNOR2x2_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_3),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_200),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_5),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_213),
.B(n_6),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_6),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_214),
.B(n_7),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_215),
.B(n_8),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_200),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_201),
.B(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_216),
.B(n_9),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_9),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_201),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_223),
.B(n_10),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_201),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_212),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_201),
.B(n_10),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_195),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_196),
.B(n_11),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_229),
.B(n_12),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_230),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_12),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_13),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_228),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_245),
.B(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_212),
.B(n_14),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_15),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_202),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_221),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g328 ( 
.A(n_210),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_259),
.B(n_15),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_250),
.B1(n_232),
.B2(n_237),
.Y(n_330)
);

CKINVDCx8_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_243),
.B1(n_226),
.B2(n_225),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_285),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_283),
.A2(n_219),
.B1(n_251),
.B2(n_231),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_238),
.Y(n_335)
);

AO22x2_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_220),
.B1(n_259),
.B2(n_270),
.Y(n_336)
);

OR2x6_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_246),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_287),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_261),
.B1(n_273),
.B2(n_272),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_328),
.A2(n_274),
.B1(n_271),
.B2(n_268),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_197),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_267),
.B1(n_266),
.B2(n_264),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_L g348 ( 
.A1(n_290),
.A2(n_263),
.B1(n_262),
.B2(n_260),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_286),
.A2(n_255),
.B1(n_253),
.B2(n_252),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_286),
.A2(n_249),
.B1(n_248),
.B2(n_247),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_204),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_206),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_280),
.A2(n_244),
.B1(n_242),
.B2(n_240),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_284),
.A2(n_239),
.B1(n_235),
.B2(n_234),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_298),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_298),
.A2(n_222),
.B1(n_218),
.B2(n_217),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_298),
.A2(n_211),
.B1(n_208),
.B2(n_207),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_L g360 ( 
.A1(n_292),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_305),
.A2(n_199),
.B1(n_20),
.B2(n_21),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_199),
.B1(n_20),
.B2(n_21),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g363 ( 
.A1(n_282),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_329),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_199),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_278),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_199),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_278),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_322),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_296),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_199),
.B1(n_32),
.B2(n_33),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_318),
.A2(n_199),
.B1(n_33),
.B2(n_34),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_313),
.B(n_199),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_319),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_31),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_42),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_296),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_279),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_302),
.A2(n_315),
.B1(n_324),
.B2(n_320),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_279),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_300),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_303),
.B(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_375),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_333),
.B(n_311),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_331),
.B(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_313),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_302),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_345),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_357),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_351),
.B(n_320),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_335),
.B(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

AND2x2_ASAP7_75t_SL g429 ( 
.A(n_378),
.B(n_302),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_358),
.B(n_317),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_351),
.B(n_315),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_363),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_358),
.B(n_302),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_359),
.B(n_323),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_355),
.B(n_312),
.Y(n_450)
);

XNOR2x2_ASAP7_75t_L g451 ( 
.A(n_332),
.B(n_293),
.Y(n_451)
);

BUFx5_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_334),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_354),
.B(n_310),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_341),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_340),
.B(n_314),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_339),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_348),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_398),
.B(n_324),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_310),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_310),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_421),
.B(n_337),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_394),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_402),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_429),
.B(n_314),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_337),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_407),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_301),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_413),
.B(n_327),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_413),
.B(n_327),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_419),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_327),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_301),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_307),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_409),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_415),
.B(n_398),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_390),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_307),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_326),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_418),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_397),
.B(n_327),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_411),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_326),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_454),
.B(n_326),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_397),
.B(n_327),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_442),
.B(n_327),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_310),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_437),
.B(n_326),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_408),
.B(n_457),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_326),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_388),
.A2(n_450),
.B(n_389),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_424),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_426),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_449),
.Y(n_512)
);

AND2x2_ASAP7_75t_SL g513 ( 
.A(n_439),
.B(n_281),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_310),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_441),
.B(n_281),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_291),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_396),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_403),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_36),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_438),
.B(n_310),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_431),
.B(n_291),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_432),
.B(n_433),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_434),
.B(n_37),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_446),
.B(n_38),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

BUFx8_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_456),
.B(n_281),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_458),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_39),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_400),
.B(n_281),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_387),
.B(n_39),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_404),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_452),
.B(n_281),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_451),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_288),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_428),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_488),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_488),
.B(n_395),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_504),
.B(n_452),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_493),
.B(n_451),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_535),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_455),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_502),
.B(n_407),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_478),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_452),
.Y(n_554)
);

CKINVDCx8_ASAP7_75t_R g555 ( 
.A(n_474),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_452),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_531),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_43),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_469),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_521),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_469),
.B(n_452),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_288),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_521),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

NAND2x1p5_ASAP7_75t_L g573 ( 
.A(n_467),
.B(n_277),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_498),
.B(n_452),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_467),
.B(n_464),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_498),
.B(n_306),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_541),
.B(n_288),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_512),
.B(n_47),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_489),
.B(n_288),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_489),
.B(n_288),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_306),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_512),
.B(n_306),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_481),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_472),
.B(n_277),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_535),
.B(n_519),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

BUFx8_ASAP7_75t_L g589 ( 
.A(n_473),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_475),
.B(n_289),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_473),
.B(n_306),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_525),
.B(n_470),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_485),
.B(n_277),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_472),
.B(n_289),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_472),
.B(n_277),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_466),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_289),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_527),
.B(n_306),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_490),
.B(n_289),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_475),
.B(n_289),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_295),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_518),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_535),
.B(n_277),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_470),
.B(n_277),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_295),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_516),
.Y(n_609)
);

BUFx4f_ASAP7_75t_SL g610 ( 
.A(n_548),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_552),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_550),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_557),
.B(n_519),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_550),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_596),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_589),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_586),
.A2(n_534),
.B1(n_483),
.B2(n_484),
.Y(n_618)
);

CKINVDCx11_ASAP7_75t_R g619 ( 
.A(n_555),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_552),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_609),
.B(n_527),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_553),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_596),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_605),
.Y(n_624)
);

INVx5_ASAP7_75t_SL g625 ( 
.A(n_586),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_562),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_596),
.Y(n_627)
);

BUFx2_ASAP7_75t_SL g628 ( 
.A(n_559),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_560),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_556),
.Y(n_632)
);

INVx3_ASAP7_75t_SL g633 ( 
.A(n_559),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_584),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_606),
.A2(n_549),
.B1(n_558),
.B2(n_531),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_545),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_561),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_561),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_568),
.B(n_467),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_563),
.Y(n_643)
);

BUFx8_ASAP7_75t_SL g644 ( 
.A(n_593),
.Y(n_644)
);

INVx3_ASAP7_75t_SL g645 ( 
.A(n_569),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_563),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_589),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_566),
.Y(n_650)
);

INVx3_ASAP7_75t_SL g651 ( 
.A(n_569),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_599),
.B(n_466),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_608),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_570),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_599),
.B(n_466),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_564),
.B(n_508),
.Y(n_656)
);

BUFx4f_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_567),
.Y(n_658)
);

CKINVDCx11_ASAP7_75t_R g659 ( 
.A(n_599),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_570),
.Y(n_661)
);

INVx6_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_600),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_565),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_565),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_593),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_602),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_573),
.Y(n_669)
);

BUFx12f_ASAP7_75t_L g670 ( 
.A(n_604),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_622),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_650),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_617),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_626),
.B(n_551),
.Y(n_675)
);

BUFx2_ASAP7_75t_SL g676 ( 
.A(n_624),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_650),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_658),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_615),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_SL g680 ( 
.A1(n_628),
.A2(n_606),
.B1(n_578),
.B2(n_598),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_611),
.B(n_546),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_617),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_619),
.Y(n_683)
);

INVx8_ASAP7_75t_L g684 ( 
.A(n_648),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

BUFx8_ASAP7_75t_L g686 ( 
.A(n_648),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_630),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_633),
.A2(n_582),
.B1(n_572),
.B2(n_547),
.Y(n_688)
);

BUFx8_ASAP7_75t_SL g689 ( 
.A(n_644),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_610),
.Y(n_690)
);

INVx6_ASAP7_75t_L g691 ( 
.A(n_631),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_633),
.A2(n_598),
.B1(n_585),
.B2(n_509),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_633),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_620),
.B(n_667),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_630),
.Y(n_695)
);

CKINVDCx11_ASAP7_75t_R g696 ( 
.A(n_659),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_637),
.A2(n_571),
.B1(n_578),
.B2(n_503),
.Y(n_697)
);

INVx6_ASAP7_75t_L g698 ( 
.A(n_631),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_642),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_642),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_636),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

BUFx8_ASAP7_75t_L g703 ( 
.A(n_638),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_628),
.A2(n_503),
.B1(n_515),
.B2(n_513),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_621),
.A2(n_585),
.B1(n_531),
.B2(n_519),
.Y(n_705)
);

BUFx4f_ASAP7_75t_SL g706 ( 
.A(n_638),
.Y(n_706)
);

CKINVDCx10_ASAP7_75t_R g707 ( 
.A(n_667),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_613),
.A2(n_503),
.B1(n_515),
.B2(n_513),
.Y(n_708)
);

INVx6_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_670),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_636),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_667),
.B(n_528),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_SL g713 ( 
.A1(n_613),
.A2(n_531),
.B1(n_528),
.B2(n_515),
.Y(n_713)
);

INVx6_ASAP7_75t_L g714 ( 
.A(n_631),
.Y(n_714)
);

CKINVDCx11_ASAP7_75t_R g715 ( 
.A(n_645),
.Y(n_715)
);

CKINVDCx11_ASAP7_75t_R g716 ( 
.A(n_645),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_656),
.B(n_587),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_670),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_636),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_641),
.A2(n_513),
.B1(n_544),
.B2(n_509),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_657),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_664),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_657),
.A2(n_618),
.B1(n_662),
.B2(n_631),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_657),
.A2(n_508),
.B1(n_592),
.B2(n_534),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_705),
.A2(n_641),
.B1(n_542),
.B2(n_539),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_705),
.A2(n_641),
.B1(n_542),
.B2(n_539),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_671),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_717),
.A2(n_631),
.B1(n_651),
.B2(n_645),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_SL g730 ( 
.A1(n_688),
.A2(n_662),
.B1(n_625),
.B2(n_663),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_713),
.A2(n_641),
.B1(n_522),
.B2(n_538),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_681),
.B(n_591),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_672),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_712),
.B(n_516),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_677),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_680),
.A2(n_547),
.B1(n_662),
.B2(n_612),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_688),
.A2(n_662),
.B1(n_625),
.B2(n_663),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_675),
.B(n_505),
.Y(n_738)
);

INVx4_ASAP7_75t_SL g739 ( 
.A(n_691),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_SL g740 ( 
.A1(n_680),
.A2(n_713),
.B(n_697),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_691),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_673),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_706),
.A2(n_612),
.B1(n_651),
.B2(n_614),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_693),
.A2(n_612),
.B1(n_651),
.B2(n_614),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

OAI222xp33_ASAP7_75t_L g746 ( 
.A1(n_723),
.A2(n_595),
.B1(n_577),
.B2(n_646),
.C1(n_668),
.C2(n_653),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_703),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_SL g749 ( 
.A1(n_693),
.A2(n_507),
.B(n_462),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_692),
.A2(n_625),
.B1(n_574),
.B2(n_554),
.Y(n_750)
);

BUFx5_ASAP7_75t_L g751 ( 
.A(n_679),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_696),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_685),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_683),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_708),
.A2(n_538),
.B1(n_522),
.B2(n_505),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_720),
.A2(n_492),
.B1(n_483),
.B2(n_486),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_725),
.A2(n_594),
.B(n_477),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_702),
.Y(n_758)
);

OAI21xp33_ASAP7_75t_L g759 ( 
.A1(n_690),
.A2(n_601),
.B(n_511),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_704),
.A2(n_484),
.B1(n_494),
.B2(n_492),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_702),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_689),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_699),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_687),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_691),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_695),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_700),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_684),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_694),
.A2(n_625),
.B1(n_653),
.B2(n_668),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_722),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_724),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_701),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_686),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_718),
.A2(n_494),
.B1(n_486),
.B2(n_646),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_676),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_703),
.A2(n_625),
.B1(n_653),
.B2(n_646),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_718),
.A2(n_471),
.B1(n_463),
.B2(n_524),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_710),
.A2(n_653),
.B1(n_669),
.B2(n_634),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_719),
.A2(n_471),
.B1(n_463),
.B2(n_668),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_721),
.A2(n_666),
.B1(n_506),
.B2(n_511),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_682),
.A2(n_669),
.B1(n_634),
.B2(n_623),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_698),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_674),
.A2(n_506),
.B1(n_597),
.B2(n_666),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_SL g785 ( 
.A1(n_698),
.A2(n_468),
.B1(n_465),
.B2(n_597),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_698),
.A2(n_583),
.B1(n_532),
.B2(n_590),
.Y(n_786)
);

OAI222xp33_ASAP7_75t_L g787 ( 
.A1(n_731),
.A2(n_674),
.B1(n_543),
.B2(n_482),
.C1(n_603),
.C2(n_581),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_734),
.B(n_715),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_732),
.A2(n_714),
.B1(n_709),
.B2(n_466),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_726),
.A2(n_714),
.B1(n_709),
.B2(n_466),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_727),
.A2(n_709),
.B1(n_714),
.B2(n_491),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_759),
.A2(n_510),
.B1(n_491),
.B2(n_716),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_SL g793 ( 
.A1(n_740),
.A2(n_684),
.B1(n_686),
.B2(n_634),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_777),
.A2(n_510),
.B1(n_482),
.B2(n_500),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_730),
.A2(n_501),
.B1(n_607),
.B2(n_669),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_730),
.A2(n_666),
.B1(n_665),
.B2(n_684),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_SL g797 ( 
.A1(n_750),
.A2(n_616),
.B1(n_643),
.B2(n_639),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_737),
.A2(n_476),
.B1(n_520),
.B2(n_529),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_736),
.A2(n_616),
.B1(n_639),
.B2(n_660),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_738),
.A2(n_616),
.B1(n_639),
.B2(n_660),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_737),
.A2(n_529),
.B1(n_580),
.B2(n_579),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_774),
.A2(n_665),
.B1(n_629),
.B2(n_640),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_755),
.A2(n_529),
.B1(n_530),
.B2(n_533),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_775),
.A2(n_643),
.B1(n_654),
.B2(n_660),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_L g805 ( 
.A1(n_749),
.A2(n_766),
.B1(n_733),
.B2(n_745),
.C(n_753),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_784),
.A2(n_623),
.B1(n_627),
.B2(n_661),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_770),
.A2(n_530),
.B1(n_533),
.B2(n_523),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_774),
.A2(n_517),
.B1(n_627),
.B2(n_661),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_784),
.A2(n_629),
.B1(n_640),
.B2(n_647),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_756),
.A2(n_647),
.B1(n_640),
.B2(n_629),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_735),
.B(n_629),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_756),
.A2(n_665),
.B1(n_640),
.B2(n_647),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_760),
.A2(n_665),
.B1(n_647),
.B2(n_655),
.Y(n_813)
);

AOI222xp33_ASAP7_75t_L g814 ( 
.A1(n_746),
.A2(n_576),
.B1(n_602),
.B2(n_536),
.C1(n_514),
.C2(n_479),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_767),
.A2(n_530),
.B1(n_533),
.B2(n_523),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_760),
.A2(n_530),
.B1(n_533),
.B2(n_523),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_728),
.A2(n_523),
.B1(n_533),
.B2(n_654),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_776),
.A2(n_707),
.B(n_655),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_781),
.A2(n_665),
.B1(n_655),
.B2(n_652),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_786),
.B(n_615),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_742),
.A2(n_523),
.B1(n_654),
.B2(n_643),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_763),
.A2(n_499),
.B1(n_495),
.B2(n_635),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_765),
.B(n_615),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_771),
.A2(n_649),
.B1(n_635),
.B2(n_632),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_768),
.A2(n_652),
.B1(n_649),
.B2(n_635),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_769),
.A2(n_649),
.B1(n_635),
.B2(n_632),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_769),
.A2(n_649),
.B1(n_635),
.B2(n_632),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_744),
.A2(n_649),
.B1(n_632),
.B2(n_615),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_764),
.B(n_632),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_768),
.A2(n_652),
.B1(n_496),
.B2(n_464),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_772),
.B(n_295),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_729),
.A2(n_496),
.B1(n_464),
.B2(n_540),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_729),
.A2(n_496),
.B1(n_304),
.B2(n_299),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_779),
.A2(n_496),
.B1(n_304),
.B2(n_299),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_765),
.B(n_783),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_785),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_776),
.A2(n_304),
.B1(n_299),
.B2(n_295),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_780),
.A2(n_304),
.B1(n_299),
.B2(n_295),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_805),
.B(n_748),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_836),
.B(n_748),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_836),
.B(n_758),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_820),
.B(n_785),
.C(n_782),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_820),
.B(n_757),
.C(n_778),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_793),
.A2(n_747),
.B1(n_743),
.B2(n_773),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_835),
.B(n_758),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_SL g846 ( 
.A(n_818),
.B(n_752),
.Y(n_846)
);

AOI221xp5_ASAP7_75t_L g847 ( 
.A1(n_787),
.A2(n_746),
.B1(n_754),
.B2(n_304),
.C(n_299),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_835),
.B(n_761),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_831),
.B(n_761),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_L g850 ( 
.A1(n_792),
.A2(n_741),
.B1(n_762),
.B2(n_739),
.C(n_751),
.Y(n_850)
);

OA211x2_ASAP7_75t_L g851 ( 
.A1(n_788),
.A2(n_751),
.B(n_739),
.C(n_741),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_SL g852 ( 
.A1(n_796),
.A2(n_741),
.B(n_739),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_831),
.B(n_811),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_828),
.B(n_751),
.Y(n_854)
);

OA211x2_ASAP7_75t_L g855 ( 
.A1(n_826),
.A2(n_751),
.B(n_741),
.C(n_51),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_829),
.B(n_751),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_SL g857 ( 
.A1(n_808),
.A2(n_751),
.B1(n_50),
.B2(n_52),
.C(n_53),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_810),
.B(n_194),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_810),
.B(n_806),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_809),
.B(n_48),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_827),
.B(n_55),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_808),
.B(n_56),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_SL g863 ( 
.A1(n_814),
.A2(n_799),
.B(n_797),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_795),
.A2(n_193),
.B1(n_58),
.B2(n_59),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_813),
.B(n_57),
.Y(n_865)
);

XNOR2xp5_ASAP7_75t_L g866 ( 
.A(n_804),
.B(n_62),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_824),
.B(n_63),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_802),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.C(n_71),
.Y(n_868)
);

NAND4xp25_ASAP7_75t_L g869 ( 
.A(n_822),
.B(n_191),
.C(n_74),
.D(n_75),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_790),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_870)
);

OAI221xp5_ASAP7_75t_SL g871 ( 
.A1(n_798),
.A2(n_833),
.B1(n_789),
.B2(n_803),
.C(n_800),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_812),
.B(n_81),
.C(n_83),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_823),
.B(n_187),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_801),
.B(n_823),
.C(n_825),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_819),
.B(n_84),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_832),
.B(n_85),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_816),
.B(n_86),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_791),
.B(n_186),
.Y(n_878)
);

AOI211xp5_ASAP7_75t_L g879 ( 
.A1(n_863),
.A2(n_830),
.B(n_837),
.C(n_90),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_853),
.B(n_821),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_857),
.B(n_834),
.C(n_815),
.Y(n_881)
);

NOR2x1_ASAP7_75t_R g882 ( 
.A(n_860),
.B(n_88),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_853),
.B(n_817),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_848),
.B(n_807),
.Y(n_884)
);

XNOR2xp5_ASAP7_75t_L g885 ( 
.A(n_844),
.B(n_794),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_860),
.A2(n_854),
.B(n_843),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_845),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_845),
.B(n_838),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_849),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_840),
.B(n_89),
.Y(n_890)
);

NAND4xp75_ASAP7_75t_L g891 ( 
.A(n_847),
.B(n_184),
.C(n_95),
.D(n_96),
.Y(n_891)
);

OAI31xp33_ASAP7_75t_L g892 ( 
.A1(n_842),
.A2(n_92),
.A3(n_99),
.B(n_100),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_849),
.B(n_104),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_856),
.B(n_105),
.Y(n_894)
);

OAI211xp5_ASAP7_75t_SL g895 ( 
.A1(n_839),
.A2(n_106),
.B(n_107),
.C(n_108),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_846),
.B(n_111),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_841),
.B(n_112),
.C(n_113),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_859),
.B(n_182),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_869),
.B(n_114),
.C(n_116),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_854),
.B(n_118),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_876),
.B(n_119),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_876),
.B(n_120),
.Y(n_902)
);

XNOR2xp5_ASAP7_75t_L g903 ( 
.A(n_885),
.B(n_879),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_889),
.B(n_852),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_899),
.A2(n_885),
.B1(n_886),
.B2(n_881),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_901),
.B(n_866),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_889),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_886),
.Y(n_908)
);

NAND4xp75_ASAP7_75t_L g909 ( 
.A(n_900),
.B(n_851),
.C(n_855),
.D(n_875),
.Y(n_909)
);

NAND4xp75_ASAP7_75t_SL g910 ( 
.A(n_892),
.B(n_861),
.C(n_867),
.D(n_875),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_893),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_886),
.B(n_858),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_887),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_861),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_898),
.A2(n_895),
.B1(n_891),
.B2(n_901),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_882),
.B(n_862),
.C(n_874),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_894),
.B(n_865),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_894),
.B(n_867),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_883),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_893),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_919),
.Y(n_921)
);

XOR2x2_ASAP7_75t_L g922 ( 
.A(n_903),
.B(n_891),
.Y(n_922)
);

XNOR2x1_ASAP7_75t_L g923 ( 
.A(n_903),
.B(n_902),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_908),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_914),
.B(n_884),
.Y(n_925)
);

OA22x2_ASAP7_75t_L g926 ( 
.A1(n_906),
.A2(n_902),
.B1(n_900),
.B2(n_880),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_904),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_908),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_912),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_927),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_928),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_925),
.Y(n_933)
);

XOR2x2_ASAP7_75t_L g934 ( 
.A(n_923),
.B(n_906),
.Y(n_934)
);

XOR2x2_ASAP7_75t_L g935 ( 
.A(n_923),
.B(n_910),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_921),
.Y(n_936)
);

OA22x2_ASAP7_75t_L g937 ( 
.A1(n_927),
.A2(n_915),
.B1(n_911),
.B2(n_920),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_924),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_929),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_936),
.Y(n_940)
);

OA22x2_ASAP7_75t_L g941 ( 
.A1(n_935),
.A2(n_922),
.B1(n_926),
.B2(n_930),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_931),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_932),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_938),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_932),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_943),
.Y(n_946)
);

OAI322xp33_ASAP7_75t_L g947 ( 
.A1(n_941),
.A2(n_937),
.A3(n_926),
.B1(n_939),
.B2(n_933),
.C1(n_934),
.C2(n_918),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_941),
.A2(n_937),
.B1(n_905),
.B2(n_943),
.Y(n_948)
);

OAI322xp33_ASAP7_75t_L g949 ( 
.A1(n_945),
.A2(n_939),
.A3(n_933),
.B1(n_917),
.B2(n_922),
.C1(n_920),
.C2(n_890),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_948),
.A2(n_944),
.B1(n_940),
.B2(n_942),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_946),
.A2(n_942),
.B1(n_907),
.B2(n_916),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_947),
.A2(n_909),
.B1(n_914),
.B2(n_896),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_SL g953 ( 
.A1(n_949),
.A2(n_864),
.B(n_873),
.C(n_877),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_950),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_951),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_952),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_953),
.B(n_913),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_950),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_952),
.B(n_913),
.Y(n_959)
);

CKINVDCx14_ASAP7_75t_R g960 ( 
.A(n_955),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_958),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_956),
.A2(n_897),
.B1(n_888),
.B2(n_890),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_957),
.A2(n_888),
.B1(n_850),
.B2(n_884),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_962),
.A2(n_957),
.B1(n_882),
.B2(n_883),
.Y(n_966)
);

AO22x2_ASAP7_75t_L g967 ( 
.A1(n_961),
.A2(n_870),
.B1(n_872),
.B2(n_878),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_964),
.Y(n_968)
);

AND4x1_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_868),
.C(n_871),
.D(n_124),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_963),
.B(n_121),
.Y(n_970)
);

AND3x4_ASAP7_75t_L g971 ( 
.A(n_969),
.B(n_960),
.C(n_125),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_122),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_966),
.A2(n_967),
.B1(n_970),
.B2(n_128),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_970),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_970),
.Y(n_975)
);

OA22x2_ASAP7_75t_L g976 ( 
.A1(n_971),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_976)
);

NAND4xp25_ASAP7_75t_L g977 ( 
.A(n_973),
.B(n_130),
.C(n_131),
.D(n_132),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_972),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_972),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_975),
.A2(n_138),
.B1(n_140),
.B2(n_142),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_976),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_979),
.B(n_974),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_977),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_981),
.A2(n_980),
.B1(n_978),
.B2(n_149),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_983),
.A2(n_982),
.B1(n_147),
.B2(n_152),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_985),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_984),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_986),
.A2(n_145),
.B1(n_155),
.B2(n_156),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_987),
.A2(n_159),
.B1(n_161),
.B2(n_166),
.Y(n_989)
);

OAI22xp33_ASAP7_75t_L g990 ( 
.A1(n_986),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_990),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_988),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_991),
.A2(n_989),
.B1(n_173),
.B2(n_174),
.C(n_175),
.Y(n_993)
);

AOI211xp5_ASAP7_75t_L g994 ( 
.A1(n_993),
.A2(n_992),
.B(n_178),
.C(n_179),
.Y(n_994)
);


endmodule