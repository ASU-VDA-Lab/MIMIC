module fake_jpeg_11739_n_509 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_87),
.Y(n_122)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_62),
.B(n_75),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_17),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_63),
.A2(n_103),
.B(n_46),
.Y(n_196)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_71),
.Y(n_200)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_23),
.A2(n_16),
.B(n_1),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_86),
.B(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_105),
.Y(n_123)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_97),
.Y(n_170)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

CKINVDCx9p33_ASAP7_75t_R g199 ( 
.A(n_99),
.Y(n_199)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_100),
.B(n_102),
.Y(n_166)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_0),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_45),
.B1(n_32),
.B2(n_40),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_110),
.A2(n_82),
.B(n_48),
.Y(n_195)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_0),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_112),
.B(n_113),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_1),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_43),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_27),
.Y(n_154)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_47),
.B1(n_31),
.B2(n_35),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_125),
.A2(n_135),
.B1(n_150),
.B2(n_157),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_47),
.B1(n_55),
.B2(n_21),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_127),
.A2(n_176),
.B1(n_191),
.B2(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_50),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_128),
.B(n_159),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_21),
.B(n_55),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_129),
.B(n_196),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_50),
.B1(n_40),
.B2(n_29),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_139),
.A2(n_165),
.B1(n_137),
.B2(n_155),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_140),
.B(n_153),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_45),
.B1(n_32),
.B2(n_29),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_27),
.B(n_5),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_152),
.B(n_167),
.C(n_126),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_154),
.B(n_126),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_73),
.B(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_71),
.B(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_161),
.B(n_175),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_163),
.B(n_172),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_58),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_167),
.A2(n_195),
.B1(n_147),
.B2(n_156),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_101),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_80),
.B(n_13),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_56),
.A2(n_13),
.B1(n_66),
.B2(n_70),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_78),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_79),
.B(n_83),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_88),
.B(n_89),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_201),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_93),
.A2(n_103),
.B1(n_63),
.B2(n_57),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_194),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_95),
.B(n_106),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_190),
.B(n_194),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_57),
.A2(n_103),
.B1(n_54),
.B2(n_52),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_57),
.B(n_62),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_57),
.B(n_62),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_197),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_86),
.Y(n_201)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_125),
.A2(n_192),
.B1(n_128),
.B2(n_177),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_207),
.A2(n_231),
.B(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_199),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_209),
.Y(n_291)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_211),
.B(n_238),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_123),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_239),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_142),
.A2(n_122),
.B(n_129),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_213),
.A2(n_271),
.B(n_204),
.Y(n_299)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_187),
.B(n_159),
.CI(n_175),
.CON(n_221),
.SN(n_221)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_221),
.B(n_222),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_161),
.A2(n_190),
.B1(n_154),
.B2(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_235),
.B1(n_255),
.B2(n_260),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_266),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_133),
.A2(n_149),
.B(n_152),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_252),
.C(n_256),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_233),
.A2(n_246),
.B1(n_269),
.B2(n_237),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_155),
.A2(n_137),
.B1(n_189),
.B2(n_132),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_141),
.A2(n_184),
.B1(n_158),
.B2(n_134),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_171),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_237),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_189),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_243),
.Y(n_289)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_167),
.A2(n_203),
.B1(n_188),
.B2(n_147),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_251),
.B1(n_205),
.B2(n_254),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_136),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_248),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_137),
.A2(n_146),
.B1(n_202),
.B2(n_144),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_247),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_143),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_268),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_146),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_185),
.A2(n_193),
.B1(n_158),
.B2(n_145),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_145),
.B(n_173),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_188),
.A2(n_203),
.B1(n_185),
.B2(n_148),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_148),
.B(n_183),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_251),
.B1(n_265),
.B2(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_183),
.C(n_193),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_259),
.B(n_262),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_131),
.A2(n_138),
.B1(n_151),
.B2(n_169),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_143),
.B(n_169),
.C(n_151),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_263),
.B(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_138),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_267),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_162),
.B(n_181),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_168),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_168),
.A2(n_195),
.B1(n_81),
.B2(n_35),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_181),
.A2(n_187),
.B1(n_191),
.B2(n_127),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_272),
.B1(n_258),
.B2(n_265),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_177),
.A2(n_196),
.B(n_198),
.C(n_194),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_214),
.B(n_215),
.C(n_261),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_187),
.A2(n_191),
.B1(n_127),
.B2(n_159),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_225),
.A2(n_231),
.B1(n_207),
.B2(n_240),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_275),
.A2(n_288),
.B1(n_315),
.B2(n_238),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_300),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_232),
.A2(n_214),
.B(n_211),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_279),
.A2(n_314),
.B(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_267),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_225),
.A2(n_261),
.B1(n_263),
.B2(n_221),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_228),
.B(n_214),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_298),
.B(n_311),
.Y(n_353)
);

OR2x2_ASAP7_75t_SL g343 ( 
.A(n_299),
.B(n_243),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_230),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_241),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_219),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_320),
.Y(n_323)
);

AOI22x1_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_250),
.B1(n_238),
.B2(n_220),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_285),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_217),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_256),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_256),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_317),
.Y(n_340)
);

AOI22x1_ASAP7_75t_SL g314 ( 
.A1(n_272),
.A2(n_258),
.B1(n_235),
.B2(n_216),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_258),
.A2(n_264),
.B1(n_259),
.B2(n_208),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_227),
.B1(n_314),
.B2(n_293),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_218),
.B(n_226),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_262),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_222),
.C(n_266),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_293),
.C(n_303),
.Y(n_378)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_292),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_330),
.Y(n_360)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_294),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_334),
.Y(n_366)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_280),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_342),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_303),
.Y(n_388)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_338),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_253),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_339),
.B(n_359),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_316),
.A2(n_247),
.B1(n_224),
.B2(n_250),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_341),
.A2(n_352),
.B1(n_315),
.B2(n_313),
.Y(n_364)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_SL g368 ( 
.A(n_343),
.B(n_347),
.C(n_351),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_206),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_354),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_287),
.Y(n_361)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_348),
.Y(n_384)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_350),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_304),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_233),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_275),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_304),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_356),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_287),
.B(n_306),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_357),
.A2(n_295),
.B(n_279),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_301),
.B(n_298),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_326),
.B(n_351),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_374),
.B(n_383),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_370),
.B1(n_371),
.B2(n_340),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_286),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_375),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_322),
.A2(n_341),
.B1(n_330),
.B2(n_354),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_322),
.A2(n_273),
.B1(n_305),
.B2(n_284),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_344),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_333),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_295),
.B(n_306),
.Y(n_374)
);

NOR3xp33_ASAP7_75t_SL g375 ( 
.A(n_329),
.B(n_273),
.C(n_297),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_324),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_306),
.B(n_273),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_283),
.B1(n_297),
.B2(n_305),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_390),
.B1(n_340),
.B2(n_337),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_388),
.B(n_389),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_276),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_323),
.A2(n_283),
.B1(n_305),
.B2(n_312),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_394),
.A2(n_395),
.B1(n_414),
.B2(n_365),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_350),
.B1(n_355),
.B2(n_326),
.Y(n_395)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_276),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_416),
.C(n_362),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_327),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_399),
.B(n_413),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_360),
.B(n_353),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_408),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_401),
.A2(n_361),
.B(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

OAI21xp33_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_343),
.B(n_329),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g408 ( 
.A1(n_379),
.A2(n_305),
.B1(n_356),
.B2(n_325),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_349),
.B1(n_331),
.B2(n_348),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_328),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_410),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_356),
.B1(n_346),
.B2(n_282),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_415),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_385),
.B(n_299),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_364),
.A2(n_370),
.B1(n_371),
.B2(n_373),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_289),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_391),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_410),
.Y(n_420)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_424),
.C(n_425),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_416),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_308),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_423),
.A2(n_436),
.B1(n_377),
.B2(n_418),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_378),
.C(n_383),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_389),
.C(n_361),
.Y(n_425)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_414),
.A2(n_365),
.B1(n_363),
.B2(n_367),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_411),
.B1(n_392),
.B2(n_413),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_393),
.A2(n_367),
.B1(n_391),
.B2(n_368),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_437),
.B1(n_412),
.B2(n_405),
.Y(n_448)
);

OR2x4_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_368),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_408),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_375),
.C(n_366),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_397),
.C(n_408),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_395),
.A2(n_402),
.B1(n_404),
.B2(n_394),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_409),
.A2(n_366),
.B1(n_375),
.B2(n_377),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_439),
.A2(n_392),
.B(n_400),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_440),
.B(n_452),
.Y(n_461)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_439),
.A2(n_417),
.B1(n_406),
.B2(n_408),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_443),
.A2(n_448),
.B1(n_426),
.B2(n_430),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_455),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_446),
.A2(n_419),
.B(n_429),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_449),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_369),
.C(n_382),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_451),
.C(n_454),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_369),
.C(n_281),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_439),
.A2(n_381),
.B(n_380),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_281),
.C(n_282),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_308),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_457),
.C(n_430),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_436),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_470),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_437),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_433),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_466),
.B(n_468),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_429),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_458),
.B(n_450),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_476),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_461),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_464),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_451),
.C(n_444),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_460),
.C(n_444),
.Y(n_490)
);

AO221x1_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_467),
.B1(n_463),
.B2(n_427),
.C(n_469),
.Y(n_478)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_478),
.Y(n_482)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_467),
.Y(n_479)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_459),
.A2(n_443),
.B(n_453),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_481),
.A2(n_441),
.B(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_480),
.A2(n_463),
.B1(n_428),
.B2(n_473),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_486),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_423),
.B1(n_459),
.B2(n_432),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_490),
.B(n_477),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_496),
.C(n_460),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_482),
.A2(n_475),
.B1(n_479),
.B2(n_431),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_494),
.A2(n_489),
.B1(n_483),
.B2(n_481),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_477),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_475),
.C(n_488),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_498),
.B(n_499),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_497),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_504),
.Y(n_505)
);

AO21x1_ASAP7_75t_L g504 ( 
.A1(n_501),
.A2(n_494),
.B(n_495),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_502),
.A2(n_498),
.B(n_483),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_505),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_438),
.Y(n_509)
);


endmodule