module fake_jpeg_2021_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_15),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

OA22x2_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_38),
.B1(n_41),
.B2(n_2),
.Y(n_62)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_62),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_35),
.C(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_47),
.C(n_36),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_55),
.B(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_40),
.B1(n_43),
.B2(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_22),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_0),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_53),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_75),
.Y(n_86)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_35),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_61),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_84),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_87),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_44),
.A3(n_52),
.B1(n_55),
.B2(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_50),
.B1(n_54),
.B2(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_4),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_70),
.C(n_72),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_103),
.C(n_107),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_102),
.B(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_76),
.C(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_16),
.B(n_28),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_76),
.Y(n_106)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_96),
.A3(n_103),
.B1(n_17),
.B2(n_20),
.C(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_116),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_93),
.B(n_94),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_113),
.B(n_8),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_14),
.B(n_27),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_26),
.C(n_25),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_117),
.C(n_116),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_6),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_11),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_24),
.C(n_23),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_115),
.C(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_124),
.C(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_120),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_134),
.B(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_120),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_130),
.Y(n_139)
);


endmodule