module fake_ibex_1073_n_993 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_993);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_993;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_980;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_439;
wire n_299;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_890;
wire n_874;
wire n_816;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_46),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_125),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_101),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_70),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_50),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_19),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_56),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_78),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_21),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_90),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_58),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_69),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_64),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_44),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_37),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_79),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_184),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_37),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_163),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_43),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_49),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_124),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_132),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_108),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_59),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_127),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_24),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_34),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_150),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_159),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_8),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_171),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_147),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_142),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_60),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_38),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_91),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_114),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_84),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_97),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_111),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_9),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_41),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_34),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_174),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_117),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_77),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_112),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_85),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_175),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_155),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_66),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_165),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_104),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_33),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_143),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_81),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_183),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_71),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_40),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_106),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_75),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_63),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_11),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_119),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_25),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_146),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_178),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_256),
.B(n_45),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_218),
.B(n_0),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_218),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_231),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_188),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_188),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_8),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_212),
.B(n_10),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_11),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_244),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_186),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_12),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_12),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_241),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_214),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_234),
.A2(n_283),
.B(n_237),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_262),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_269),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_212),
.B(n_14),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_290),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g350 ( 
.A1(n_234),
.A2(n_88),
.B(n_185),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_239),
.B(n_16),
.Y(n_351)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_244),
.Y(n_352)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_270),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_270),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_223),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_227),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_196),
.B(n_48),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_237),
.A2(n_92),
.B(n_180),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_283),
.A2(n_87),
.B(n_179),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_295),
.B(n_17),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_189),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_207),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_R g367 ( 
.A1(n_257),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_190),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_241),
.B(n_196),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_241),
.B(n_22),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_233),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_281),
.B(n_22),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_193),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_253),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_270),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_295),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_250),
.B(n_23),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_310),
.A2(n_96),
.B(n_177),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_199),
.Y(n_384)
);

CKINVDCx11_ASAP7_75t_R g385 ( 
.A(n_191),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_263),
.B(n_24),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_332),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_202),
.C(n_200),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_205),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_387),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_284),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_323),
.A2(n_289),
.B1(n_245),
.B2(n_191),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_347),
.B(n_337),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_261),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_264),
.B1(n_272),
.B2(n_308),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

BUFx6f_ASAP7_75t_SL g412 ( 
.A(n_311),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_203),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_337),
.B(n_208),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_209),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_339),
.B(n_205),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_345),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_348),
.B(n_273),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_279),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_364),
.B(n_201),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_349),
.A2(n_255),
.B1(n_198),
.B2(n_245),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_352),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_318),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

NAND3xp33_ASAP7_75t_L g438 ( 
.A(n_364),
.B(n_221),
.C(n_219),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_368),
.B(n_222),
.Y(n_439)
);

AND3x2_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_215),
.C(n_211),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_362),
.A2(n_310),
.B(n_228),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_319),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_368),
.B(n_204),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_369),
.B(n_206),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_314),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_369),
.A2(n_282),
.B1(n_285),
.B2(n_306),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_373),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_374),
.B(n_210),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_314),
.B(n_291),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_374),
.B(n_213),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_373),
.B(n_294),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_326),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_380),
.B(n_217),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_380),
.B(n_220),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_384),
.A2(n_302),
.B1(n_307),
.B2(n_305),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_318),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_356),
.B(n_281),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_384),
.B(n_225),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_359),
.A2(n_309),
.B1(n_303),
.B2(n_224),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_343),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_322),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_313),
.B(n_232),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_322),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_322),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_335),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_334),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_367),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_343),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_322),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_315),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_342),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_330),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_330),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_325),
.A2(n_194),
.B1(n_259),
.B2(n_255),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_358),
.B(n_226),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_330),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_391),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_340),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_391),
.A2(n_338),
.B1(n_346),
.B2(n_289),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_342),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_427),
.A2(n_360),
.B(n_350),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_357),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_409),
.B(n_198),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_400),
.B(n_382),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_427),
.A2(n_357),
.B1(n_375),
.B2(n_312),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_375),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_375),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_409),
.B(n_451),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_428),
.A2(n_386),
.B1(n_333),
.B2(n_315),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_417),
.A2(n_420),
.B(n_439),
.C(n_455),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_316),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_399),
.B(n_316),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_428),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_425),
.B(n_324),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_432),
.B(n_229),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_433),
.A2(n_360),
.B(n_350),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_433),
.A2(n_333),
.B1(n_324),
.B2(n_328),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_399),
.B(n_328),
.Y(n_507)
);

AO22x1_ASAP7_75t_L g508 ( 
.A1(n_431),
.A2(n_365),
.B1(n_259),
.B2(n_230),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_408),
.B(n_329),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_432),
.B(n_235),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_329),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_444),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_390),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_412),
.A2(n_280),
.B1(n_249),
.B2(n_251),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_412),
.B(n_236),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_402),
.B(n_293),
.C(n_243),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_434),
.B(n_350),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_394),
.B(n_396),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_430),
.B(n_238),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_401),
.B(n_350),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_446),
.B(n_242),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_398),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_447),
.B(n_248),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_456),
.B(n_258),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_445),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_265),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_414),
.B(n_246),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_409),
.B(n_247),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_401),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_412),
.A2(n_299),
.B1(n_266),
.B2(n_286),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_360),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_445),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_267),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_454),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_405),
.B(n_271),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2x1_ASAP7_75t_L g542 ( 
.A(n_451),
.B(n_360),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_451),
.B(n_277),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_461),
.B(n_278),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_453),
.B(n_288),
.Y(n_547)
);

AND3x1_ASAP7_75t_L g548 ( 
.A(n_440),
.B(n_195),
.C(n_216),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_477),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_464),
.B(n_296),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_415),
.B(n_297),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_457),
.B(n_298),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_393),
.A2(n_383),
.B(n_361),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_457),
.B(n_301),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_429),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

AND2x6_ASAP7_75t_SL g560 ( 
.A(n_469),
.B(n_195),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_469),
.B(n_361),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_361),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_482),
.B(n_383),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_462),
.B(n_383),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_454),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_410),
.B(n_26),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_415),
.B(n_343),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_443),
.A2(n_393),
.B1(n_438),
.B2(n_466),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_388),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_389),
.B(n_353),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_562),
.A2(n_397),
.B(n_389),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_502),
.A2(n_426),
.B(n_411),
.Y(n_573)
);

CKINVDCx10_ASAP7_75t_R g574 ( 
.A(n_512),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_567),
.A2(n_469),
.B1(n_481),
.B2(n_419),
.Y(n_575)
);

CKINVDCx8_ASAP7_75t_R g576 ( 
.A(n_541),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_469),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_485),
.B(n_424),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_502),
.A2(n_411),
.B(n_419),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_505),
.A2(n_442),
.B(n_395),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_542),
.A2(n_489),
.B(n_555),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_450),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_392),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_557),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

O2A1O1Ixp5_ASAP7_75t_L g586 ( 
.A1(n_563),
.A2(n_403),
.B(n_404),
.C(n_406),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_503),
.B(n_392),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_492),
.B(n_474),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_516),
.A2(n_407),
.B1(n_421),
.B2(n_418),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_513),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_497),
.A2(n_543),
.B(n_532),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_498),
.A2(n_474),
.B1(n_407),
.B2(n_416),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_523),
.B(n_404),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_503),
.B(n_406),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_529),
.B(n_416),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_558),
.Y(n_596)
);

BUFx8_ASAP7_75t_L g597 ( 
.A(n_533),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_423),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_423),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_487),
.A2(n_467),
.B1(n_353),
.B2(n_354),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_550),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_495),
.B(n_467),
.Y(n_603)
);

OAI22x1_ASAP7_75t_L g604 ( 
.A1(n_514),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_27),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_496),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_501),
.B(n_28),
.Y(n_607)
);

HB1xp67_ASAP7_75t_SL g608 ( 
.A(n_516),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_528),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_538),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_508),
.Y(n_612)
);

AO21x1_ASAP7_75t_L g613 ( 
.A1(n_520),
.A2(n_476),
.B(n_435),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_509),
.B(n_30),
.Y(n_614)
);

A2O1A1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_540),
.A2(n_331),
.B(n_376),
.C(n_354),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_498),
.A2(n_353),
.B1(n_354),
.B2(n_331),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_32),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_531),
.B(n_32),
.Y(n_619)
);

AO21x1_ASAP7_75t_L g620 ( 
.A1(n_520),
.A2(n_471),
.B(n_435),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_33),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_506),
.A2(n_354),
.B1(n_331),
.B2(n_376),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_35),
.Y(n_623)
);

OAI22x1_ASAP7_75t_L g624 ( 
.A1(n_534),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_545),
.A2(n_331),
.B(n_376),
.C(n_479),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_36),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_546),
.A2(n_564),
.B(n_517),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_517),
.A2(n_468),
.B(n_480),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_488),
.B(n_39),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_557),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_535),
.A2(n_331),
.B1(n_376),
.B2(n_479),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_556),
.B(n_42),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_547),
.B(n_475),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_569),
.B(n_475),
.C(n_376),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_504),
.B(n_475),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_547),
.B(n_475),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_569),
.B(n_463),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_548),
.A2(n_476),
.B1(n_471),
.B2(n_470),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_553),
.Y(n_641)
);

NOR2x1_ASAP7_75t_SL g642 ( 
.A(n_561),
.B(n_463),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_559),
.Y(n_643)
);

AO32x2_ASAP7_75t_L g644 ( 
.A1(n_561),
.A2(n_483),
.A3(n_463),
.B1(n_53),
.B2(n_54),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_51),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_536),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_494),
.B(n_52),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_565),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_486),
.A2(n_65),
.B(n_68),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_570),
.A2(n_526),
.B1(n_522),
.B2(n_527),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_490),
.A2(n_72),
.B(n_74),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_597),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_578),
.B(n_530),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_597),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_577),
.A2(n_525),
.B1(n_519),
.B2(n_521),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_627),
.A2(n_537),
.B(n_524),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_580),
.A2(n_571),
.B(n_552),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_518),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_585),
.B(n_598),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_586),
.A2(n_568),
.B(n_510),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_620),
.A2(n_560),
.A3(n_80),
.B(n_82),
.Y(n_663)
);

NOR4xp25_ASAP7_75t_L g664 ( 
.A(n_575),
.B(n_619),
.C(n_621),
.D(n_614),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_590),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_SL g666 ( 
.A1(n_647),
.A2(n_76),
.B(n_83),
.C(n_86),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_587),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_592),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_577),
.B(n_99),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_577),
.B(n_102),
.Y(n_671)
);

AO32x2_ASAP7_75t_L g672 ( 
.A1(n_640),
.A2(n_120),
.A3(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_572),
.A2(n_128),
.B(n_130),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_643),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_642),
.A2(n_131),
.A3(n_133),
.B(n_136),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_607),
.A2(n_137),
.B(n_138),
.C(n_139),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_595),
.B(n_140),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_588),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_595),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_649),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_582),
.B(n_157),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_583),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_162),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_SL g684 ( 
.A(n_576),
.B(n_168),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_591),
.A2(n_170),
.B(n_172),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_612),
.B(n_606),
.Y(n_687)
);

BUFx2_ASAP7_75t_R g688 ( 
.A(n_574),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_625),
.A2(n_616),
.A3(n_615),
.B(n_622),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_632),
.B(n_624),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_618),
.A2(n_623),
.B(n_626),
.C(n_630),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_645),
.A2(n_652),
.A3(n_650),
.B(n_604),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_573),
.A2(n_579),
.B(n_594),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_600),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_574),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_635),
.A2(n_638),
.B(n_601),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_617),
.Y(n_698)
);

BUFx12f_ASAP7_75t_L g699 ( 
.A(n_637),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_SL g700 ( 
.A(n_648),
.B(n_584),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_SL g701 ( 
.A1(n_602),
.A2(n_599),
.B(n_633),
.C(n_646),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

AO32x2_ASAP7_75t_L g703 ( 
.A1(n_644),
.A2(n_648),
.A3(n_608),
.B1(n_589),
.B2(n_651),
.Y(n_703)
);

BUFx5_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_603),
.A2(n_611),
.B(n_593),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_641),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_631),
.B(n_644),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_644),
.B(n_578),
.Y(n_709)
);

AO31x2_ASAP7_75t_L g710 ( 
.A1(n_613),
.A2(n_620),
.A3(n_581),
.B(n_627),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_577),
.A2(n_587),
.B1(n_594),
.B2(n_585),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_588),
.A2(n_431),
.B1(n_492),
.B2(n_612),
.Y(n_712)
);

INVx6_ASAP7_75t_L g713 ( 
.A(n_597),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_533),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_577),
.A2(n_587),
.B1(n_594),
.B2(n_585),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_596),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_583),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_578),
.B(n_485),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_590),
.Y(n_719)
);

AO31x2_ASAP7_75t_L g720 ( 
.A1(n_613),
.A2(n_620),
.A3(n_581),
.B(n_627),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_597),
.Y(n_721)
);

AO21x2_ASAP7_75t_L g722 ( 
.A1(n_581),
.A2(n_639),
.B(n_636),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_581),
.A2(n_580),
.B(n_629),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_581),
.A2(n_580),
.B(n_629),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_578),
.B(n_533),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_578),
.B(n_533),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_597),
.B(n_492),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_578),
.B(n_485),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_577),
.A2(n_587),
.B1(n_594),
.B2(n_585),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_607),
.A2(n_618),
.B(n_499),
.C(n_614),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_590),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_607),
.A2(n_618),
.B(n_499),
.C(n_614),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_628),
.B(n_529),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_607),
.A2(n_618),
.B(n_499),
.C(n_614),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_590),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_578),
.B(n_485),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_628),
.B(n_529),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_581),
.A2(n_580),
.B(n_629),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_718),
.B(n_728),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_736),
.B(n_733),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_723),
.A2(n_724),
.B(n_738),
.Y(n_741)
);

AND2x2_ASAP7_75t_SL g742 ( 
.A(n_721),
.B(n_679),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_658),
.A2(n_691),
.B(n_701),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_702),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_665),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_667),
.B(n_661),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_706),
.Y(n_747)
);

CKINVDCx6p67_ASAP7_75t_R g748 ( 
.A(n_665),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_716),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_677),
.B(n_737),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_664),
.B(n_655),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_694),
.A2(n_730),
.B(n_734),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_677),
.B(n_713),
.Y(n_753)
);

AOI221xp5_ASAP7_75t_L g754 ( 
.A1(n_714),
.A2(n_725),
.B1(n_726),
.B2(n_711),
.C(n_729),
.Y(n_754)
);

NAND2x1p5_ASAP7_75t_L g755 ( 
.A(n_665),
.B(n_721),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_732),
.A2(n_709),
.B(n_697),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_674),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_680),
.B(n_687),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_713),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_681),
.A2(n_722),
.B(n_708),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_656),
.Y(n_762)
);

AOI222xp33_ASAP7_75t_L g763 ( 
.A1(n_715),
.A2(n_727),
.B1(n_693),
.B2(n_696),
.C1(n_671),
.C2(n_660),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_698),
.Y(n_765)
);

BUFx8_ASAP7_75t_SL g766 ( 
.A(n_719),
.Y(n_766)
);

AO21x2_ASAP7_75t_L g767 ( 
.A1(n_662),
.A2(n_673),
.B(n_695),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_700),
.B(n_690),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_670),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_717),
.B(n_657),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_683),
.A2(n_685),
.B(n_705),
.Y(n_771)
);

INVx4_ASAP7_75t_SL g772 ( 
.A(n_719),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_688),
.Y(n_773)
);

OA21x2_ASAP7_75t_L g774 ( 
.A1(n_676),
.A2(n_703),
.B(n_710),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_666),
.A2(n_659),
.B(n_669),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_707),
.B(n_735),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_690),
.Y(n_777)
);

OA21x2_ASAP7_75t_L g778 ( 
.A1(n_703),
.A2(n_710),
.B(n_720),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_684),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_678),
.A2(n_707),
.B(n_712),
.Y(n_781)
);

BUFx6f_ASAP7_75t_SL g782 ( 
.A(n_731),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_699),
.Y(n_783)
);

AO31x2_ASAP7_75t_L g784 ( 
.A1(n_663),
.A2(n_672),
.A3(n_692),
.B(n_689),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_686),
.B(n_672),
.Y(n_785)
);

AND2x6_ASAP7_75t_L g786 ( 
.A(n_704),
.B(n_686),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_704),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_675),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_675),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_668),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_668),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_714),
.B(n_578),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_677),
.B(n_713),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_665),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_733),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_714),
.B(n_578),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_668),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_714),
.B(n_578),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_706),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_665),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_677),
.B(n_713),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_668),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_733),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_668),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_702),
.Y(n_805)
);

AOI221xp5_ASAP7_75t_L g806 ( 
.A1(n_718),
.A2(n_736),
.B1(n_728),
.B2(n_516),
.C(n_575),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_668),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_SL g808 ( 
.A1(n_711),
.A2(n_431),
.B1(n_588),
.B2(n_715),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_718),
.B(n_431),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_677),
.B(n_713),
.Y(n_810)
);

CKINVDCx6p67_ASAP7_75t_R g811 ( 
.A(n_748),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_741),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_752),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_751),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_765),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_753),
.B(n_793),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_808),
.A2(n_754),
.B(n_809),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_751),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_746),
.B(n_758),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_740),
.B(n_762),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_746),
.B(n_744),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_786),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_747),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_747),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_749),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_750),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_753),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_753),
.B(n_793),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_793),
.Y(n_829)
);

BUFx12f_ASAP7_75t_L g830 ( 
.A(n_759),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_757),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_787),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_801),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_801),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_754),
.A2(n_806),
.B(n_743),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_801),
.B(n_810),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_810),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_790),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_806),
.A2(n_781),
.B(n_771),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_791),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_786),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_739),
.A2(n_796),
.B1(n_792),
.B2(n_798),
.C(n_769),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_797),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_802),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_755),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_805),
.B(n_807),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_739),
.B(n_763),
.Y(n_847)
);

OA21x2_ASAP7_75t_L g848 ( 
.A1(n_775),
.A2(n_756),
.B(n_761),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_804),
.Y(n_849)
);

BUFx4f_ASAP7_75t_SL g850 ( 
.A(n_759),
.Y(n_850)
);

OA21x2_ASAP7_75t_L g851 ( 
.A1(n_756),
.A2(n_788),
.B(n_789),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_785),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_764),
.B(n_770),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_770),
.B(n_777),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_810),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_786),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_763),
.B(n_778),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_779),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_795),
.B(n_750),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_803),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_766),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_742),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_795),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_857),
.B(n_778),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_857),
.B(n_784),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_819),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_832),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_812),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_862),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_813),
.B(n_774),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_819),
.B(n_768),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_814),
.B(n_767),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_818),
.B(n_781),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_821),
.B(n_780),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_847),
.B(n_760),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_842),
.B(n_747),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_821),
.B(n_799),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_817),
.A2(n_745),
.B1(n_794),
.B2(n_800),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_852),
.B(n_799),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_859),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_846),
.B(n_783),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_839),
.B(n_776),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_835),
.A2(n_776),
.B1(n_773),
.B2(n_782),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_853),
.B(n_772),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_853),
.B(n_772),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_854),
.B(n_782),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_865),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_845),
.Y(n_890)
);

INVx4_ASAP7_75t_R g891 ( 
.A(n_845),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_846),
.B(n_825),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_815),
.B(n_831),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_861),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_R g895 ( 
.A(n_811),
.B(n_863),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_866),
.B(n_851),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_871),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_866),
.B(n_854),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_894),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_867),
.B(n_851),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_870),
.B(n_822),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_869),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_875),
.B(n_851),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_868),
.B(n_840),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_875),
.B(n_848),
.Y(n_905)
);

INVxp33_ASAP7_75t_L g906 ( 
.A(n_895),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_877),
.B(n_838),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_869),
.B(n_838),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_892),
.B(n_848),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_883),
.B(n_824),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_869),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_890),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_890),
.B(n_864),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_899),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_874),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_910),
.A2(n_884),
.B1(n_878),
.B2(n_816),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_912),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_898),
.B(n_874),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_907),
.B(n_892),
.Y(n_919)
);

AND2x4_ASAP7_75t_SL g920 ( 
.A(n_911),
.B(n_816),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_900),
.B(n_909),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_897),
.Y(n_922)
);

NOR2x1_ASAP7_75t_L g923 ( 
.A(n_913),
.B(n_816),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_909),
.B(n_872),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_902),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_897),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_896),
.B(n_901),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_907),
.B(n_889),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_904),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_915),
.B(n_896),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_929),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_922),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_922),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_903),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_926),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_915),
.B(n_908),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_923),
.B(n_912),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_914),
.B(n_904),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_921),
.B(n_905),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_917),
.Y(n_940)
);

NOR2x1_ASAP7_75t_L g941 ( 
.A(n_938),
.B(n_816),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_934),
.B(n_918),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_931),
.A2(n_916),
.B1(n_927),
.B2(n_928),
.Y(n_943)
);

CKINVDCx14_ASAP7_75t_R g944 ( 
.A(n_934),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_939),
.B(n_924),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_940),
.A2(n_927),
.B1(n_836),
.B2(n_828),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_936),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_930),
.B(n_906),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_937),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_940),
.A2(n_927),
.B(n_919),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_939),
.B(n_924),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_937),
.A2(n_836),
.B1(n_828),
.B2(n_881),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_932),
.A2(n_884),
.B1(n_828),
.B2(n_836),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_L g954 ( 
.A(n_944),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_948),
.A2(n_881),
.B1(n_836),
.B2(n_828),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_949),
.B(n_917),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_949),
.A2(n_863),
.B1(n_850),
.B2(n_864),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_SL g958 ( 
.A1(n_950),
.A2(n_891),
.B(n_826),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_R g959 ( 
.A(n_947),
.B(n_811),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_942),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_959),
.B(n_941),
.Y(n_961)
);

AOI221xp5_ASAP7_75t_L g962 ( 
.A1(n_957),
.A2(n_943),
.B1(n_945),
.B2(n_951),
.C(n_953),
.Y(n_962)
);

AOI221xp5_ASAP7_75t_L g963 ( 
.A1(n_956),
.A2(n_933),
.B1(n_935),
.B2(n_946),
.C(n_858),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_SL g964 ( 
.A1(n_962),
.A2(n_954),
.B1(n_955),
.B2(n_960),
.C(n_885),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_961),
.B(n_952),
.Y(n_965)
);

NAND3x1_ASAP7_75t_L g966 ( 
.A(n_964),
.B(n_963),
.C(n_860),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_L g967 ( 
.A(n_965),
.B(n_823),
.C(n_837),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_966),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_967),
.B(n_830),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_969),
.A2(n_958),
.B(n_955),
.Y(n_970)
);

XNOR2xp5_ASAP7_75t_L g971 ( 
.A(n_968),
.B(n_827),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_971),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_970),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_970),
.A2(n_830),
.B1(n_880),
.B2(n_888),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_973),
.A2(n_888),
.B(n_855),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_972),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_974),
.A2(n_823),
.B1(n_833),
.B2(n_834),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_973),
.A2(n_829),
.B1(n_925),
.B2(n_882),
.Y(n_978)
);

OAI22x1_ASAP7_75t_L g979 ( 
.A1(n_973),
.A2(n_820),
.B1(n_841),
.B2(n_856),
.Y(n_979)
);

NAND4xp25_ASAP7_75t_SL g980 ( 
.A(n_976),
.B(n_879),
.C(n_886),
.D(n_887),
.Y(n_980)
);

XNOR2xp5_ASAP7_75t_L g981 ( 
.A(n_978),
.B(n_886),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_975),
.B(n_876),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_979),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_977),
.A2(n_893),
.B(n_843),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_980),
.A2(n_890),
.B1(n_887),
.B2(n_841),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_985),
.A2(n_844),
.B(n_849),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_983),
.B(n_920),
.Y(n_988)
);

XNOR2xp5_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_876),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_988),
.B(n_982),
.Y(n_990)
);

AO21x2_ASAP7_75t_L g991 ( 
.A1(n_987),
.A2(n_984),
.B(n_873),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_989),
.A2(n_986),
.B(n_849),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_990),
.A2(n_991),
.B1(n_992),
.B2(n_920),
.Y(n_993)
);


endmodule