module fake_jpeg_10376_n_24 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_2),
.A2(n_6),
.B1(n_1),
.B2(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_4),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_9),
.B1(n_13),
.B2(n_8),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_14),
.C(n_15),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.Y(n_23)
);

AOI221xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_20),
.B1(n_21),
.B2(n_19),
.C(n_18),
.Y(n_24)
);


endmodule