module real_jpeg_28667_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_286;
wire n_166;
wire n_221;
wire n_300;
wire n_176;
wire n_215;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_293;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_283;
wire n_85;
wire n_81;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx5_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_0),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_1),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_1),
.A2(n_77),
.B1(n_78),
.B2(n_152),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_152),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_152),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_73),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_29),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_2),
.A2(n_29),
.B(n_196),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_156),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_48),
.B(n_52),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_2),
.B(n_122),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_2),
.A2(n_90),
.B1(n_93),
.B2(n_244),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_41),
.B1(n_48),
.B2(n_51),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_7),
.A2(n_48),
.B1(n_51),
.B2(n_58),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_77),
.B1(n_78),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_8),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_128),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_9),
.A2(n_45),
.B1(n_77),
.B2(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_10),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_174)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_12),
.A2(n_77),
.B1(n_78),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_12),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_158),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_158),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_48),
.B1(n_51),
.B2(n_158),
.Y(n_244)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_87),
.B2(n_88),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_24),
.B(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_70),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_25),
.A2(n_32),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_25),
.A2(n_32),
.B1(n_151),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_25),
.A2(n_32),
.B1(n_183),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_27),
.B(n_34),
.Y(n_197)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_30),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_29),
.B(n_74),
.Y(n_172)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_30),
.A2(n_82),
.B1(n_155),
.B2(n_172),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_30),
.A2(n_33),
.A3(n_36),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_32),
.B(n_169),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_34),
.A2(n_50),
.B(n_156),
.C(n_223),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_38),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_43),
.A2(n_55),
.B(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_47),
.A2(n_55),
.B1(n_99),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_47),
.A2(n_53),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_47),
.A2(n_55),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_47),
.A2(n_55),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_47),
.A2(n_55),
.B1(n_203),
.B2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_47),
.B(n_156),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_51),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_55),
.A2(n_64),
.B(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_85),
.B2(n_86),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_67),
.A2(n_69),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_80),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_72),
.A2(n_126),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_72),
.A2(n_126),
.B1(n_127),
.B2(n_164),
.Y(n_280)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_73),
.B(n_102),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_81),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_78),
.Y(n_82)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_78),
.B(n_156),
.CON(n_155),
.SN(n_155)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_97),
.B(n_101),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_89),
.A2(n_98),
.B1(n_108),
.B2(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_90),
.A2(n_93),
.B1(n_141),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_90),
.A2(n_117),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_90),
.A2(n_236),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_91),
.A2(n_96),
.B(n_143),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_91),
.A2(n_118),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_94),
.A2(n_114),
.B(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_94),
.B(n_156),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_98),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_105),
.B(n_109),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_110),
.A2(n_111),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.C(n_124),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_112),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_113),
.B(n_119),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_144),
.Y(n_143)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_118),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_300),
.B(n_305),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_287),
.B(n_299),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_187),
.B(n_268),
.C(n_286),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_175),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_136),
.B(n_175),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_159),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_138),
.B(n_146),
.C(n_159),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_139),
.B(n_140),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_154),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_170),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_161),
.B(n_166),
.C(n_170),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_176),
.A2(n_177),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_267),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_260),
.B(n_266),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_214),
.B(n_259),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_205),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_191),
.B(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.C(n_201),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_192),
.A2(n_193),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_212),
.C(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_253),
.B(n_258),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_232),
.B(n_252),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_224),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_240),
.B(n_251),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_238),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_246),
.B(n_250),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_284),
.B2(n_285),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_276),
.C(n_285),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_279),
.C(n_282),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.C(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);


endmodule