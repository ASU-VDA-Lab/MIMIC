module fake_jpeg_7967_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_40),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_30),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_84)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_23),
.B1(n_29),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_26),
.B1(n_36),
.B2(n_28),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_32),
.B1(n_21),
.B2(n_19),
.Y(n_83)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_20),
.Y(n_82)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_39),
.B1(n_25),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_83),
.B1(n_16),
.B2(n_21),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_72),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_54),
.C(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_86),
.B(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_30),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_37),
.C(n_42),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_37),
.C(n_42),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_94),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_97),
.B(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_112),
.B1(n_88),
.B2(n_52),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_69),
.B(n_70),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_40),
.B(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_48),
.B1(n_39),
.B2(n_16),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_71),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_88),
.B1(n_64),
.B2(n_68),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_43),
.B1(n_67),
.B2(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_126),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_122),
.B(n_81),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_131),
.B1(n_68),
.B2(n_52),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_56),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_132),
.B1(n_89),
.B2(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_53),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_58),
.Y(n_152)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_57),
.B1(n_45),
.B2(n_65),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_134),
.B1(n_101),
.B2(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_112),
.B1(n_98),
.B2(n_90),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_98),
.B(n_117),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_145),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_103),
.B(n_97),
.C(n_109),
.D(n_96),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_96),
.C(n_40),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_146),
.C(n_158),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_40),
.B(n_38),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_105),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_122),
.B(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_59),
.B1(n_68),
.B2(n_81),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_113),
.B1(n_126),
.B2(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_2),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_35),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_30),
.B(n_22),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_174),
.B1(n_147),
.B2(n_159),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_177),
.B1(n_140),
.B2(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_135),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_124),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_162),
.B(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_146),
.C(n_136),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_144),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_155),
.B1(n_154),
.B2(n_131),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_190),
.B1(n_192),
.B2(n_170),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_173),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_151),
.B1(n_147),
.B2(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_125),
.B1(n_145),
.B2(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_58),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_194),
.C(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_78),
.C(n_22),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_78),
.C(n_22),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_165),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_78),
.C(n_22),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_177),
.C(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_207),
.B1(n_211),
.B2(n_213),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_203),
.B(n_208),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_170),
.B(n_167),
.C(n_161),
.Y(n_205)
);

OA21x2_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_167),
.B(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.C(n_194),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_18),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g215 ( 
.A(n_204),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_6),
.B(n_7),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.C(n_221),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_196),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_193),
.B1(n_198),
.B2(n_18),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_18),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_3),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_5),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_201),
.C(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_232),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_5),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_15),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_219),
.B1(n_224),
.B2(n_8),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_239),
.B1(n_230),
.B2(n_226),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_15),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_10),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_7),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_9),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_240),
.Y(n_241)
);

AOI21x1_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_243),
.B(n_238),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_10),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_10),
.C(n_11),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_246),
.A2(n_11),
.B(n_12),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_238),
.A3(n_237),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_11),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_251),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_247),
.Y(n_254)
);


endmodule