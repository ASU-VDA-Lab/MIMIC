module real_jpeg_31577_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

OAI22x1_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_58),
.B1(n_72),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_58),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_1),
.A2(n_58),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_4),
.Y(n_236)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_4),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_167),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_5),
.A2(n_167),
.B1(n_225),
.B2(n_302),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_5),
.A2(n_167),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_6),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_6),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_69),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_11),
.A2(n_25),
.B1(n_124),
.B2(n_128),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g233 ( 
.A1(n_11),
.A2(n_25),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g297 ( 
.A(n_11),
.B(n_55),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_11),
.B(n_209),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g359 ( 
.A1(n_11),
.A2(n_292),
.A3(n_360),
.B1(n_365),
.B2(n_371),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_274),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_272),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_239),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_15),
.B(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_171),
.C(n_219),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_17),
.B(n_219),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_86),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_SL g269 ( 
.A(n_18),
.B(n_270),
.C(n_271),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_52),
.B(n_63),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_19),
.B(n_325),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_19),
.B(n_52),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_20),
.B(n_53),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_20),
.A2(n_30),
.B(n_53),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_24),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_25),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_25),
.A2(n_199),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_25),
.B(n_204),
.Y(n_284)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_25),
.A2(n_292),
.A3(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_25),
.B(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_25),
.B(n_40),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_25),
.B(n_76),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_27),
.Y(n_224)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_30),
.B(n_54),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_30),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_30),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_40),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_36),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_47),
.Y(n_238)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_52),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_52),
.B(n_300),
.Y(n_339)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_53),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_53),
.B(n_301),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_55),
.B(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_57),
.Y(n_227)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_64),
.B(n_414),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_74),
.B(n_80),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_65),
.A2(n_174),
.B(n_177),
.Y(n_173)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_73),
.Y(n_349)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_73),
.Y(n_364)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_73),
.Y(n_370)
);

AO21x2_ASAP7_75t_L g260 ( 
.A1(n_74),
.A2(n_261),
.B(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_84),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_75),
.B(n_233),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_75),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_76),
.Y(n_382)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_77),
.Y(n_232)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_80),
.B(n_344),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_131),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_88),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_107),
.B(n_123),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_90),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_108),
.B(n_117),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_100),
.B2(n_104),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_107),
.B(n_123),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_111),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_117),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_123),
.Y(n_210)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_163),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_143),
.B(n_255),
.Y(n_309)
);

NOR2x1p5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_156),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B1(n_151),
.B2(n_154),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

AO22x2_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_163),
.B(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_171),
.B(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_201),
.C(n_206),
.Y(n_171)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_172),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_173),
.B(n_178),
.Y(n_318)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_177),
.B(n_381),
.Y(n_380)
);

OAI31xp33_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.A3(n_186),
.B(n_189),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B(n_198),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_201),
.B(n_207),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_254),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_209),
.B(n_213),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2x1_ASAP7_75t_L g313 ( 
.A(n_212),
.B(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2x2_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_229),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_228),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

AND2x4_ASAP7_75t_SL g343 ( 
.A(n_230),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_235),
.Y(n_347)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx4f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_269),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_259),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

OAI21x1_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2x2_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_260),
.A2(n_291),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_405),
.B(n_424),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_320),
.B(n_404),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_306),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_278),
.B(n_306),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_290),
.C(n_298),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_280),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_284),
.C(n_289),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_286),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_298),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_317),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_307),
.B(n_318),
.C(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_308),
.B(n_311),
.C(n_315),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

OAI21x1_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_336),
.B(n_403),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_333),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_333),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.C(n_329),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_352),
.B(n_402),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_350),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_338),
.B(n_350),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.C(n_342),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_378),
.B(n_401),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_357),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_377),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_384),
.B(n_400),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_383),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_390),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_388),
.B(n_399),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_387),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_398),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_419),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_426),
.Y(n_425)
);

NAND2x1_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_417),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_417),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.C(n_415),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_416),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_422),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.Y(n_424)
);


endmodule