module fake_jpeg_3891_n_143 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_18),
.C(n_13),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_11),
.B1(n_18),
.B2(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_16),
.B1(n_10),
.B2(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_28),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_23),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_29),
.C(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_40),
.C(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_60),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_40),
.B1(n_47),
.B2(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_72),
.B1(n_50),
.B2(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_49),
.B1(n_39),
.B2(n_30),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_39),
.B1(n_30),
.B2(n_44),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_22),
.B1(n_37),
.B2(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_83),
.C(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_56),
.B(n_55),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_39),
.B(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_64),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_54),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_89),
.B(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_67),
.B1(n_69),
.B2(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_16),
.B1(n_10),
.B2(n_14),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_92),
.C(n_77),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_73),
.B(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_25),
.B(n_11),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_52),
.B1(n_51),
.B2(n_22),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_58),
.B(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_34),
.B1(n_36),
.B2(n_75),
.C(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_100),
.C(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_75),
.C(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_34),
.C(n_15),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_95),
.C(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_20),
.C(n_16),
.Y(n_114)
);

AOI31xp67_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_87),
.A3(n_93),
.B(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_104),
.B(n_86),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_116),
.B(n_19),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.C(n_15),
.Y(n_119)
);

AOI31xp67_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_20),
.A3(n_10),
.B(n_15),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_15),
.B(n_19),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_108),
.B1(n_106),
.B2(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_124),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_19),
.C(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_0),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_110),
.B(n_2),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_6),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_134),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_3),
.B(n_4),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_4),
.B(n_6),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_3),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_3),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_133),
.B(n_7),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_140),
.B1(n_7),
.B2(n_8),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_9),
.Y(n_143)
);


endmodule