module fake_ariane_818_n_864 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_864);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_864;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_779;
wire n_754;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_99),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_59),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_89),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_100),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_70),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_L g206 ( 
.A(n_105),
.B(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_74),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_20),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_56),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_50),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_83),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_94),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_15),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_66),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_84),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_87),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_77),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_109),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_25),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_150),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_8),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_174),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_44),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_91),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_64),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_30),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_97),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_204),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_23),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_211),
.B(n_1),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_194),
.B(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_219),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_203),
.A2(n_92),
.B(n_180),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_202),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_197),
.B(n_3),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_211),
.B(n_3),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_239),
.B(n_4),
.Y(n_278)
);

OAI22x1_ASAP7_75t_SL g279 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_5),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_204),
.A2(n_220),
.B1(n_216),
.B2(n_251),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_209),
.A2(n_96),
.B(n_179),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_7),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_225),
.B(n_8),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_220),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_9),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_224),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_298)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_193),
.Y(n_302)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_274),
.B(n_193),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_294),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_217),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

AND3x2_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_237),
.C(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

BUFx6f_ASAP7_75t_SL g314 ( 
.A(n_270),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_286),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

NOR2x1p5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_281),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_286),
.B(n_217),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

NOR2x1p5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

NOR2x1p5_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_228),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_255),
.B(n_253),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_254),
.C(n_187),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_278),
.B(n_233),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_L g347 ( 
.A(n_262),
.B(n_266),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_278),
.B(n_252),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

BUFx4f_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g353 ( 
.A(n_264),
.B(n_206),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_344),
.A2(n_258),
.B1(n_283),
.B2(n_298),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_296),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_296),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_353),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_275),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_321),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_293),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_351),
.B(n_264),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_331),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_255),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_257),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_349),
.A2(n_290),
.B1(n_293),
.B2(n_277),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_257),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_261),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_304),
.B(n_289),
.C(n_288),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_297),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_351),
.B(n_277),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_262),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_261),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_269),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_262),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_269),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_277),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_314),
.A2(n_292),
.B1(n_299),
.B2(n_279),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_320),
.B(n_267),
.Y(n_391)
);

BUFx6f_ASAP7_75t_SL g392 ( 
.A(n_340),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_314),
.A2(n_308),
.B1(n_347),
.B2(n_292),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_273),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_299),
.B1(n_301),
.B2(n_300),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_323),
.B(n_299),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_276),
.B1(n_300),
.B2(n_295),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_309),
.B(n_284),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_319),
.B(n_186),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_303),
.A2(n_287),
.B1(n_295),
.B2(n_226),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_306),
.B(n_287),
.Y(n_408)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_303),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_307),
.A2(n_262),
.B1(n_285),
.B2(n_271),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_312),
.B(n_188),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_307),
.B(n_189),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_311),
.B(n_316),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_311),
.B(n_198),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_316),
.B(n_200),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_317),
.B(n_201),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_329),
.B(n_208),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_317),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_302),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_285),
.B(n_271),
.C(n_339),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_213),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_357),
.A2(n_222),
.B(n_221),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_306),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_345),
.B(n_342),
.C(n_339),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_366),
.A2(n_223),
.B1(n_229),
.B2(n_232),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_410),
.A2(n_262),
.B(n_342),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_234),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_238),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_391),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_240),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_379),
.A2(n_345),
.B(n_337),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_12),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_366),
.B(n_396),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_244),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_379),
.A2(n_335),
.B(n_334),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_388),
.A2(n_335),
.B(n_334),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_361),
.B(n_249),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_360),
.A2(n_333),
.B(n_330),
.C(n_328),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_405),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_388),
.A2(n_333),
.B(n_330),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_324),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_380),
.A2(n_328),
.B(n_327),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_395),
.A2(n_324),
.B1(n_327),
.B2(n_15),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_374),
.A2(n_371),
.B(n_369),
.Y(n_451)
);

NOR3xp33_ASAP7_75t_L g452 ( 
.A(n_355),
.B(n_13),
.C(n_14),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_407),
.B(n_329),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_397),
.B(n_329),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_329),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_400),
.B(n_13),
.Y(n_456)
);

AO21x1_ASAP7_75t_L g457 ( 
.A1(n_385),
.A2(n_104),
.B(n_177),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_373),
.A2(n_102),
.B(n_175),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_14),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_375),
.B(n_399),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_24),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_355),
.B(n_16),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_364),
.B(n_16),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_376),
.B(n_17),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_383),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_398),
.A2(n_362),
.B(n_367),
.C(n_370),
.Y(n_468)
);

BUFx4f_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_384),
.A2(n_107),
.B(n_173),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_402),
.A2(n_106),
.B(n_172),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_381),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_404),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_382),
.B(n_21),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_410),
.A2(n_22),
.B(n_28),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_362),
.A2(n_111),
.B(n_29),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_387),
.B(n_404),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_406),
.A2(n_112),
.B(n_31),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_413),
.A2(n_113),
.B(n_32),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_416),
.A2(n_114),
.B(n_33),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_367),
.B(n_22),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_370),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_417),
.A2(n_34),
.B(n_35),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

O2A1O1Ixp5_ASAP7_75t_L g485 ( 
.A1(n_421),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_485)
);

AO21x1_ASAP7_75t_L g486 ( 
.A1(n_414),
.A2(n_421),
.B(n_422),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_L g487 ( 
.A1(n_386),
.A2(n_40),
.B(n_41),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_390),
.B(n_42),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g489 ( 
.A(n_389),
.B(n_43),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_389),
.B(n_45),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_394),
.B(n_47),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_394),
.A2(n_48),
.B(n_49),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_SL g493 ( 
.A(n_411),
.B(n_51),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_411),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_449),
.A2(n_420),
.B(n_419),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_415),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_431),
.A2(n_420),
.B(n_419),
.Y(n_497)
);

INVx6_ASAP7_75t_SL g498 ( 
.A(n_448),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_440),
.B(n_448),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_431),
.A2(n_414),
.B(n_55),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

AOI221x1_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.C(n_60),
.Y(n_502)
);

AOI222xp33_ASAP7_75t_L g503 ( 
.A1(n_463),
.A2(n_392),
.B1(n_62),
.B2(n_65),
.C1(n_68),
.C2(n_69),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_61),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_72),
.Y(n_505)
);

NAND2x2_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_392),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_469),
.B(n_73),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_451),
.A2(n_436),
.B(n_447),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_458),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_443),
.A2(n_75),
.B(n_76),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_491),
.A2(n_78),
.B(n_79),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_475),
.A2(n_80),
.B(n_81),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_438),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_445),
.A2(n_82),
.B(n_86),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_427),
.B(n_88),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_432),
.A2(n_90),
.B(n_93),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_SL g519 ( 
.A(n_452),
.B(n_98),
.C(n_108),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_469),
.B(n_115),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_476),
.A2(n_116),
.B(n_117),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_472),
.B(n_118),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_442),
.A2(n_480),
.B(n_479),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_439),
.B(n_185),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_489),
.B(n_455),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_119),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_490),
.B(n_122),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_474),
.B(n_123),
.C(n_124),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_489),
.A2(n_126),
.B(n_127),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_430),
.A2(n_128),
.B1(n_131),
.B2(n_133),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_435),
.A2(n_134),
.B(n_135),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_425),
.B(n_136),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_424),
.A2(n_137),
.B(n_138),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_433),
.B(n_140),
.Y(n_535)
);

AOI21xp33_ASAP7_75t_L g536 ( 
.A1(n_450),
.A2(n_141),
.B(n_142),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_454),
.B(n_144),
.Y(n_537)
);

AO31x2_ASAP7_75t_L g538 ( 
.A1(n_486),
.A2(n_145),
.A3(n_146),
.B(n_147),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_459),
.A2(n_149),
.B(n_151),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_478),
.A2(n_152),
.B(n_153),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_485),
.A2(n_154),
.B(n_155),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_448),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_456),
.B(n_156),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_481),
.Y(n_544)
);

A2O1A1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_473),
.A2(n_157),
.B(n_159),
.C(n_162),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_462),
.A2(n_453),
.B(n_492),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_464),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

O2A1O1Ixp5_ASAP7_75t_L g549 ( 
.A1(n_460),
.A2(n_163),
.B(n_165),
.C(n_167),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_493),
.A2(n_168),
.B(n_170),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_468),
.A2(n_429),
.B(n_465),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_457),
.A2(n_470),
.B(n_471),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_441),
.A2(n_488),
.B(n_487),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_500),
.A2(n_513),
.B(n_497),
.Y(n_554)
);

NOR2x1_ASAP7_75t_R g555 ( 
.A(n_499),
.B(n_466),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_514),
.B(n_426),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_534),
.A2(n_505),
.B(n_551),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_501),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_498),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_524),
.A2(n_526),
.B(n_552),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_496),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_534),
.A2(n_508),
.B(n_546),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_495),
.A2(n_522),
.B(n_515),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_520),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_506),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_510),
.A2(n_541),
.B(n_530),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_505),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_511),
.A2(n_537),
.B(n_540),
.Y(n_574)
);

AO21x2_ASAP7_75t_L g575 ( 
.A1(n_551),
.A2(n_537),
.B(n_523),
.Y(n_575)
);

NOR2x1_ASAP7_75t_R g576 ( 
.A(n_507),
.B(n_521),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_539),
.A2(n_550),
.B(n_553),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_512),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_527),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_544),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_503),
.B(n_535),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_525),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_502),
.C(n_536),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_523),
.A2(n_543),
.B(n_533),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_543),
.A2(n_504),
.B(n_527),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_528),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_528),
.B(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_538),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_519),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_549),
.A2(n_517),
.B(n_532),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_529),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_529),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_501),
.B(n_463),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_548),
.B(n_294),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_500),
.A2(n_475),
.B(n_363),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_500),
.A2(n_524),
.B(n_526),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_559),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_560),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_580),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_581),
.A2(n_599),
.B1(n_583),
.B2(n_585),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_602),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_567),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_581),
.A2(n_596),
.B1(n_593),
.B2(n_589),
.Y(n_612)
);

OAI33xp33_ASAP7_75t_L g613 ( 
.A1(n_557),
.A2(n_603),
.A3(n_592),
.B1(n_569),
.B2(n_567),
.B3(n_588),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_602),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_604),
.B(n_556),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_563),
.A2(n_601),
.B(n_591),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_559),
.B(n_598),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_568),
.A2(n_577),
.B(n_563),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_598),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_573),
.A2(n_596),
.B1(n_589),
.B2(n_578),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_570),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_557),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

AO21x1_ASAP7_75t_SL g630 ( 
.A1(n_592),
.A2(n_597),
.B(n_584),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_562),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_604),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_588),
.Y(n_634)
);

BUFx2_ASAP7_75t_SL g635 ( 
.A(n_561),
.Y(n_635)
);

CKINVDCx6p67_ASAP7_75t_R g636 ( 
.A(n_562),
.Y(n_636)
);

BUFx8_ASAP7_75t_L g637 ( 
.A(n_571),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_566),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_561),
.B(n_578),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_578),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_571),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_579),
.B(n_596),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_595),
.B(n_558),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_600),
.B(n_590),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_565),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_582),
.A2(n_565),
.B1(n_594),
.B2(n_554),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_586),
.A2(n_558),
.B(n_575),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_612),
.B(n_558),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_644),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_608),
.A2(n_582),
.B1(n_575),
.B2(n_587),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_631),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_624),
.A2(n_582),
.B1(n_575),
.B2(n_587),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_644),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_611),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_565),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_644),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_623),
.B(n_601),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_624),
.A2(n_568),
.B1(n_574),
.B2(n_572),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_634),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_627),
.B(n_577),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_618),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_617),
.B(n_574),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_618),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_618),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_610),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_650),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_647),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_572),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_621),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_625),
.B(n_626),
.Y(n_673)
);

BUFx4f_ASAP7_75t_SL g674 ( 
.A(n_637),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_645),
.A2(n_642),
.B1(n_605),
.B2(n_635),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_639),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_643),
.A2(n_609),
.B(n_638),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_607),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_607),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_650),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_646),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_637),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_630),
.B(n_640),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_628),
.B(n_629),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_610),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_610),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_648),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_648),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_614),
.A2(n_632),
.B1(n_633),
.B2(n_649),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_616),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_616),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_SL g693 ( 
.A1(n_631),
.A2(n_636),
.B(n_613),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_615),
.B(n_620),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_622),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_614),
.B(n_616),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_613),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_614),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_641),
.B(n_612),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_612),
.B(n_611),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_612),
.B(n_611),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_608),
.A2(n_581),
.B1(n_463),
.B2(n_585),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_670),
.B(n_658),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_676),
.B(n_702),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_664),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_674),
.B(n_677),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_702),
.B(n_670),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_670),
.B(n_672),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_670),
.B(n_658),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_700),
.A2(n_701),
.B1(n_699),
.B2(n_697),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_652),
.B(n_659),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_664),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_689),
.B(n_697),
.C(n_653),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_693),
.B(n_675),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_672),
.B(n_662),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_664),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_700),
.B(n_701),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_688),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_652),
.B(n_659),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_657),
.B(n_662),
.Y(n_722)
);

OAI222xp33_ASAP7_75t_L g723 ( 
.A1(n_699),
.A2(n_651),
.B1(n_681),
.B2(n_696),
.C1(n_673),
.C2(n_678),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_652),
.B(n_659),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_698),
.B(n_683),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_652),
.B(n_659),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_656),
.B(n_687),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_657),
.B(n_687),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_681),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_687),
.B(n_665),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_665),
.B(n_671),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_673),
.B(n_660),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_684),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_651),
.A2(n_691),
.B1(n_694),
.B2(n_679),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_684),
.B(n_694),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_666),
.B(n_667),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_667),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_667),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_683),
.B(n_685),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_738),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_706),
.B(n_685),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_703),
.B(n_655),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_741),
.B(n_692),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_703),
.B(n_690),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_741),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_738),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_722),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_713),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_709),
.B(n_690),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_741),
.Y(n_752)
);

AND2x4_ASAP7_75t_SL g753 ( 
.A(n_711),
.B(n_692),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_713),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_728),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_718),
.B(n_669),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_721),
.B(n_685),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_719),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_709),
.B(n_695),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_719),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_718),
.B(n_732),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_708),
.B(n_680),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_732),
.B(n_695),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_724),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_729),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_711),
.B(n_692),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_730),
.B(n_695),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_734),
.B(n_686),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_711),
.B(n_692),
.Y(n_771)
);

NAND2x1_ASAP7_75t_L g772 ( 
.A(n_711),
.B(n_690),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_730),
.B(n_727),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_727),
.B(n_661),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_715),
.B(n_698),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_750),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_761),
.B(n_773),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_761),
.B(n_726),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_768),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_755),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_768),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_750),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_773),
.B(n_726),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_756),
.B(n_733),
.Y(n_784)
);

NAND2x1_ASAP7_75t_L g785 ( 
.A(n_765),
.B(n_721),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_749),
.B(n_707),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_758),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_743),
.B(n_698),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_747),
.B(n_720),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_758),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_747),
.B(n_720),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_762),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_764),
.B(n_724),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_764),
.B(n_736),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_752),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_756),
.B(n_716),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_742),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_762),
.B(n_710),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_714),
.B1(n_744),
.B2(n_704),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_765),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_776),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_782),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_777),
.A2(n_714),
.B1(n_775),
.B2(n_744),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_786),
.A2(n_752),
.B1(n_698),
.B2(n_691),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_793),
.B(n_765),
.Y(n_805)
);

OAI21xp33_ASAP7_75t_L g806 ( 
.A1(n_780),
.A2(n_774),
.B(n_770),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_795),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_779),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_787),
.Y(n_809)
);

AOI22x1_ASAP7_75t_SL g810 ( 
.A1(n_807),
.A2(n_654),
.B1(n_682),
.B2(n_792),
.Y(n_810)
);

OAI222xp33_ASAP7_75t_L g811 ( 
.A1(n_799),
.A2(n_784),
.B1(n_796),
.B2(n_785),
.C1(n_774),
.C2(n_794),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_808),
.Y(n_812)
);

AOI222xp33_ASAP7_75t_L g813 ( 
.A1(n_803),
.A2(n_806),
.B1(n_723),
.B2(n_804),
.C1(n_797),
.C2(n_801),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_803),
.A2(n_788),
.B(n_785),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_L g815 ( 
.A1(n_802),
.A2(n_784),
.B1(n_796),
.B2(n_797),
.C(n_790),
.Y(n_815)
);

AO22x1_ASAP7_75t_L g816 ( 
.A1(n_807),
.A2(n_745),
.B1(n_795),
.B2(n_771),
.Y(n_816)
);

OA22x2_ASAP7_75t_L g817 ( 
.A1(n_814),
.A2(n_800),
.B1(n_809),
.B2(n_805),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_814),
.A2(n_757),
.B(n_682),
.Y(n_818)
);

OAI221xp5_ASAP7_75t_L g819 ( 
.A1(n_813),
.A2(n_763),
.B1(n_766),
.B2(n_781),
.C(n_779),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_815),
.Y(n_820)
);

OAI222xp33_ASAP7_75t_L g821 ( 
.A1(n_810),
.A2(n_811),
.B1(n_812),
.B2(n_816),
.C1(n_742),
.C2(n_748),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_815),
.Y(n_822)
);

AOI221xp5_ASAP7_75t_SL g823 ( 
.A1(n_814),
.A2(n_791),
.B1(n_789),
.B2(n_778),
.C(n_783),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_821),
.A2(n_819),
.B(n_818),
.Y(n_824)
);

NAND4xp25_ASAP7_75t_L g825 ( 
.A(n_823),
.B(n_725),
.C(n_778),
.D(n_760),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_SL g826 ( 
.A1(n_818),
.A2(n_757),
.B(n_791),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_820),
.B(n_754),
.C(n_772),
.Y(n_827)
);

NAND4xp25_ASAP7_75t_L g828 ( 
.A(n_824),
.B(n_822),
.C(n_817),
.D(n_789),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_827),
.A2(n_757),
.B(n_783),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_826),
.B(n_772),
.C(n_737),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_828),
.B(n_825),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_830),
.A2(n_698),
.B1(n_745),
.B2(n_781),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_SL g833 ( 
.A(n_829),
.B(n_793),
.C(n_735),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_829),
.B(n_751),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_833),
.A2(n_745),
.B1(n_769),
.B2(n_767),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_834),
.B(n_737),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_832),
.B(n_759),
.Y(n_838)
);

NOR2x1_ASAP7_75t_L g839 ( 
.A(n_831),
.B(n_771),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_835),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_838),
.B(n_759),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_839),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_837),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_836),
.A2(n_748),
.B1(n_767),
.B2(n_771),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_835),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_751),
.B1(n_746),
.B2(n_728),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_842),
.A2(n_739),
.B1(n_668),
.B2(n_740),
.C(n_731),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_845),
.A2(n_769),
.B1(n_767),
.B2(n_746),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_843),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_841),
.Y(n_850)
);

XNOR2x1_ASAP7_75t_L g851 ( 
.A(n_849),
.B(n_844),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_850),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

AOI21xp33_ASAP7_75t_L g854 ( 
.A1(n_846),
.A2(n_844),
.B(n_739),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_853),
.A2(n_848),
.B1(n_740),
.B2(n_717),
.C(n_731),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_724),
.B(n_753),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_852),
.A2(n_668),
.B(n_740),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_854),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_858),
.A2(n_668),
.B1(n_740),
.B2(n_753),
.Y(n_859)
);

OAI21x1_ASAP7_75t_SL g860 ( 
.A1(n_856),
.A2(n_712),
.B(n_731),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_859),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_861),
.B(n_857),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_862),
.B(n_860),
.Y(n_863)
);

AOI211xp5_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_855),
.B(n_712),
.C(n_717),
.Y(n_864)
);


endmodule