module fake_jpeg_15333_n_393 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_41),
.B(n_50),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_26),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_28),
.B1(n_23),
.B2(n_4),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_19),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_26),
.B1(n_15),
.B2(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_69),
.A2(n_76),
.B1(n_90),
.B2(n_103),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_20),
.C(n_29),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_78),
.Y(n_127)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_26),
.B1(n_15),
.B2(n_17),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_25),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_80),
.B(n_86),
.Y(n_159)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_99),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_28),
.B1(n_17),
.B2(n_23),
.Y(n_90)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_16),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_28),
.B1(n_37),
.B2(n_36),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_16),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_37),
.Y(n_110)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_38),
.B(n_36),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_156)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_123),
.B(n_151),
.Y(n_214)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_124),
.B(n_129),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_82),
.A2(n_64),
.B1(n_56),
.B2(n_34),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_141),
.Y(n_205)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_142),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_29),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_155),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_69),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_123),
.B1(n_127),
.B2(n_165),
.Y(n_182)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_5),
.B(n_6),
.Y(n_179)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_105),
.B(n_29),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_162),
.B1(n_164),
.B2(n_101),
.Y(n_187)
);

BUFx12f_ASAP7_75t_SL g157 ( 
.A(n_73),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_161),
.B(n_159),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_169),
.Y(n_193)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

OR2x2_ASAP7_75t_SL g161 ( 
.A(n_85),
.B(n_30),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_90),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_76),
.B(n_19),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_89),
.A2(n_35),
.B1(n_19),
.B2(n_29),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_79),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_72),
.B(n_40),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_142),
.C(n_145),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_119),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_98),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_152),
.B(n_138),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_3),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_178),
.A2(n_183),
.B(n_199),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_179),
.A2(n_182),
.B(n_140),
.C(n_146),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_5),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_29),
.C(n_77),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_209),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_187),
.A2(n_197),
.B1(n_204),
.B2(n_179),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_212),
.B1(n_151),
.B2(n_150),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_84),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_207),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_68),
.B1(n_83),
.B2(n_107),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_7),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_131),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_11),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_131),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_139),
.B(n_8),
.C(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_138),
.A2(n_11),
.B1(n_160),
.B2(n_137),
.Y(n_211)
);

OAI22x1_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_148),
.B1(n_130),
.B2(n_143),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_166),
.B1(n_121),
.B2(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_226),
.B(n_230),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_171),
.B(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_218),
.B(n_219),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_222),
.Y(n_275)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_231),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_225),
.A2(n_240),
.B(n_216),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_146),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_236),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_182),
.A2(n_130),
.B(n_148),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_235),
.A2(n_230),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_149),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_183),
.A2(n_199),
.B1(n_178),
.B2(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_244),
.B1(n_245),
.B2(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_207),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_250),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_191),
.A2(n_178),
.B(n_195),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_193),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_214),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_191),
.A2(n_212),
.B1(n_183),
.B2(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_200),
.A2(n_175),
.B1(n_210),
.B2(n_177),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_177),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_186),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_175),
.A2(n_176),
.B1(n_203),
.B2(n_198),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_209),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_180),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_206),
.A2(n_180),
.B1(n_181),
.B2(n_192),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_255),
.B1(n_249),
.B2(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_206),
.B1(n_190),
.B2(n_181),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_194),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_246),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_264),
.B(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_271),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_272),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_281),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_277),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_215),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_264),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_240),
.A2(n_234),
.B1(n_226),
.B2(n_224),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_284),
.B1(n_261),
.B2(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_229),
.B(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_285),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_289),
.B(n_258),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_224),
.B1(n_227),
.B2(n_244),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_260),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_292),
.C(n_303),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_250),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_237),
.B1(n_251),
.B2(n_222),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_293),
.A2(n_294),
.B1(n_269),
.B2(n_275),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_251),
.B1(n_232),
.B2(n_248),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_228),
.B1(n_263),
.B2(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_301),
.A2(n_302),
.B(n_312),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_280),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_309),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_316),
.B1(n_314),
.B2(n_295),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_260),
.C(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_258),
.B(n_289),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_277),
.A2(n_257),
.B1(n_281),
.B2(n_272),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_256),
.B(n_279),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_266),
.B1(n_267),
.B2(n_259),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_287),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_333),
.Y(n_345)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_328),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_307),
.B(n_309),
.CI(n_299),
.CON(n_328),
.SN(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_335),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_270),
.B1(n_288),
.B2(n_308),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_337),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_339),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_299),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_291),
.C(n_303),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_346),
.C(n_349),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_314),
.B1(n_302),
.B2(n_312),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_331),
.B1(n_338),
.B2(n_334),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_292),
.C(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_297),
.C(n_293),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_300),
.C(n_301),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_357),
.C(n_320),
.Y(n_366)
);

FAx1_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_302),
.CI(n_313),
.CON(n_352),
.SN(n_352)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_325),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_336),
.Y(n_353)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_335),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_330),
.C(n_321),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_362),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_365),
.B(n_369),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_333),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_364),
.C(n_366),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_326),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_323),
.C(n_320),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_370),
.C(n_357),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_323),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_373),
.B(n_364),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_350),
.C(n_345),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_361),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_368),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_376),
.A2(n_377),
.B(n_344),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_358),
.A2(n_342),
.B(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_380),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_381),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_374),
.A2(n_341),
.B1(n_355),
.B2(n_348),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_359),
.B(n_343),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_382),
.B(n_371),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_367),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_387),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_383),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_389),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_390),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_383),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_392),
.A2(n_380),
.B(n_318),
.C(n_352),
.Y(n_393)
);


endmodule