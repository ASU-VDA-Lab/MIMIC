module real_jpeg_11408_n_16 (n_5, n_4, n_8, n_0, n_12, n_398, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_397, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_398;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_397;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_3),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_3),
.B(n_28),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_3),
.B(n_51),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_39),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_31),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_106),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_28),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_5),
.B(n_39),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_5),
.B(n_44),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_25),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_28),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_6),
.B(n_93),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_6),
.B(n_31),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_6),
.B(n_51),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_6),
.B(n_39),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_6),
.B(n_44),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_7),
.B(n_51),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_7),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_7),
.B(n_39),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_28),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_51),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_10),
.B(n_25),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_10),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_10),
.B(n_39),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_12),
.B(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_106),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_93),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_12),
.B(n_25),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_12),
.B(n_28),
.Y(n_343)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_93),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_13),
.B(n_31),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_13),
.B(n_25),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_28),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_14),
.B(n_39),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_14),
.B(n_25),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_106),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_14),
.B(n_93),
.Y(n_206)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_116),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_20),
.B(n_77),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.C(n_53),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_22),
.B(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_36),
.C(n_40),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.C(n_30),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_24),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_55),
.C(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_24),
.A2(n_30),
.B1(n_61),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_24),
.A2(n_61),
.B1(n_107),
.B2(n_108),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_24),
.B(n_107),
.C(n_250),
.Y(n_270)
);

INVx5_ASAP7_75t_SL g146 ( 
.A(n_25),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_27),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_27),
.A2(n_81),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_27),
.B(n_288),
.C(n_291),
.Y(n_336)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_29),
.B(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_30),
.B(n_91),
.C(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_30),
.A2(n_84),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_30),
.B(n_198),
.C(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_30),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_32),
.B(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_32),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_32),
.B(n_42),
.Y(n_267)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_37),
.B(n_134),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_43),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_43),
.B(n_177),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_43),
.B(n_135),
.Y(n_327)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_46),
.A2(n_53),
.B1(n_54),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_47),
.B(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_55),
.A2(n_56),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.C(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_59),
.A2(n_60),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_60),
.B(n_96),
.C(n_262),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_76),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_87),
.C(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_65),
.A2(n_69),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_67),
.A2(n_68),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_68),
.B(n_301),
.C(n_303),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_111),
.C(n_112),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_78),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_97),
.C(n_101),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_79),
.B(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_86),
.C(n_90),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_87),
.B(n_88),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_89),
.B(n_132),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_103),
.C(n_109),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_92),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_91),
.A2(n_92),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_91),
.A2(n_92),
.B1(n_109),
.B2(n_358),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_92),
.B(n_158),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_92),
.B(n_341),
.C(n_343),
.Y(n_359)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_94),
.B(n_177),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_96),
.A2(n_259),
.B1(n_260),
.B2(n_263),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_96),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_96),
.A2(n_263),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_97),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_103),
.A2(n_104),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_105),
.B(n_137),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_105),
.A2(n_139),
.B1(n_205),
.B2(n_206),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_139),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_105),
.B(n_206),
.C(n_304),
.Y(n_341)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_109),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_111),
.Y(n_391)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_380),
.A3(n_388),
.B1(n_392),
.B2(n_393),
.C(n_397),
.Y(n_117)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_312),
.A3(n_346),
.B1(n_374),
.B2(n_379),
.C(n_398),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_253),
.C(n_307),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_224),
.B(n_252),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_192),
.B(n_223),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_161),
.B(n_191),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_124),
.B(n_140),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_136),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_143),
.B1(n_144),
.B2(n_152),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_188),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.CI(n_128),
.CON(n_125),
.SN(n_125)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_129),
.A2(n_130),
.B1(n_136),
.B2(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_134),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_146),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_153),
.B2(n_160),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_152),
.C(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_158),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_158),
.A2(n_159),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_158),
.B(n_275),
.C(n_278),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_185),
.B(n_190),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_174),
.B(n_184),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_209),
.B2(n_210),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_211),
.C(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_207),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_221),
.B2(n_222),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_220),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_217),
.C(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_226),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_242),
.B2(n_251),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_241),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_241),
.C(n_251),
.Y(n_308)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_237),
.B2(n_238),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_239),
.C(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_233),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.CI(n_236),
.CON(n_233),
.SN(n_233)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_242),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.CI(n_248),
.CON(n_242),
.SN(n_242)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_244),
.C(n_248),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B(n_247),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_254),
.A2(n_376),
.B(n_377),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_284),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_255),
.B(n_284),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_272),
.C(n_283),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_264),
.C(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_268),
.C(n_270),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_273),
.B1(n_283),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_280),
.C(n_282),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_306),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_295),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_295),
.C(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_293),
.C(n_294),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_308),
.B(n_309),
.Y(n_376)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_313),
.A2(n_375),
.B(n_378),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_314),
.B(n_315),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_345),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_318),
.C(n_345),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_337),
.B2(n_338),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_339),
.C(n_340),
.Y(n_373)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_329),
.B2(n_330),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_331),
.C(n_336),
.Y(n_352)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_325),
.C(n_327),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_335),
.B2(n_336),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_343),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_348),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_373),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_360),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_360),
.C(n_373),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_355),
.C(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_365),
.B2(n_366),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_367),
.C(n_372),
.Y(n_383)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_381),
.B(n_382),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_389),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_384),
.CI(n_387),
.CON(n_382),
.SN(n_382)
);


endmodule