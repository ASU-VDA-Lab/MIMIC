module fake_netlist_1_11358_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
NAND2xp33_ASAP7_75t_SL g16 ( .A(n_11), .B(n_9), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_1), .A2(n_5), .B(n_2), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_8), .B(n_3), .Y(n_18) );
AOI22xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_14), .Y(n_20) );
CKINVDCx12_ASAP7_75t_R g21 ( .A(n_19), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
OAI211xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_16), .B(n_13), .C(n_18), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_17), .B1(n_15), .B2(n_14), .Y(n_25) );
XNOR2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_0), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_26), .Y(n_27) );
CKINVDCx16_ASAP7_75t_R g28 ( .A(n_25), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AOI322xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_4), .A3(n_12), .B1(n_17), .B2(n_27), .C1(n_28), .C2(n_16), .Y(n_30) );
endmodule