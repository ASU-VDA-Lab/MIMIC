module fake_ibex_34_n_539 (n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_539);

input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_539;

wire n_151;
wire n_85;
wire n_507;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_86;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_134;
wire n_94;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_88;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_89;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_275;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_480;
wire n_416;
wire n_365;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_214;
wire n_238;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_318;
wire n_291;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_425;

INVx1_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_13),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_26),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_44),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_29),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_38),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_36),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_10),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_30),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_5),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_34),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_19),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_11),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_16),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_50),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_25),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_18),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_80),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_9),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_43),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_77),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_40),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_0),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_89),
.B(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

AOI22x1_ASAP7_75t_SL g169 ( 
.A1(n_86),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_87),
.B(n_3),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_91),
.B(n_7),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_107),
.B(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_7),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_8),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_56),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_125),
.A2(n_60),
.B(n_82),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_90),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_112),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_116),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_127),
.B(n_15),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_101),
.B(n_21),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_93),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_84),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_95),
.A2(n_24),
.B(n_32),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_165),
.B(n_164),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_104),
.Y(n_215)
);

OR2x6_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_111),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_148),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_145),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_152),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_103),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_128),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_105),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2x1p5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_106),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_182),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_154),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_120),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

NOR2x1p5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_146),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_206),
.B(n_142),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_206),
.B(n_139),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_156),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_147),
.C(n_124),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_198),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_212),
.B(n_210),
.Y(n_254)
);

CKINVDCx11_ASAP7_75t_R g255 ( 
.A(n_205),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_48),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_181),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_202),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_65),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_70),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_160),
.B(n_71),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_166),
.B(n_72),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_168),
.B(n_74),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

BUFx6f_ASAP7_75t_SL g273 ( 
.A(n_216),
.Y(n_273)
);

OR2x6_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_211),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_231),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_207),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_173),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_163),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_221),
.B(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_186),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_184),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_231),
.B(n_183),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_220),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_199),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

O2A1O1Ixp5_ASAP7_75t_L g297 ( 
.A1(n_213),
.A2(n_165),
.B(n_174),
.C(n_194),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_261),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_224),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_153),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_215),
.B(n_170),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_150),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_191),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_151),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_267),
.B(n_258),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_272),
.B1(n_178),
.B2(n_177),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_158),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_234),
.A2(n_169),
.B1(n_176),
.B2(n_177),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_149),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_223),
.A2(n_185),
.B(n_188),
.C(n_193),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_185),
.Y(n_317)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_250),
.A2(n_185),
.B1(n_188),
.B2(n_193),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_243),
.B(n_188),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_223),
.B(n_244),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_216),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_241),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_273),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_297),
.A2(n_228),
.B(n_230),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_277),
.A2(n_303),
.B(n_308),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_281),
.A2(n_218),
.B(n_226),
.C(n_265),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_277),
.A2(n_249),
.B(n_229),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_240),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_255),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_252),
.B(n_264),
.C(n_237),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_200),
.B(n_253),
.C(n_239),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_274),
.B1(n_307),
.B2(n_309),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_291),
.Y(n_349)
);

CKINVDCx11_ASAP7_75t_R g350 ( 
.A(n_274),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_274),
.A2(n_257),
.B1(n_245),
.B2(n_246),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_257),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_248),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_273),
.A2(n_260),
.B1(n_263),
.B2(n_270),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_287),
.B(n_293),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_247),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_247),
.B(n_312),
.C(n_278),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_347),
.A2(n_319),
.B1(n_321),
.B2(n_317),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_321),
.Y(n_364)
);

NOR2x1_ASAP7_75t_SL g365 ( 
.A(n_325),
.B(n_289),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_317),
.Y(n_366)
);

BUFx4f_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_316),
.B(n_315),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_320),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_344),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_356),
.B1(n_332),
.B2(n_360),
.Y(n_373)
);

OAI21x1_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_348),
.B(n_361),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_342),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_356),
.B1(n_335),
.B2(n_329),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_362),
.B1(n_357),
.B2(n_345),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_328),
.Y(n_379)
);

AO21x1_ASAP7_75t_L g380 ( 
.A1(n_333),
.A2(n_354),
.B(n_339),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

AO22x1_ASAP7_75t_L g383 ( 
.A1(n_325),
.A2(n_341),
.B1(n_324),
.B2(n_343),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_341),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_338),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_251),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_340),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_340),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_251),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_251),
.Y(n_393)
);

NAND2x1_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_356),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_347),
.A2(n_298),
.B1(n_310),
.B2(n_311),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_SL g396 ( 
.A(n_327),
.B(n_222),
.C(n_286),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_331),
.A2(n_297),
.B(n_330),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_334),
.B(n_292),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_359),
.A2(n_282),
.B(n_347),
.C(n_281),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_331),
.A2(n_297),
.B(n_330),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_358),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_331),
.A2(n_297),
.B(n_330),
.Y(n_402)
);

AO31x2_ASAP7_75t_L g403 ( 
.A1(n_347),
.A2(n_362),
.A3(n_353),
.B(n_331),
.Y(n_403)
);

NOR2x1_ASAP7_75t_SL g404 ( 
.A(n_325),
.B(n_340),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

AO31x2_ASAP7_75t_L g406 ( 
.A1(n_347),
.A2(n_362),
.A3(n_353),
.B(n_331),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_251),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_251),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_251),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_325),
.B(n_340),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_334),
.B(n_292),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_351),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_379),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_388),
.A2(n_413),
.B1(n_405),
.B2(n_408),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_367),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_395),
.A2(n_366),
.B1(n_382),
.B2(n_370),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_414),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_389),
.Y(n_422)
);

NAND2x1p5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_367),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_378),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_395),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_404),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_393),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_409),
.B1(n_364),
.B2(n_368),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_371),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_397),
.A2(n_400),
.B(n_402),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_410),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_401),
.Y(n_434)
);

NOR3xp33_ASAP7_75t_SL g435 ( 
.A(n_363),
.B(n_376),
.C(n_377),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_369),
.A2(n_394),
.B(n_380),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_406),
.B(n_384),
.Y(n_438)
);

AO31x2_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_406),
.A3(n_365),
.B(n_386),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_385),
.A2(n_390),
.B1(n_391),
.B2(n_411),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_381),
.A2(n_403),
.B1(n_406),
.B2(n_383),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_388),
.A2(n_326),
.B1(n_413),
.B2(n_405),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

AO22x2_ASAP7_75t_L g445 ( 
.A1(n_395),
.A2(n_347),
.B1(n_373),
.B2(n_376),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_347),
.B1(n_298),
.B2(n_395),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_414),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_413),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_432),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_SL g451 ( 
.A1(n_421),
.A2(n_429),
.B(n_418),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_444),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_418),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_434),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_425),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

OAI22xp33_ASAP7_75t_L g464 ( 
.A1(n_443),
.A2(n_416),
.B1(n_427),
.B2(n_446),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_432),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_435),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_436),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_422),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_445),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_430),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_460),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_453),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_470),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_461),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_455),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_469),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_477),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_471),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_482),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_467),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_474),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_476),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_483),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_475),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_454),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_492),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_496),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_476),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_496),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_491),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_498),
.A2(n_451),
.B(n_464),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_497),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_499),
.A2(n_481),
.B(n_484),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_493),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_490),
.B(n_467),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_464),
.B(n_424),
.C(n_486),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_504),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_504),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_491),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_502),
.B(n_448),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_508),
.B(n_505),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_511),
.Y(n_518)
);

OAI211xp5_ASAP7_75t_L g519 ( 
.A1(n_513),
.A2(n_459),
.B(n_451),
.C(n_417),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_SL g520 ( 
.A(n_517),
.B(n_423),
.C(n_415),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_518),
.A2(n_509),
.B(n_514),
.Y(n_521)
);

NOR3x1_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_519),
.C(n_472),
.Y(n_522)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_463),
.Y(n_523)
);

NOR2x1_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_463),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_522),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_431),
.C(n_433),
.Y(n_526)
);

XNOR2x1_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_449),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_527),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_526),
.B1(n_507),
.B2(n_487),
.Y(n_529)
);

OAI22x1_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_420),
.B1(n_449),
.B2(n_465),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_428),
.B(n_463),
.Y(n_531)
);

XNOR2x2_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_440),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_532),
.B(n_530),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_531),
.A2(n_440),
.B(n_437),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_462),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_533),
.B(n_535),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_462),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_465),
.B(n_450),
.Y(n_539)
);


endmodule