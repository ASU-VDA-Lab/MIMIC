module fake_jpeg_26605_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

OR2x2_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_32),
.B1(n_27),
.B2(n_17),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_47),
.B1(n_39),
.B2(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_53),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_32),
.B1(n_22),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_37),
.B1(n_23),
.B2(n_18),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_16),
.B(n_36),
.C(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_39),
.B1(n_32),
.B2(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_74),
.B1(n_84),
.B2(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_85),
.B1(n_16),
.B2(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_73),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_39),
.B1(n_37),
.B2(n_34),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_81),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_26),
.B1(n_18),
.B2(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_96),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_109),
.B1(n_48),
.B2(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_45),
.B1(n_62),
.B2(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_17),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_53),
.C(n_43),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_36),
.C(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_110),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_57),
.B(n_55),
.C(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_25),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_116),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_80),
.B(n_82),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_118),
.B(n_121),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_135),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_67),
.B(n_19),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_124),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_70),
.B(n_74),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_109),
.B1(n_101),
.B2(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_74),
.B(n_0),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_103),
.B(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_130),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_133),
.B1(n_108),
.B2(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_114),
.Y(n_163)
);

OAI22x1_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_109),
.B1(n_97),
.B2(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_99),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_142),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_141),
.B1(n_131),
.B2(n_87),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_133),
.A2(n_106),
.B1(n_96),
.B2(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_103),
.C(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_156),
.C(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_151),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_24),
.B(n_21),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_93),
.C(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_55),
.B1(n_57),
.B2(n_19),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_117),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_135),
.B1(n_112),
.B2(n_87),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_93),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_20),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_138),
.C(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_186),
.C(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_171),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_172),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_125),
.B(n_119),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_183),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_185),
.B1(n_145),
.B2(n_144),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_95),
.B1(n_89),
.B2(n_74),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_178),
.B1(n_181),
.B2(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_75),
.B1(n_77),
.B2(n_69),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_150),
.B1(n_137),
.B2(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_57),
.B1(n_20),
.B2(n_21),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_24),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_29),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_71),
.C(n_36),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_22),
.B(n_24),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_138),
.B(n_31),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_0),
.C(n_31),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_1),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_204),
.B1(n_177),
.B2(n_29),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_164),
.C(n_146),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.C(n_200),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_155),
.C(n_151),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_178),
.B1(n_180),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_210),
.B1(n_179),
.B2(n_187),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.C(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_159),
.B1(n_153),
.B2(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_160),
.C(n_36),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_30),
.C(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_206),
.B1(n_210),
.B2(n_207),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_188),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_200),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_223),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_192),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_198),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_235),
.C(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_234),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_193),
.C(n_196),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_222),
.B1(n_219),
.B2(n_224),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_214),
.B1(n_216),
.B2(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_217),
.B(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_245),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_238),
.B(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_3),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_3),
.C(n_4),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_229),
.C(n_236),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_14),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_256),
.C(n_247),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_230),
.B1(n_5),
.B2(n_6),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_7),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_252),
.A2(n_255),
.B(n_7),
.C(n_8),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_257),
.Y(n_261)
);

AOI211xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_248),
.Y(n_259)
);

NAND4xp25_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_243),
.C(n_244),
.D(n_246),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_9),
.B(n_10),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.B1(n_261),
.B2(n_10),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_253),
.B(n_246),
.C(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_266),
.B(n_9),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_9),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_10),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_267),
.C(n_11),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_11),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_12),
.Y(n_273)
);


endmodule