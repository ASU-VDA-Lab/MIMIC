module real_jpeg_24628_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_0),
.B(n_43),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_0),
.B(n_40),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_0),
.B(n_50),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_0),
.B(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_2),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_43),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_2),
.B(n_50),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_131),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_2),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_3),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_3),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_3),
.B(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_50),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_3),
.B(n_167),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_4),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_4),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_50),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_167),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx8_ASAP7_75t_SL g133 ( 
.A(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_8),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_9),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_36),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_40),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_50),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_9),
.B(n_167),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_61),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_43),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_10),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_10),
.B(n_40),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_10),
.B(n_50),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_10),
.B(n_329),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_11),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_11),
.B(n_61),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_11),
.B(n_43),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_11),
.B(n_36),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_11),
.B(n_40),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_11),
.B(n_50),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_11),
.B(n_131),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_11),
.B(n_329),
.Y(n_378)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_13),
.B(n_43),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_13),
.B(n_36),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_13),
.B(n_40),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_13),
.B(n_50),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_13),
.B(n_131),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_13),
.B(n_329),
.Y(n_365)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_16),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_50),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_16),
.B(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_16),
.B(n_167),
.Y(n_209)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_384),
.B(n_385),
.C(n_390),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_374),
.C(n_383),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_359),
.C(n_360),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_337),
.C(n_338),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_304),
.C(n_305),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_279),
.C(n_280),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_247),
.C(n_248),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_211),
.C(n_212),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_174),
.C(n_175),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_140),
.C(n_141),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_111),
.C(n_112),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_72),
.C(n_83),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_64),
.C(n_65),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_71),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_82),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_107),
.C(n_108),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.C(n_97),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.C(n_102),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_126),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_127),
.C(n_139),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_121),
.C(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_120),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_122),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.CI(n_125),
.CON(n_122),
.SN(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_139),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_137),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_132),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_132),
.B(n_218),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_132),
.B(n_233),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.C(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_152),
.C(n_155),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_147),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.CI(n_150),
.CON(n_147),
.SN(n_147)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_164),
.C(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B(n_163),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_163),
.B(n_200),
.C(n_201),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_170),
.C(n_171),
.Y(n_195)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_168),
.Y(n_331)
);

INVx8_ASAP7_75t_L g389 ( 
.A(n_168),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_196),
.B2(n_210),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_197),
.C(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_180),
.C(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_183),
.B(n_233),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_193),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_243),
.C(n_244),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.CI(n_209),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_245),
.B2(n_246),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_237),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_237),
.C(n_245),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_225),
.C(n_226),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_236),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_227),
.Y(n_236)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_231),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_235),
.C(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_230),
.B(n_254),
.C(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_251),
.C(n_278),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_265),
.B2(n_278),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_260),
.C(n_261),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_257),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_258),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_SL g319 ( 
.A(n_257),
.B(n_284),
.C(n_287),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_261),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.CI(n_264),
.CON(n_261),
.SN(n_261)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_277),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_273),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_275),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_301),
.C(n_302),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_303),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_294),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_294),
.C(n_303),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_289),
.C(n_290),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_287),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_SL g348 ( 
.A(n_287),
.B(n_312),
.C(n_314),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_290),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.CI(n_293),
.CON(n_290),
.SN(n_290)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_308),
.C(n_321),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_320),
.B2(n_321),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_316),
.B2(n_317),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_318),
.C(n_319),
.Y(n_340)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_314),
.A2(n_315),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_353),
.C(n_354),
.Y(n_366)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_324),
.C(n_327),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_333),
.C(n_336),
.Y(n_346)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_335),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_341),
.C(n_358),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_348),
.C(n_349),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_361),
.C(n_363),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.CI(n_346),
.CON(n_343),
.SN(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_354),
.B2(n_355),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_352),
.A2(n_353),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_370),
.C(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_366),
.C(n_367),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_372),
.B2(n_373),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_370),
.A2(n_371),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g391 ( 
.A(n_371),
.B(n_378),
.C(n_381),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_372),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_377),
.C(n_382),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_381),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_381),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_388),
.Y(n_390)
);


endmodule