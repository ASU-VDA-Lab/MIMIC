module fake_jpeg_25087_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_152;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_18),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_40),
.B1(n_36),
.B2(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_51),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_20),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_28),
.B(n_33),
.C(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_40),
.B1(n_16),
.B2(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_74),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_18),
.B1(n_26),
.B2(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_27),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_26),
.B1(n_39),
.B2(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_40),
.B1(n_39),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_30),
.B1(n_38),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_51),
.B1(n_58),
.B2(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_38),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_28),
.B1(n_17),
.B2(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_17),
.B(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_35),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_28),
.A3(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_84),
.B(n_87),
.C(n_81),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_63),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_35),
.C(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_85),
.C(n_62),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_60),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_29),
.B1(n_17),
.B2(n_30),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_117),
.B1(n_65),
.B2(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_63),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_21),
.B1(n_35),
.B2(n_22),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_76),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_22),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_123),
.Y(n_158)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_132),
.B1(n_146),
.B2(n_115),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_125),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_73),
.B1(n_89),
.B2(n_63),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_131),
.B1(n_145),
.B2(n_95),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_139),
.B(n_107),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_71),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_88),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_89),
.B1(n_63),
.B2(n_62),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_141),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_140),
.Y(n_164)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_93),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_83),
.B1(n_76),
.B2(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_95),
.B1(n_117),
.B2(n_118),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_61),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_110),
.C(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_76),
.B1(n_90),
.B2(n_2),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_151),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_133),
.B(n_128),
.C(n_137),
.D(n_104),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_0),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_108),
.B(n_113),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_173),
.B1(n_106),
.B2(n_96),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_172),
.B1(n_154),
.B2(n_148),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_176),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_123),
.B(n_124),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_168),
.B(n_169),
.Y(n_199)
);

BUFx12f_ASAP7_75t_SL g163 ( 
.A(n_119),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_110),
.C(n_100),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_178),
.B(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_97),
.B(n_61),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_136),
.B1(n_142),
.B2(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_134),
.B1(n_143),
.B2(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_205),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_186),
.B1(n_196),
.B2(n_165),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_61),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_171),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_106),
.B1(n_96),
.B2(n_97),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_188),
.B(n_193),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_97),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_14),
.C(n_2),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_177),
.C(n_168),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_3),
.C(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_201),
.C(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_5),
.C(n_6),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_203),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_214),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_198),
.B1(n_191),
.B2(n_188),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_183),
.B1(n_187),
.B2(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_175),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_216),
.Y(n_232)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_166),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_154),
.B(n_149),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_155),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_151),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_159),
.B1(n_176),
.B2(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_231),
.B1(n_233),
.B2(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_170),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_241),
.B1(n_218),
.B2(n_214),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_209),
.A2(n_203),
.B1(n_199),
.B2(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_181),
.B1(n_201),
.B2(n_182),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_150),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_185),
.C(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_238),
.C(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_197),
.C(n_178),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_188),
.B1(n_192),
.B2(n_150),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_211),
.B1(n_217),
.B2(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_216),
.C(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_231),
.B1(n_233),
.B2(n_242),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_252),
.B1(n_256),
.B2(n_243),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_224),
.B1(n_192),
.B2(n_153),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_232),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_224),
.B1(n_190),
.B2(n_152),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_152),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_167),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_248),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_234),
.B(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_254),
.B1(n_249),
.B2(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_246),
.C(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_240),
.C(n_253),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_7),
.B(n_8),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_284),
.Y(n_288)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_262),
.A3(n_266),
.B1(n_269),
.B2(n_240),
.C1(n_261),
.C2(n_153),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_285),
.B1(n_276),
.B2(n_275),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_174),
.C2(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_174),
.C(n_10),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_289),
.C(n_290),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_9),
.B(n_10),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_281),
.C(n_10),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_288),
.C(n_11),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_291),
.C(n_11),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_9),
.B(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_12),
.B(n_289),
.Y(n_296)
);


endmodule