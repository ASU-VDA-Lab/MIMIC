module fake_jpeg_27324_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_44),
.B1(n_47),
.B2(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_20),
.B1(n_32),
.B2(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_34),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_27),
.B1(n_32),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_85)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_77),
.Y(n_99)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_86),
.B1(n_92),
.B2(n_57),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_84),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_39),
.B1(n_20),
.B2(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_91),
.B1(n_57),
.B2(n_67),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_39),
.B1(n_20),
.B2(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_93),
.Y(n_125)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_39),
.B(n_40),
.C(n_33),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_67),
.B1(n_50),
.B2(n_57),
.Y(n_90)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_62),
.B(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_29),
.B1(n_36),
.B2(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_24),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_43),
.C(n_38),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_46),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_38),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_25),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_121),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_127),
.B1(n_68),
.B2(n_88),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_74),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_26),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_66),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_60),
.B1(n_59),
.B2(n_43),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_91),
.B(n_26),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx10_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_147),
.B1(n_119),
.B2(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_68),
.B1(n_69),
.B2(n_97),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_43),
.B1(n_38),
.B2(n_37),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_155),
.B1(n_119),
.B2(n_111),
.Y(n_160)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_98),
.C(n_118),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_117),
.A3(n_108),
.B1(n_104),
.B2(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_144),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_99),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_139),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_174),
.B1(n_178),
.B2(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_99),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_133),
.B1(n_154),
.B2(n_147),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_105),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_122),
.B1(n_112),
.B2(n_114),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_182),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_123),
.B1(n_33),
.B2(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_123),
.B1(n_80),
.B2(n_76),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_145),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_197),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_157),
.B(n_23),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_194),
.B(n_208),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_214),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_131),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_137),
.C(n_37),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_215),
.C(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_148),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_152),
.Y(n_204)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_11),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_82),
.Y(n_207)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_23),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_152),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_24),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_156),
.C(n_164),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_165),
.Y(n_216)
);

NOR4xp25_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_171),
.C(n_170),
.D(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_24),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_185),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_208),
.B1(n_211),
.B2(n_188),
.Y(n_258)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_229),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_193),
.B1(n_197),
.B2(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_34),
.C(n_29),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_214),
.C(n_201),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_29),
.B1(n_0),
.B2(n_2),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_193),
.B1(n_191),
.B2(n_202),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_233),
.C(n_224),
.Y(n_266)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_202),
.B1(n_191),
.B2(n_192),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_262),
.B1(n_231),
.B2(n_239),
.Y(n_273)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_196),
.C(n_218),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_263),
.C(n_244),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_259),
.B(n_219),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_205),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_260),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_227),
.A2(n_196),
.B1(n_0),
.B2(n_2),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_22),
.C(n_1),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_22),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_243),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_8),
.C(n_1),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_222),
.C(n_232),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_232),
.C(n_238),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_271),
.B(n_277),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_259),
.B(n_261),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_273),
.A2(n_265),
.B1(n_3),
.B2(n_5),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_231),
.C(n_227),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_230),
.C(n_236),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_230),
.C(n_1),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_9),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_298),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_277),
.B(n_278),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_251),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_299),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_245),
.B1(n_262),
.B2(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

BUFx12_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_269),
.C(n_3),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_303),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_8),
.C(n_3),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_10),
.B(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_312),
.C(n_294),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_11),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_6),
.C(n_7),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_300),
.B1(n_284),
.B2(n_309),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_318),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_319),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_304),
.A2(n_286),
.B(n_294),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_7),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_325),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_302),
.B(n_310),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_321),
.C(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_7),
.C(n_8),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_12),
.C(n_13),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_323),
.Y(n_334)
);

AOI311xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_331),
.A3(n_327),
.B(n_326),
.C(n_332),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_325),
.B(n_12),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_13),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_0),
.B(n_15),
.C(n_334),
.Y(n_339)
);


endmodule