module fake_jpeg_23187_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_16),
.B1(n_23),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_41),
.B1(n_50),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_18),
.B1(n_16),
.B2(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_48),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_25),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_52),
.C(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_21),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_21),
.B(n_15),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_28),
.B(n_20),
.C(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_70),
.B(n_43),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_0),
.C(n_1),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_54),
.B1(n_60),
.B2(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_67),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_43),
.B1(n_46),
.B2(n_42),
.Y(n_76)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_61),
.B(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_45),
.B1(n_24),
.B2(n_13),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_45),
.B1(n_20),
.B2(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_82),
.B1(n_56),
.B2(n_69),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_20),
.B1(n_27),
.B2(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_62),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_91),
.C(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_92),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_96),
.B(n_75),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_68),
.C(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR4xp25_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_63),
.C(n_55),
.D(n_62),
.Y(n_95)
);

NOR4xp25_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_97),
.C(n_85),
.D(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_109),
.B(n_110),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_71),
.C(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_105),
.C(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_75),
.C(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_94),
.B(n_86),
.Y(n_109)
);

AO221x1_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_73),
.B1(n_58),
.B2(n_20),
.C(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_117),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_107),
.B(n_110),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_107),
.B(n_105),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_77),
.C(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_27),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_123),
.B1(n_124),
.B2(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_109),
.B1(n_84),
.B2(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_67),
.B1(n_73),
.B2(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_4),
.Y(n_131)
);

AOI222xp33_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_115),
.C(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_121),
.B(n_120),
.Y(n_132)
);

AOI31xp67_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_4),
.A3(n_7),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_133),
.B(n_122),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_137),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_122),
.B(n_11),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_7),
.C(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_9),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_139),
.Y(n_141)
);


endmodule