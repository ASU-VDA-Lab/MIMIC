module fake_jpeg_31268_n_532 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_532);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_21),
.B(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_66),
.Y(n_150)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_0),
.C(n_1),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_72),
.B(n_20),
.C(n_37),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_96),
.Y(n_134)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_1),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_102),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_18),
.B(n_2),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_109),
.Y(n_129)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_43),
.B1(n_54),
.B2(n_53),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_113),
.A2(n_133),
.B1(n_157),
.B2(n_165),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_43),
.B1(n_82),
.B2(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_58),
.A2(n_22),
.B1(n_40),
.B2(n_54),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_143),
.B1(n_149),
.B2(n_161),
.Y(n_186)
);

BUFx16f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_28),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_62),
.A2(n_81),
.B1(n_102),
.B2(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_29),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_144),
.B(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_68),
.A2(n_22),
.B1(n_54),
.B2(n_50),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_19),
.C(n_46),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_155),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_69),
.B(n_37),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_56),
.A2(n_22),
.B1(n_50),
.B2(n_47),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_33),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_168),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_75),
.A2(n_50),
.B1(n_38),
.B2(n_47),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_83),
.A2(n_43),
.B1(n_53),
.B2(n_38),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_76),
.B(n_20),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_41),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_175),
.B(n_216),
.Y(n_257)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_114),
.A2(n_78),
.B1(n_55),
.B2(n_53),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_177),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_33),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_217),
.C(n_218),
.Y(n_232)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_181),
.Y(n_255)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_183),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_122),
.A2(n_86),
.B1(n_77),
.B2(n_90),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_185),
.A2(n_215),
.B1(n_163),
.B2(n_169),
.Y(n_251)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_187),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_29),
.B1(n_49),
.B2(n_46),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_192),
.Y(n_248)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_200),
.Y(n_261)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_89),
.B1(n_84),
.B2(n_50),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_203),
.B1(n_208),
.B2(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_125),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_109),
.B1(n_107),
.B2(n_87),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_206),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_139),
.A2(n_47),
.B1(n_42),
.B2(n_32),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_210),
.Y(n_241)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_213),
.Y(n_254)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_123),
.A2(n_49),
.B1(n_45),
.B2(n_41),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

NAND2xp67_ASAP7_75t_SL g217 ( 
.A(n_113),
.B(n_26),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_142),
.B(n_45),
.Y(n_218)
);

BUFx8_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_134),
.B(n_25),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_134),
.Y(n_235)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_130),
.A2(n_47),
.B1(n_42),
.B2(n_25),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_26),
.B1(n_19),
.B2(n_42),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_133),
.B1(n_157),
.B2(n_145),
.Y(n_250)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_145),
.B1(n_146),
.B2(n_117),
.Y(n_258)
);

OR2x4_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_116),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_230),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_226),
.A2(n_137),
.B1(n_163),
.B2(n_169),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_231),
.A2(n_251),
.B1(n_252),
.B2(n_256),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_235),
.B(n_184),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_166),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_246),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_150),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_240),
.B(n_26),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_186),
.B1(n_203),
.B2(n_137),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_250),
.B1(n_177),
.B2(n_201),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_130),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_150),
.B(n_114),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_175),
.B(n_141),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_260),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_204),
.B(n_141),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_189),
.B(n_123),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_185),
.A2(n_152),
.B(n_146),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_185),
.B(n_225),
.C(n_227),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_136),
.B1(n_162),
.B2(n_167),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_271),
.A2(n_282),
.B1(n_288),
.B2(n_290),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_274),
.B1(n_277),
.B2(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_185),
.B1(n_162),
.B2(n_167),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_251),
.B(n_243),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_276),
.B(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_197),
.B1(n_159),
.B2(n_195),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_279),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_280),
.B(n_300),
.Y(n_328)
);

BUFx24_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_180),
.B1(n_223),
.B2(n_214),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_176),
.B1(n_170),
.B2(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_211),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_292),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_170),
.B1(n_42),
.B2(n_216),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_198),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_248),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_268),
.A2(n_26),
.B1(n_219),
.B2(n_188),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_299),
.B1(n_243),
.B2(n_264),
.Y(n_323)
);

INVx11_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_268),
.A2(n_219),
.B1(n_26),
.B2(n_6),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_26),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_308),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_232),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_239),
.C(n_257),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_311),
.A2(n_321),
.B(n_234),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_251),
.B1(n_257),
.B2(n_245),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_312),
.A2(n_316),
.B1(n_287),
.B2(n_297),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_292),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_325),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_323),
.B(n_327),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_287),
.A2(n_251),
.B1(n_257),
.B2(n_253),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_265),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_278),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_243),
.B(n_237),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_323),
.A2(n_330),
.B1(n_273),
.B2(n_286),
.Y(n_340)
);

OAI221xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_235),
.B1(n_229),
.B2(n_241),
.C(n_239),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_272),
.A2(n_239),
.B1(n_236),
.B2(n_228),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_234),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_236),
.B1(n_255),
.B2(n_261),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_261),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_262),
.C(n_267),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_333),
.A2(n_334),
.B(n_308),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_286),
.B(n_280),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_306),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_338),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_348),
.B1(n_322),
.B2(n_309),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_302),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_345),
.B1(n_359),
.B2(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_289),
.B1(n_275),
.B2(n_270),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_300),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_347),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_312),
.A2(n_277),
.B1(n_291),
.B2(n_275),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_353),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_269),
.Y(n_350)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_351),
.B(n_352),
.Y(n_370)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_265),
.C(n_266),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_332),
.C(n_329),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_328),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_356),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_360),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_315),
.B1(n_330),
.B2(n_316),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_228),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_324),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_362),
.B(n_281),
.Y(n_381)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_381),
.C(n_382),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_368),
.B(n_391),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_335),
.B(n_331),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_369),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_384),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_374),
.A2(n_376),
.B1(n_378),
.B2(n_392),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_317),
.B1(n_309),
.B2(n_324),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_356),
.A2(n_317),
.B1(n_319),
.B2(n_326),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_333),
.A2(n_319),
.B(n_281),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_336),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_344),
.A2(n_281),
.B(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_380),
.B(n_388),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_262),
.C(n_293),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_279),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_298),
.B(n_279),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_385),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_389),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_351),
.A2(n_298),
.B(n_188),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_334),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_259),
.B1(n_267),
.B2(n_233),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_233),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_362),
.C(n_339),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_337),
.C(n_346),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_398),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_377),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_415),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_390),
.B(n_341),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_401),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_383),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_406),
.Y(n_443)
);

AO32x1_ASAP7_75t_L g405 ( 
.A1(n_364),
.A2(n_340),
.A3(n_350),
.B1(n_348),
.B2(n_342),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_405),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_354),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_362),
.Y(n_408)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_408),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_382),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_413),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_385),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_353),
.C(n_361),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_420),
.C(n_393),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_418),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_369),
.A2(n_343),
.B1(n_358),
.B2(n_8),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_419),
.A2(n_422),
.B1(n_372),
.B2(n_365),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_358),
.C(n_247),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_358),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_366),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_380),
.B(n_188),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_434),
.C(n_413),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_370),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_428),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_370),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_368),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_445),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_SL g430 ( 
.A(n_402),
.B(n_388),
.C(n_385),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_430),
.A2(n_403),
.B(n_414),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_367),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_432),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_420),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_427),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_376),
.C(n_379),
.Y(n_434)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_400),
.A2(n_371),
.B1(n_375),
.B2(n_387),
.Y(n_441)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_375),
.B1(n_387),
.B2(n_374),
.Y(n_445)
);

FAx1_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_394),
.CI(n_405),
.CON(n_446),
.SN(n_446)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_461),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_247),
.C(n_5),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_401),
.B(n_407),
.Y(n_450)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_454),
.A2(n_463),
.B(n_444),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_412),
.C(n_416),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_460),
.C(n_432),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_405),
.B1(n_410),
.B2(n_414),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_456),
.A2(n_457),
.B1(n_434),
.B2(n_392),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_412),
.B1(n_398),
.B2(n_418),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_418),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_462),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_L g463 ( 
.A1(n_440),
.A2(n_397),
.B(n_409),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_436),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_453),
.A2(n_444),
.B1(n_458),
.B2(n_442),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_471),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_480),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_475),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_462),
.A2(n_397),
.B1(n_445),
.B2(n_404),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_478),
.B1(n_452),
.B2(n_446),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_16),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_378),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_431),
.C(n_433),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_477),
.C(n_481),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_428),
.C(n_426),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_404),
.B1(n_421),
.B2(n_365),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_372),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_247),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_452),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_466),
.B(n_471),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_463),
.B1(n_459),
.B2(n_460),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_487),
.B(n_491),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_476),
.B(n_459),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_489),
.Y(n_506)
);

XOR2x1_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_451),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_490),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_451),
.C(n_247),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_484),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_480),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_472),
.A2(n_3),
.B(n_5),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_495),
.B(n_493),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_8),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_467),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_477),
.C(n_465),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_498),
.B(n_501),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_494),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_467),
.C(n_473),
.Y(n_501)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_504),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_8),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_505),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_10),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_490),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_492),
.A2(n_10),
.B(n_12),
.Y(n_508)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_508),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_489),
.Y(n_510)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_513),
.Y(n_521)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_511),
.A2(n_509),
.B(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_520),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_497),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_497),
.C(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_516),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_525),
.C(n_519),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_513),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g528 ( 
.A1(n_526),
.A2(n_527),
.B(n_500),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_524),
.A2(n_519),
.B(n_515),
.C(n_510),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_10),
.B(n_13),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_13),
.B(n_14),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_15),
.C(n_13),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_14),
.B1(n_15),
.B2(n_469),
.Y(n_532)
);


endmodule