module fake_jpeg_26318_n_311 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_19),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_46),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_25),
.B1(n_28),
.B2(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_54),
.B1(n_57),
.B2(n_60),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_47),
.B1(n_31),
.B2(n_33),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_45),
.B1(n_44),
.B2(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_63),
.B1(n_44),
.B2(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_21),
.B1(n_17),
.B2(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_40),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_38),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_86),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_93),
.B(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_97),
.B(n_101),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_55),
.B1(n_63),
.B2(n_50),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_98),
.A2(n_116),
.B1(n_41),
.B2(n_55),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_86),
.B1(n_79),
.B2(n_80),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_65),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_64),
.B1(n_67),
.B2(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_61),
.B1(n_92),
.B2(n_56),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_65),
.C(n_44),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_32),
.C(n_36),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_38),
.A3(n_46),
.B1(n_65),
.B2(n_43),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_43),
.A3(n_42),
.B1(n_91),
.B2(n_75),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_107),
.Y(n_124)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_64),
.B1(n_84),
.B2(n_67),
.Y(n_119)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_112),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_118),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_46),
.B1(n_44),
.B2(n_51),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_120),
.A2(n_123),
.B(n_125),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_71),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_127),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_79),
.B(n_77),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_100),
.B(n_94),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_132),
.B(n_135),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_134),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_87),
.B1(n_91),
.B2(n_57),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_32),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_41),
.B1(n_55),
.B2(n_37),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_98),
.B1(n_109),
.B2(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_148),
.B1(n_102),
.B2(n_108),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_109),
.B1(n_98),
.B2(n_105),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_147),
.B1(n_108),
.B2(n_111),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_101),
.B(n_96),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_32),
.B(n_24),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_98),
.A2(n_41),
.B1(n_37),
.B2(n_48),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_37),
.B1(n_56),
.B2(n_17),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_118),
.B1(n_96),
.B2(n_99),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_157),
.B1(n_184),
.B2(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_155),
.B(n_170),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_148),
.B1(n_140),
.B2(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_48),
.B1(n_37),
.B2(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_22),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_22),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_22),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_23),
.Y(n_176)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_37),
.B1(n_68),
.B2(n_16),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_12),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_23),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_169),
.B(n_146),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_68),
.B1(n_18),
.B2(n_16),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_192),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_183),
.B1(n_179),
.B2(n_158),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_134),
.C(n_130),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_193),
.C(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_150),
.C(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_196),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_125),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_156),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_153),
.B1(n_177),
.B2(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_36),
.C(n_12),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_23),
.B(n_24),
.Y(n_209)
);

AND3x1_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_183),
.C(n_161),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_165),
.B1(n_160),
.B2(n_157),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_184),
.B1(n_178),
.B2(n_175),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_173),
.B1(n_168),
.B2(n_166),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_230),
.B1(n_207),
.B2(n_199),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_229),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_224),
.B1(n_231),
.B2(n_188),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_180),
.B(n_166),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_193),
.C(n_197),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_227),
.C(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_181),
.C(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_200),
.B1(n_195),
.B2(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_153),
.B1(n_177),
.B2(n_68),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_12),
.C(n_18),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_247),
.B1(n_248),
.B2(n_6),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_227),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_198),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_201),
.B1(n_210),
.B2(n_192),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_7),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_205),
.B1(n_208),
.B2(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_203),
.C(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_189),
.C(n_206),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_194),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_231),
.B1(n_223),
.B2(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_218),
.B1(n_199),
.B2(n_232),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_209),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_253),
.B(n_246),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_216),
.B(n_212),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_250),
.B(n_238),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_189),
.B1(n_217),
.B2(n_18),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_260),
.B1(n_7),
.B2(n_10),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_24),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_18),
.C(n_16),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_24),
.C(n_1),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_24),
.C(n_1),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_5),
.B1(n_10),
.B2(n_2),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_238),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_240),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_275),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_6),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_11),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_251),
.B1(n_254),
.B2(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_289),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_262),
.B1(n_259),
.B2(n_3),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_5),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_7),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_8),
.B(n_10),
.C(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_271),
.C(n_276),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_271),
.B(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_281),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_3),
.Y(n_299)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_296),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_283),
.B(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_283),
.B(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.C(n_0),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_300),
.B(n_4),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_4),
.B(n_8),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_305),
.A3(n_9),
.B1(n_11),
.B2(n_4),
.C1(n_8),
.C2(n_0),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_302),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_301),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_296),
.B1(n_9),
.B2(n_1),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_0),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_0),
.Y(n_311)
);


endmodule