module fake_netlist_5_1117_n_1906 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1906);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1906;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_97),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_98),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_102),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_45),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_7),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_47),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_21),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_131),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_113),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_95),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_71),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_30),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_68),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_5),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_153),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_138),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_25),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_89),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_91),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_62),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_6),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_86),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_106),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_54),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_85),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_137),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_44),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_54),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_11),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_79),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_47),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_57),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_55),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_126),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_60),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_165),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_112),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_67),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_80),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_62),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_16),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_78),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_51),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_0),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_68),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_10),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_83),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_21),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_100),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_26),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_3),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_139),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_108),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_175),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_111),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_20),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_63),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_128),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_135),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_94),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_120),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_101),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_152),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_74),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_155),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_84),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_121),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_26),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_124),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_149),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_34),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_35),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_40),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_61),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_50),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_30),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_77),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_69),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_48),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_20),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_23),
.Y(n_317)
);

BUFx2_ASAP7_75t_SL g318 ( 
.A(n_22),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_117),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_40),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_57),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_61),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_10),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_169),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_24),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_42),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_125),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_114),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_93),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_75),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_109),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_19),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_87),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_39),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_76),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_63),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_136),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_4),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_65),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_146),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_38),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_19),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_115),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_28),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_56),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_49),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_16),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_130),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_2),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_193),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_193),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_198),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_215),
.B(n_178),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_352),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_219),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_232),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_215),
.B(n_1),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_177),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_180),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_352),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_181),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_244),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_245),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_232),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_182),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_244),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_221),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_250),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_250),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

BUFx6f_ASAP7_75t_SL g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_183),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_178),
.B(n_1),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_184),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_188),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_184),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_280),
.B(n_179),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_286),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_280),
.B(n_2),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_184),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_256),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_289),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_325),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_338),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_268),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_185),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_191),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_202),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_256),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_185),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_268),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_196),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_241),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_196),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_211),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_238),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_190),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_241),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_229),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_312),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_204),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_312),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_229),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_241),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_205),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_233),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_233),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_199),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_209),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_179),
.B(n_4),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_245),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_213),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_260),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_260),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_265),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_241),
.B(n_9),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_214),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_186),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_265),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_195),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_216),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_218),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_186),
.B(n_247),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_266),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_227),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_230),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_186),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_355),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_368),
.B(n_247),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_356),
.B(n_361),
.C(n_438),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_247),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_231),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_255),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_426),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_377),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_354),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_357),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_236),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_387),
.B(n_239),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_384),
.B(n_248),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_359),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_359),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_380),
.B(n_197),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_384),
.B(n_255),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_362),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_362),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_388),
.B(n_252),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_367),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_371),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_371),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_373),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_374),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_374),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_375),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_425),
.B(n_261),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_400),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_410),
.B(n_208),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_360),
.B(n_255),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_271),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

OA21x2_ASAP7_75t_L g513 ( 
.A1(n_406),
.A2(n_267),
.B(n_266),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_505),
.B(n_415),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_453),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_443),
.B(n_435),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_512),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_446),
.B(n_245),
.Y(n_526)
);

AND3x2_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_408),
.C(n_306),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_475),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_363),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_457),
.A2(n_365),
.B1(n_210),
.B2(n_235),
.Y(n_533)
);

BUFx4f_ASAP7_75t_L g534 ( 
.A(n_513),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_457),
.B(n_411),
.C(n_397),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_446),
.A2(n_358),
.B1(n_310),
.B2(n_308),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_477),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_470),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_364),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_475),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_477),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_189),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_505),
.B(n_415),
.C(n_309),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_502),
.A2(n_369),
.B1(n_376),
.B2(n_360),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_446),
.A2(n_310),
.B1(n_308),
.B2(n_378),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_492),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_492),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_459),
.B(n_360),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_443),
.B(n_366),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_491),
.B(n_369),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_508),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_370),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_446),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_444),
.B(n_379),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_513),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_456),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_459),
.B(n_369),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_441),
.B(n_417),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_446),
.B(n_245),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_491),
.B(n_376),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_456),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_453),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_476),
.B(n_382),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_441),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_463),
.A2(n_378),
.B1(n_311),
.B2(n_307),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_462),
.B(n_395),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_463),
.A2(n_267),
.B1(n_269),
.B2(n_272),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_462),
.B(n_396),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_508),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_476),
.B(n_398),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_510),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_463),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_508),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_517),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_510),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_473),
.B(n_399),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_473),
.B(n_416),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_459),
.B(n_376),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_479),
.B(n_407),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_445),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_479),
.B(n_420),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_488),
.B(n_407),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_445),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_424),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_517),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_245),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_501),
.B(n_427),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_507),
.B(n_437),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_445),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_501),
.B(n_407),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_507),
.B(n_463),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_503),
.B(n_432),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_517),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_441),
.B(n_423),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_448),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_441),
.B(n_436),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_463),
.B(n_228),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_517),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_517),
.Y(n_628)
);

BUFx8_ASAP7_75t_SL g629 ( 
.A(n_448),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_483),
.B(n_414),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_453),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_454),
.B(n_439),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_503),
.B(n_467),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_467),
.B(n_206),
.C(n_418),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_506),
.B(n_509),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_517),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_509),
.B(n_511),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_483),
.B(n_189),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_445),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_511),
.Y(n_643)
);

BUFx4f_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_453),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_483),
.B(n_421),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_506),
.B(n_245),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_480),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_483),
.B(n_200),
.C(n_194),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_483),
.A2(n_311),
.B1(n_281),
.B2(n_285),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_445),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_483),
.B(n_421),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_441),
.B(n_238),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_511),
.B(n_372),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_497),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g658 ( 
.A(n_454),
.B(n_203),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_441),
.B(n_238),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_511),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_486),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_478),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_442),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_458),
.B(n_238),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_486),
.B(n_383),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_489),
.B(n_386),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_458),
.B(n_328),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_506),
.B(n_274),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_489),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_578),
.B(n_458),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_531),
.B(n_520),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_661),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_561),
.B(n_506),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_578),
.B(n_458),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_521),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_661),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_526),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_556),
.A2(n_391),
.B1(n_392),
.B2(n_390),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_535),
.B(n_582),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_670),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_535),
.B(n_584),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_578),
.B(n_458),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_521),
.B(n_478),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_557),
.A2(n_269),
.B1(n_272),
.B2(n_349),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_614),
.B(n_207),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_600),
.B(n_506),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_609),
.B(n_212),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_618),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_561),
.A2(n_328),
.B1(n_331),
.B2(n_334),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_600),
.B(n_485),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_667),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_572),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_578),
.B(n_458),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_555),
.B(n_478),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_593),
.B(n_331),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_607),
.B(n_485),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_523),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_607),
.B(n_485),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_593),
.B(n_334),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_606),
.B(n_485),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_593),
.B(n_277),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_525),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_591),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_551),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_617),
.B(n_485),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_572),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_560),
.B(n_217),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_562),
.B(n_616),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_616),
.B(n_518),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_555),
.B(n_490),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_223),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_567),
.B(n_490),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_567),
.B(n_490),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_523),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_593),
.B(n_288),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_599),
.B(n_490),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_599),
.B(n_626),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_529),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_558),
.B(n_499),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_592),
.B(n_490),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_596),
.B(n_514),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_SL g726 ( 
.A1(n_533),
.A2(n_622),
.B1(n_662),
.B2(n_603),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_571),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_596),
.B(n_514),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_665),
.B(n_666),
.C(n_658),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_529),
.B(n_530),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_530),
.B(n_514),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_541),
.B(n_514),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_541),
.B(n_452),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_534),
.A2(n_447),
.B(n_442),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_613),
.B(n_226),
.C(n_225),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_655),
.B(n_240),
.C(n_237),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_545),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_545),
.B(n_452),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_525),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_540),
.A2(n_292),
.B1(n_350),
.B2(n_345),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_538),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_552),
.B(n_452),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_538),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_571),
.B(n_243),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_534),
.B(n_290),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_630),
.B(n_499),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_552),
.B(n_455),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_542),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_554),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_597),
.A2(n_296),
.B1(n_342),
.B2(n_336),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_554),
.B(n_455),
.Y(n_751)
);

INVx3_ASAP7_75t_R g752 ( 
.A(n_634),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_630),
.B(n_646),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_598),
.A2(n_319),
.B1(n_314),
.B2(n_329),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_557),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_634),
.B(n_515),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_563),
.A2(n_281),
.B1(n_349),
.B2(n_347),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_533),
.B(n_515),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_667),
.B(n_300),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_563),
.B(n_565),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_542),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_565),
.B(n_566),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_566),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_526),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_543),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_543),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_653),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_602),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_649),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_534),
.B(n_305),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_586),
.B(n_330),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_635),
.B(n_516),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_568),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_591),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_577),
.B(n_246),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_589),
.A2(n_546),
.B1(n_547),
.B2(n_654),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_568),
.B(n_455),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_639),
.B(n_469),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_612),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_615),
.B(n_469),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_527),
.B(n_249),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_633),
.B(n_253),
.C(n_251),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_586),
.B(n_332),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_632),
.B(n_258),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_649),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_586),
.B(n_497),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_537),
.B(n_516),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_583),
.A2(n_347),
.B(n_285),
.C(n_307),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_659),
.A2(n_279),
.B1(n_194),
.B2(n_304),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_544),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_652),
.B(n_469),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_667),
.B(n_526),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_636),
.B(n_471),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_624),
.B(n_497),
.Y(n_797)
);

AO221x1_ASAP7_75t_L g798 ( 
.A1(n_564),
.A2(n_320),
.B1(n_321),
.B2(n_335),
.C(n_294),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_636),
.B(n_471),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_544),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_641),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_641),
.B(n_471),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_612),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_643),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_643),
.B(n_472),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_647),
.B(n_472),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_591),
.Y(n_807)
);

NOR3xp33_ASAP7_75t_L g808 ( 
.A(n_625),
.B(n_262),
.C(n_259),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_669),
.A2(n_335),
.B(n_321),
.C(n_320),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_647),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_660),
.B(n_472),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_660),
.B(n_474),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_544),
.B(n_474),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_544),
.B(n_564),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_664),
.B(n_548),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_612),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_453),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_580),
.B(n_200),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_602),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_624),
.B(n_497),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_621),
.B(n_224),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_605),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_640),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_569),
.A2(n_278),
.B1(n_224),
.B2(n_304),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_481),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_640),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_605),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_605),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_564),
.B(n_474),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_573),
.B(n_497),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_605),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_650),
.B(n_481),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_573),
.B(n_497),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_624),
.B(n_497),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_629),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_602),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_644),
.B(n_528),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_573),
.B(n_242),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_640),
.A2(n_242),
.B1(n_254),
.B2(n_257),
.Y(n_839)
);

AND2x2_ASAP7_75t_SL g840 ( 
.A(n_644),
.B(n_254),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_644),
.B(n_257),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_672),
.B(n_620),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_723),
.B(n_651),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_672),
.A2(n_579),
.B1(n_573),
.B2(n_637),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_681),
.B(n_608),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_696),
.B(n_187),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_694),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_694),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_608),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_837),
.A2(n_576),
.B(n_528),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_781),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_683),
.B(n_278),
.C(n_275),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_690),
.B(n_187),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_708),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_711),
.B(n_187),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_709),
.Y(n_856)
);

NOR2x2_ASAP7_75t_L g857 ( 
.A(n_685),
.B(n_187),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_837),
.A2(n_576),
.B(n_528),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_707),
.A2(n_576),
.B(n_528),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_753),
.B(n_621),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_814),
.A2(n_764),
.B(n_762),
.Y(n_861)
);

AOI21xp33_ASAP7_75t_L g862 ( 
.A1(n_683),
.A2(n_279),
.B(n_275),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_721),
.A2(n_648),
.B(n_302),
.C(n_294),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_688),
.A2(n_585),
.B(n_581),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_692),
.A2(n_588),
.B(n_576),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_711),
.B(n_608),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_735),
.B(n_621),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_710),
.B(n_608),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_712),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_709),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_710),
.B(n_591),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_713),
.B(n_752),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_698),
.A2(n_604),
.B(n_588),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_781),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_687),
.B(n_591),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_687),
.B(n_642),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_234),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_700),
.A2(n_604),
.B(n_588),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_804),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_631),
.B(n_604),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_714),
.A2(n_645),
.B(n_631),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_716),
.A2(n_645),
.B(n_631),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_713),
.A2(n_689),
.B1(n_815),
.B2(n_753),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_745),
.A2(n_287),
.B(n_284),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_689),
.B(n_642),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_727),
.Y(n_888)
);

OAI321xp33_ASAP7_75t_L g889 ( 
.A1(n_778),
.A2(n_303),
.A3(n_302),
.B1(n_291),
.B2(n_287),
.C(n_284),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_645),
.B(n_631),
.Y(n_890)
);

NOR2x1p5_ASAP7_75t_SL g891 ( 
.A(n_755),
.B(n_559),
.Y(n_891)
);

NOR2x1_ASAP7_75t_R g892 ( 
.A(n_835),
.B(n_264),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_673),
.B(n_678),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_815),
.A2(n_758),
.B(n_686),
.C(n_777),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_686),
.A2(n_291),
.B(n_303),
.C(n_668),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_682),
.B(n_642),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_804),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_720),
.A2(n_645),
.B(n_519),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_781),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_677),
.B(n_579),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_803),
.B(n_668),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_810),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_746),
.B(n_755),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_765),
.B(n_642),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_697),
.A2(n_519),
.B(n_549),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_697),
.A2(n_519),
.B(n_549),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_790),
.A2(n_668),
.B(n_559),
.C(n_574),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_810),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_787),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_734),
.A2(n_590),
.B(n_587),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_758),
.A2(n_422),
.B(n_428),
.C(n_429),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_701),
.A2(n_519),
.B(n_550),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_765),
.B(n_587),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_803),
.B(n_816),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_759),
.B(n_757),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_775),
.B(n_590),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_775),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_701),
.A2(n_519),
.B(n_550),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_779),
.A2(n_794),
.B(n_772),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_756),
.B(n_595),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_760),
.B(n_769),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_772),
.A2(n_519),
.B(n_522),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_761),
.A2(n_797),
.B(n_788),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_788),
.A2(n_524),
.B(n_522),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_797),
.A2(n_524),
.B(n_522),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_813),
.A2(n_623),
.B(n_595),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_786),
.B(n_623),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_790),
.A2(n_841),
.B(n_691),
.C(n_719),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_820),
.A2(n_532),
.B(n_524),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_715),
.B(n_270),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_744),
.B(n_273),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_841),
.A2(n_559),
.B(n_574),
.C(n_575),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_777),
.A2(n_422),
.B(n_428),
.C(n_429),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_786),
.B(n_627),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_820),
.A2(n_834),
.B(n_800),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_627),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_774),
.B(n_276),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_834),
.A2(n_532),
.B(n_539),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_792),
.A2(n_532),
.B(n_539),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_770),
.B(n_430),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_699),
.B(n_638),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_675),
.A2(n_536),
.B(n_553),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_685),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_685),
.B(n_234),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_718),
.B(n_638),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_675),
.A2(n_539),
.B(n_553),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_703),
.A2(n_601),
.B(n_574),
.C(n_575),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_840),
.A2(n_579),
.B1(n_575),
.B2(n_610),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_722),
.B(n_663),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_680),
.B(n_430),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_737),
.B(n_663),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_770),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_749),
.B(n_663),
.Y(n_955)
);

O2A1O1Ixp5_ASAP7_75t_SL g956 ( 
.A1(n_839),
.A2(n_440),
.B(n_434),
.C(n_504),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_724),
.A2(n_619),
.B(n_594),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_675),
.A2(n_536),
.B(n_553),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_693),
.A2(n_536),
.B(n_628),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_795),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_818),
.A2(n_611),
.B1(n_570),
.B2(n_526),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_789),
.B(n_663),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_818),
.A2(n_434),
.B(n_440),
.C(n_481),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_801),
.Y(n_964)
);

NOR2x1_ASAP7_75t_L g965 ( 
.A(n_819),
.B(n_836),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_703),
.A2(n_601),
.B(n_594),
.C(n_610),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_840),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_782),
.B(n_594),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_803),
.B(n_601),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_822),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_693),
.A2(n_610),
.B(n_628),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_830),
.A2(n_619),
.B(n_628),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_793),
.B(n_619),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_780),
.A2(n_657),
.B(n_656),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_823),
.B(n_667),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_667),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_726),
.B(n_282),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_677),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_693),
.A2(n_657),
.B(n_656),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_674),
.A2(n_657),
.B(n_656),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_729),
.B(n_824),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_773),
.A2(n_442),
.B(n_447),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_730),
.A2(n_611),
.B(n_526),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_773),
.A2(n_442),
.B(n_447),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_829),
.A2(n_611),
.B(n_526),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_526),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_736),
.B(n_234),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_827),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_570),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_816),
.B(n_480),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_784),
.B(n_783),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_785),
.A2(n_447),
.B(n_460),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_833),
.A2(n_611),
.B(n_570),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_785),
.A2(n_468),
.B(n_466),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_816),
.A2(n_466),
.B(n_468),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_783),
.B(n_283),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_816),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_828),
.B(n_831),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_821),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_808),
.B(n_484),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_821),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_825),
.B(n_570),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_719),
.A2(n_611),
.B1(n_570),
.B2(n_579),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_791),
.B(n_293),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_705),
.A2(n_451),
.B(n_460),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_838),
.A2(n_484),
.B(n_494),
.C(n_504),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_705),
.A2(n_451),
.B(n_460),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_832),
.B(n_570),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_733),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_796),
.B(n_570),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_679),
.B(n_480),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_776),
.A2(n_461),
.B(n_466),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_731),
.A2(n_611),
.B(n_451),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_732),
.A2(n_611),
.B(n_451),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_738),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_704),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_SL g1017 ( 
.A1(n_809),
.A2(n_504),
.B(n_484),
.C(n_498),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_799),
.B(n_500),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_802),
.B(n_500),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_776),
.A2(n_468),
.B(n_460),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_671),
.A2(n_346),
.B1(n_297),
.B2(n_298),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_R g1022 ( 
.A(n_671),
.B(n_295),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_807),
.A2(n_468),
.B(n_461),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_805),
.B(n_500),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_807),
.A2(n_461),
.B(n_464),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_679),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_806),
.B(n_299),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_742),
.A2(n_461),
.B(n_464),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_747),
.Y(n_1029)
);

AND2x4_ASAP7_75t_SL g1030 ( 
.A(n_771),
.B(n_234),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1009),
.B(n_811),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_873),
.A2(n_817),
.B(n_679),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_842),
.B(n_679),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_894),
.A2(n_684),
.B1(n_676),
.B2(n_695),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1009),
.B(n_812),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_885),
.B(n_766),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_862),
.A2(n_798),
.B1(n_751),
.B2(n_263),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_916),
.B(n_725),
.Y(n_1038)
);

BUFx4_ASAP7_75t_SL g1039 ( 
.A(n_978),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_900),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_916),
.B(n_728),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_886),
.A2(n_695),
.B(n_684),
.C(n_676),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_877),
.A2(n_768),
.B(n_767),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_861),
.A2(n_887),
.B(n_878),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_R g1045 ( 
.A(n_842),
.B(n_766),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_860),
.B(n_766),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_894),
.A2(n_740),
.B(n_750),
.C(n_754),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_931),
.B(n_739),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_967),
.A2(n_766),
.B1(n_763),
.B2(n_748),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_896),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_866),
.B(n_741),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_931),
.A2(n_743),
.B(n_494),
.C(n_498),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_920),
.A2(n_858),
.B(n_850),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_888),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_932),
.B(n_494),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_932),
.B(n_496),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_848),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_967),
.A2(n_344),
.B1(n_315),
.B2(n_316),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1015),
.B(n_496),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_888),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1029),
.B(n_496),
.Y(n_1061)
);

CKINVDCx11_ASAP7_75t_R g1062 ( 
.A(n_892),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_874),
.B(n_313),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_981),
.A2(n_938),
.B(n_929),
.C(n_996),
.Y(n_1064)
);

BUFx8_ASAP7_75t_L g1065 ( 
.A(n_991),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_860),
.B(n_941),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_874),
.B(n_317),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_843),
.B(n_498),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_854),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_909),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_855),
.B(n_480),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_981),
.B(n_322),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_854),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1027),
.B(n_487),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_918),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_901),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_918),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_904),
.A2(n_351),
.B1(n_327),
.B2(n_333),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_847),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_852),
.A2(n_938),
.B(n_977),
.C(n_996),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_944),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_870),
.B(n_263),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1027),
.B(n_487),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_954),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_SL g1085 ( 
.A1(n_893),
.A2(n_960),
.B(n_867),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_977),
.A2(n_495),
.B(n_493),
.C(n_487),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1004),
.A2(n_348),
.B(n_324),
.C(n_337),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_L g1088 ( 
.A(n_1004),
.B(n_339),
.C(n_341),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_879),
.A2(n_849),
.B1(n_845),
.B2(n_964),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_922),
.B(n_487),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_882),
.A2(n_465),
.B(n_464),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_846),
.B(n_263),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_900),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_941),
.B(n_493),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_924),
.A2(n_465),
.B(n_464),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_859),
.A2(n_465),
.B(n_466),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_987),
.B(n_340),
.C(n_343),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_856),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_869),
.A2(n_500),
.B1(n_495),
.B2(n_493),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_962),
.B(n_495),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_944),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_945),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_883),
.A2(n_450),
.B(n_449),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_903),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_936),
.A2(n_495),
.B(n_493),
.C(n_450),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_902),
.A2(n_449),
.B1(n_134),
.B2(n_132),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_910),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_965),
.B(n_123),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_972),
.A2(n_449),
.B(n_453),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_954),
.B(n_453),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_872),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_952),
.B(n_174),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_900),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_896),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_900),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_902),
.A2(n_119),
.B1(n_81),
.B2(n_172),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_876),
.B(n_166),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_881),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_853),
.B(n_301),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_884),
.A2(n_453),
.B(n_162),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_898),
.Y(n_1121)
);

OAI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_1030),
.A2(n_301),
.B(n_263),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_876),
.B(n_301),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_964),
.B(n_301),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_937),
.B(n_9),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_896),
.B(n_11),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_921),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_901),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_963),
.B(n_12),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_963),
.B(n_12),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1030),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1000),
.B(n_968),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1000),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1001),
.B(n_970),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_988),
.B(n_13),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_890),
.A2(n_161),
.B(n_150),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_L g1137 ( 
.A(n_1021),
.B(n_14),
.C(n_15),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_999),
.A2(n_143),
.B1(n_141),
.B2(n_118),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_951),
.B(n_116),
.Y(n_1139)
);

AO32x2_ASAP7_75t_L g1140 ( 
.A1(n_949),
.A2(n_14),
.A3(n_15),
.B1(n_18),
.B2(n_22),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_857),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_868),
.A2(n_999),
.B1(n_915),
.B2(n_986),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_1022),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_908),
.A2(n_18),
.B(n_25),
.C(n_27),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_915),
.A2(n_99),
.B1(n_92),
.B2(n_90),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_989),
.A2(n_88),
.B1(n_73),
.B2(n_33),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_997),
.B(n_31),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_889),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_865),
.A2(n_37),
.B(n_41),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_875),
.A2(n_42),
.B(n_43),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_880),
.A2(n_67),
.B(n_46),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_934),
.A2(n_43),
.B(n_48),
.C(n_49),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1016),
.B(n_50),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_851),
.A2(n_66),
.B1(n_53),
.B2(n_55),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_905),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1026),
.A2(n_66),
.B(n_58),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_997),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_851),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_871),
.B(n_52),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_871),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_897),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_928),
.B(n_52),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_935),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_R g1165 ( 
.A(n_975),
.B(n_59),
.Y(n_1165)
);

CKINVDCx8_ASAP7_75t_R g1166 ( 
.A(n_934),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_998),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_895),
.A2(n_64),
.B(n_65),
.C(n_912),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1026),
.A2(n_64),
.B(n_844),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_973),
.B(n_895),
.Y(n_1170)
);

CKINVDCx16_ASAP7_75t_R g1171 ( 
.A(n_1003),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_899),
.A2(n_911),
.B(n_947),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_943),
.A2(n_958),
.B(n_959),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_969),
.A2(n_971),
.B(n_979),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1010),
.A2(n_983),
.B(n_939),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_942),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_969),
.A2(n_976),
.B(n_974),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_946),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_914),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_917),
.A2(n_864),
.B(n_1018),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_SL g1181 ( 
.A1(n_990),
.A2(n_957),
.B(n_927),
.C(n_1024),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_961),
.B(n_1002),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1019),
.B(n_912),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_994),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_990),
.B(n_1011),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_1008),
.B(n_961),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1173),
.A2(n_1174),
.B(n_1053),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_1115),
.B(n_1011),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1101),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1064),
.A2(n_950),
.B1(n_953),
.B2(n_955),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1038),
.B(n_891),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1041),
.B(n_1006),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_1172),
.B(n_1180),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1080),
.A2(n_863),
.B(n_948),
.C(n_966),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_1169),
.A3(n_1177),
.B(n_1144),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1166),
.A2(n_985),
.B1(n_993),
.B2(n_1013),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1085),
.A2(n_923),
.B(n_980),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_1043),
.A2(n_984),
.B(n_982),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1088),
.A2(n_940),
.B(n_933),
.C(n_992),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1175),
.A2(n_1017),
.B(n_930),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1109),
.A2(n_1095),
.B(n_1091),
.Y(n_1201)
);

AOI221x1_ASAP7_75t_L g1202 ( 
.A1(n_1137),
.A2(n_926),
.B1(n_925),
.B2(n_1028),
.C(n_1014),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1092),
.B(n_956),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1184),
.A2(n_1007),
.B(n_1023),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1033),
.A2(n_906),
.B(n_907),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1050),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1137),
.A2(n_1012),
.B1(n_1020),
.B2(n_1025),
.C(n_1005),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1046),
.Y(n_1208)
);

AO22x2_ASAP7_75t_L g1209 ( 
.A1(n_1088),
.A2(n_1163),
.B1(n_1164),
.B2(n_1072),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1047),
.A2(n_1067),
.B(n_1063),
.C(n_1112),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1052),
.A2(n_1042),
.B(n_1089),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1048),
.A2(n_913),
.B(n_919),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1046),
.Y(n_1213)
);

NAND2x1_ASAP7_75t_L g1214 ( 
.A(n_1158),
.B(n_995),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1074),
.A2(n_1017),
.B(n_1083),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1119),
.B(n_1063),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1115),
.B(n_1158),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1040),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_1032),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1081),
.B(n_1054),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1105),
.A2(n_1099),
.A3(n_1152),
.B(n_1150),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1170),
.A2(n_1071),
.B(n_1132),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1181),
.A2(n_1089),
.B(n_1052),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1151),
.A2(n_1183),
.A3(n_1125),
.B(n_1103),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1031),
.B(n_1035),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_SL g1227 ( 
.A1(n_1163),
.A2(n_1130),
.B(n_1129),
.C(n_1182),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1067),
.A2(n_1097),
.B1(n_1171),
.B2(n_1133),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1082),
.A2(n_1076),
.B1(n_1143),
.B2(n_1131),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1036),
.A2(n_1042),
.B(n_1100),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1054),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1066),
.B(n_1060),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1108),
.B(n_1117),
.Y(n_1234)
);

AO32x1_ASAP7_75t_L g1235 ( 
.A1(n_1140),
.A2(n_1106),
.A3(n_1116),
.B1(n_1058),
.B2(n_1138),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1097),
.A2(n_1149),
.B(n_1122),
.C(n_1176),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1049),
.A2(n_1120),
.A3(n_1096),
.B(n_1136),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1068),
.A2(n_1090),
.B(n_1179),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1059),
.A2(n_1061),
.B1(n_1178),
.B2(n_1111),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_1128),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1066),
.A2(n_1148),
.B1(n_1126),
.B2(n_1160),
.Y(n_1241)
);

OAI22x1_ASAP7_75t_L g1242 ( 
.A1(n_1148),
.A2(n_1134),
.B1(n_1143),
.B2(n_1155),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1134),
.B(n_1060),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1178),
.A2(n_1098),
.B1(n_1121),
.B2(n_1162),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1117),
.A2(n_1142),
.B(n_1139),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1115),
.A2(n_1156),
.B(n_1162),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1050),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1115),
.A2(n_1094),
.B(n_1086),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1185),
.A2(n_1045),
.B(n_1110),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1057),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1040),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1087),
.A2(n_1153),
.B(n_1135),
.C(n_1126),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1084),
.B(n_1123),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1084),
.B(n_1124),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1045),
.A2(n_1123),
.B(n_1069),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1062),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1147),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1051),
.B(n_1118),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1070),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_1165),
.B1(n_1154),
.B2(n_1104),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1078),
.B(n_1114),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1186),
.A2(n_1165),
.B(n_1145),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_SL g1263 ( 
.A1(n_1157),
.A2(n_1146),
.B(n_1077),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1073),
.A2(n_1075),
.B(n_1168),
.Y(n_1264)
);

AOI221x1_ASAP7_75t_L g1265 ( 
.A1(n_1140),
.A2(n_1113),
.B1(n_1093),
.B2(n_1107),
.C(n_1040),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1159),
.A2(n_1140),
.A3(n_1037),
.B(n_1186),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1140),
.A2(n_1037),
.B(n_1040),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1161),
.B(n_1093),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1113),
.B(n_1102),
.Y(n_1269)
);

BUFx4f_ASAP7_75t_SL g1270 ( 
.A(n_1065),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1065),
.A2(n_1039),
.B(n_1141),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1039),
.B(n_672),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1034),
.A2(n_1064),
.A3(n_886),
.B(n_1044),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1064),
.A2(n_672),
.B1(n_683),
.B2(n_681),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1080),
.B(n_672),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1070),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1064),
.B(n_672),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1101),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1062),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1046),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1054),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1101),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1066),
.B(n_1114),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1290)
);

INVx3_ASAP7_75t_SL g1291 ( 
.A(n_1128),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1292)
);

AO22x1_ASAP7_75t_L g1293 ( 
.A1(n_1088),
.A2(n_672),
.B1(n_842),
.B2(n_683),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1101),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1064),
.A2(n_894),
.B(n_1080),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1080),
.B(n_672),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1064),
.B(n_672),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1080),
.B(n_672),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1080),
.A2(n_842),
.B(n_672),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1080),
.B(n_672),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_L g1302 ( 
.A1(n_1064),
.A2(n_1137),
.B1(n_862),
.B2(n_1034),
.C(n_1088),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1064),
.A2(n_894),
.B(n_1034),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1080),
.A2(n_672),
.B(n_683),
.C(n_681),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1054),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1080),
.A2(n_672),
.B(n_1064),
.C(n_842),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1064),
.A2(n_672),
.B1(n_683),
.B2(n_681),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1063),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1034),
.A2(n_1064),
.A3(n_886),
.B(n_1044),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_L g1311 ( 
.A(n_1115),
.B(n_885),
.Y(n_1311)
);

AOI221x1_ASAP7_75t_L g1312 ( 
.A1(n_1064),
.A2(n_1137),
.B1(n_862),
.B2(n_1034),
.C(n_1088),
.Y(n_1312)
);

OAI22x1_ASAP7_75t_L g1313 ( 
.A1(n_1072),
.A2(n_842),
.B1(n_672),
.B2(n_778),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1034),
.A2(n_1064),
.A3(n_886),
.B(n_1044),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1066),
.B(n_1114),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1054),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1034),
.A2(n_1064),
.A3(n_886),
.B(n_1044),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1063),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1054),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1092),
.B(n_696),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1322)
);

AO32x2_ASAP7_75t_L g1323 ( 
.A1(n_1034),
.A2(n_1164),
.A3(n_691),
.B1(n_1099),
.B2(n_1140),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1064),
.B(n_672),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1070),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1133),
.B(n_1147),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1044),
.A2(n_693),
.B(n_675),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1173),
.A2(n_972),
.B(n_1174),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1080),
.B(n_672),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1080),
.A2(n_672),
.B(n_683),
.C(n_681),
.Y(n_1334)
);

INVx3_ASAP7_75t_SL g1335 ( 
.A(n_1128),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1031),
.B(n_672),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1064),
.A2(n_894),
.B(n_1080),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1101),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1080),
.A2(n_672),
.B(n_683),
.C(n_681),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1039),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1034),
.A2(n_1064),
.A3(n_886),
.B(n_1044),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1092),
.B(n_696),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1064),
.B(n_672),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1064),
.A2(n_672),
.B1(n_894),
.B2(n_842),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1080),
.B(n_672),
.C(n_1064),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1070),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1044),
.A2(n_1052),
.B(n_1175),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_1345),
.B2(n_1299),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1283),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1220),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1233),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1256),
.Y(n_1352)
);

CKINVDCx11_ASAP7_75t_R g1353 ( 
.A(n_1240),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1345),
.A2(n_1301),
.B1(n_1333),
.B2(n_1296),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1206),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1296),
.A2(n_1337),
.B1(n_1276),
.B2(n_1308),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1340),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1309),
.A2(n_1319),
.B1(n_1216),
.B2(n_1209),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1280),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1206),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1309),
.A2(n_1319),
.B1(n_1209),
.B2(n_1344),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1228),
.A2(n_1308),
.B(n_1276),
.Y(n_1362)
);

INVx6_ASAP7_75t_L g1363 ( 
.A(n_1247),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1337),
.A2(n_1344),
.B1(n_1300),
.B2(n_1313),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1247),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1291),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1281),
.A2(n_1324),
.B1(n_1298),
.B2(n_1343),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1250),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1328),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1240),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1336),
.A2(n_1334),
.B1(n_1339),
.B2(n_1305),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1281),
.A2(n_1298),
.B1(n_1343),
.B2(n_1324),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1189),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1346),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1229),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1242),
.A2(n_1262),
.B1(n_1228),
.B2(n_1260),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1335),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1293),
.A2(n_1321),
.B1(n_1342),
.B2(n_1272),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1286),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1257),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1247),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1254),
.B(n_1288),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1251),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1210),
.A2(n_1241),
.B1(n_1226),
.B2(n_1307),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1267),
.A2(n_1262),
.B1(n_1234),
.B2(n_1239),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1244),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1234),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1234),
.A2(n_1239),
.B1(n_1196),
.B2(n_1192),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_SL g1389 ( 
.A(n_1282),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1243),
.B(n_1234),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1270),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1295),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1253),
.A2(n_1252),
.B1(n_1261),
.B2(n_1236),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1306),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1203),
.A2(n_1230),
.B1(n_1196),
.B2(n_1338),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1288),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1244),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1258),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1263),
.A2(n_1311),
.B1(n_1192),
.B2(n_1329),
.Y(n_1399)
);

BUFx2_ASAP7_75t_SL g1400 ( 
.A(n_1257),
.Y(n_1400)
);

BUFx2_ASAP7_75t_SL g1401 ( 
.A(n_1315),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1269),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1271),
.A2(n_1302),
.B1(n_1312),
.B2(n_1303),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1311),
.A2(n_1315),
.B1(n_1329),
.B2(n_1213),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1329),
.A2(n_1284),
.B1(n_1208),
.B2(n_1213),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1221),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1320),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1223),
.A2(n_1238),
.B1(n_1316),
.B2(n_1232),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1316),
.A2(n_1224),
.B1(n_1285),
.B2(n_1190),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1190),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1245),
.A2(n_1191),
.B1(n_1255),
.B2(n_1246),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1265),
.A2(n_1194),
.B(n_1224),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1211),
.A2(n_1284),
.B1(n_1208),
.B2(n_1191),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1268),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1218),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1249),
.A2(n_1248),
.B1(n_1219),
.B2(n_1217),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1218),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1266),
.Y(n_1418)
);

OAI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1264),
.A2(n_1202),
.B1(n_1231),
.B2(n_1235),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1188),
.A2(n_1199),
.B1(n_1197),
.B2(n_1347),
.Y(n_1420)
);

CKINVDCx11_ASAP7_75t_R g1421 ( 
.A(n_1227),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1214),
.B2(n_1193),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1274),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1200),
.A2(n_1215),
.B1(n_1235),
.B2(n_1212),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1275),
.A2(n_1290),
.B1(n_1277),
.B2(n_1331),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1200),
.A2(n_1215),
.B1(n_1323),
.B2(n_1198),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1225),
.B(n_1341),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1323),
.A2(n_1198),
.B1(n_1187),
.B2(n_1332),
.Y(n_1428)
);

AOI21xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1273),
.A2(n_1325),
.B(n_1322),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1323),
.A2(n_1195),
.B1(n_1292),
.B2(n_1294),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1304),
.A2(n_1330),
.B1(n_1204),
.B2(n_1327),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1279),
.A2(n_1287),
.B1(n_1326),
.B2(n_1317),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1195),
.A2(n_1289),
.B1(n_1341),
.B2(n_1274),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1207),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1225),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1201),
.A2(n_1310),
.B1(n_1314),
.B2(n_1318),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1310),
.A2(n_1314),
.B1(n_1318),
.B2(n_1341),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1225),
.Y(n_1438)
);

INVx8_ASAP7_75t_L g1439 ( 
.A(n_1318),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1222),
.B(n_1237),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1222),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1222),
.A2(n_672),
.B1(n_1308),
.B2(n_1276),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1237),
.A2(n_672),
.B1(n_1308),
.B2(n_1276),
.Y(n_1443)
);

BUFx4f_ASAP7_75t_L g1444 ( 
.A(n_1206),
.Y(n_1444)
);

BUFx4_ASAP7_75t_SL g1445 ( 
.A(n_1340),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_681),
.B2(n_683),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1278),
.A2(n_672),
.B1(n_1297),
.B2(n_683),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1206),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_681),
.B2(n_683),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1336),
.B2(n_1297),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1276),
.A2(n_672),
.B1(n_1308),
.B2(n_842),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1336),
.B2(n_1297),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_681),
.B2(n_683),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1278),
.A2(n_672),
.B1(n_1297),
.B2(n_842),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1233),
.Y(n_1455)
);

CKINVDCx6p67_ASAP7_75t_R g1456 ( 
.A(n_1256),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1283),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1206),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1336),
.B(n_672),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1321),
.B(n_1342),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1276),
.A2(n_672),
.B1(n_1308),
.B2(n_842),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1220),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1336),
.B2(n_1297),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_681),
.B2(n_683),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1220),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1278),
.A2(n_672),
.B1(n_1297),
.B2(n_683),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1189),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1220),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_681),
.B2(n_683),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1311),
.B(n_1115),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1259),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1233),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1321),
.B(n_1342),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1256),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1220),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1220),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1336),
.B(n_672),
.Y(n_1477)
);

BUFx4_ASAP7_75t_SL g1478 ( 
.A(n_1340),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_672),
.B2(n_1088),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1283),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1425),
.A2(n_1431),
.B(n_1432),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1427),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1387),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1387),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1443),
.A2(n_1442),
.A3(n_1420),
.B(n_1438),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1418),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1447),
.B(n_1466),
.Y(n_1488)
);

AO21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1385),
.A2(n_1376),
.B(n_1356),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1364),
.B(n_1356),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1410),
.A2(n_1479),
.B1(n_1454),
.B2(n_1469),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1460),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1386),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1387),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1364),
.B(n_1440),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1362),
.A2(n_1453),
.B(n_1446),
.C(n_1469),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1446),
.A2(n_1464),
.B1(n_1453),
.B2(n_1449),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1449),
.A2(n_1464),
.B1(n_1393),
.B2(n_1451),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1438),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1348),
.B(n_1354),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1435),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1439),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1397),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1439),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1439),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1375),
.B(n_1459),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1429),
.A2(n_1419),
.B(n_1416),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1368),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1407),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1473),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1350),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1406),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1411),
.A2(n_1422),
.B(n_1371),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1387),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1348),
.B(n_1437),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1354),
.B(n_1395),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1434),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1394),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1462),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1434),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1465),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1468),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1419),
.A2(n_1412),
.B(n_1463),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1404),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1431),
.A2(n_1432),
.B(n_1436),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1476),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1423),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1436),
.A2(n_1428),
.B(n_1424),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1396),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1421),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1428),
.A2(n_1424),
.B(n_1437),
.Y(n_1532)
);

NOR3xp33_ASAP7_75t_L g1533 ( 
.A(n_1461),
.B(n_1384),
.C(n_1403),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1426),
.A2(n_1385),
.B(n_1409),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1349),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1433),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1351),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1405),
.B(n_1399),
.Y(n_1538)
);

BUFx2_ASAP7_75t_SL g1539 ( 
.A(n_1398),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1470),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1409),
.B(n_1450),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1430),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1450),
.A2(n_1452),
.B(n_1463),
.Y(n_1543)
);

CKINVDCx6p67_ASAP7_75t_R g1544 ( 
.A(n_1457),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1396),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1361),
.A2(n_1452),
.B1(n_1358),
.B2(n_1378),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1455),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1413),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1388),
.B(n_1367),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1359),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1401),
.B(n_1390),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1388),
.A2(n_1408),
.B(n_1372),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1367),
.B(n_1372),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1472),
.B(n_1414),
.Y(n_1554)
);

AOI21xp33_ASAP7_75t_L g1555 ( 
.A1(n_1477),
.A2(n_1408),
.B(n_1379),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1415),
.A2(n_1374),
.B(n_1471),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1369),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1382),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1417),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1444),
.A2(n_1402),
.B(n_1392),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1389),
.A2(n_1370),
.B1(n_1396),
.B2(n_1400),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_SL g1562 ( 
.A(n_1474),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1383),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1355),
.B(n_1467),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1373),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1360),
.B(n_1458),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1458),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1458),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1363),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1389),
.A2(n_1444),
.B(n_1448),
.Y(n_1570)
);

AOI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1363),
.A2(n_1381),
.B(n_1448),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1353),
.Y(n_1572)
);

AND2x6_ASAP7_75t_L g1573 ( 
.A(n_1484),
.B(n_1381),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1562),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1526),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1542),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1488),
.B(n_1366),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_R g1578 ( 
.A(n_1535),
.B(n_1480),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1543),
.A2(n_1391),
.B(n_1377),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1553),
.B(n_1365),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1533),
.A2(n_1365),
.B(n_1478),
.C(n_1445),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1495),
.B(n_1456),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1496),
.A2(n_1380),
.B(n_1445),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1509),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1526),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1494),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1552),
.A2(n_1478),
.B(n_1474),
.C(n_1352),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1491),
.A2(n_1357),
.B1(n_1498),
.B2(n_1546),
.C(n_1497),
.Y(n_1588)
);

BUFx2_ASAP7_75t_R g1589 ( 
.A(n_1523),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1498),
.A2(n_1552),
.B1(n_1555),
.B2(n_1541),
.C(n_1560),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_SL g1593 ( 
.A(n_1539),
.B(n_1551),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1565),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1483),
.B(n_1495),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1541),
.A2(n_1528),
.B1(n_1531),
.B2(n_1516),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1518),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1508),
.B(n_1511),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_L g1599 ( 
.A(n_1516),
.B(n_1513),
.C(n_1500),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1490),
.A2(n_1500),
.B(n_1549),
.C(n_1539),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1492),
.B(n_1510),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1513),
.B(n_1481),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1512),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1528),
.A2(n_1515),
.B(n_1506),
.C(n_1563),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1525),
.A2(n_1481),
.B(n_1529),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1531),
.A2(n_1561),
.B1(n_1524),
.B2(n_1490),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1525),
.A2(n_1529),
.B(n_1499),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_SL g1609 ( 
.A(n_1551),
.B(n_1489),
.Y(n_1609)
);

AO32x2_ASAP7_75t_L g1610 ( 
.A1(n_1519),
.A2(n_1522),
.A3(n_1494),
.B1(n_1568),
.B2(n_1530),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1548),
.B(n_1549),
.C(n_1524),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1548),
.A2(n_1515),
.B(n_1538),
.C(n_1532),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1518),
.A2(n_1547),
.B1(n_1537),
.B2(n_1554),
.C(n_1538),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1538),
.A2(n_1501),
.B(n_1569),
.C(n_1545),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1531),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1538),
.A2(n_1570),
.B(n_1556),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1531),
.A2(n_1551),
.B1(n_1564),
.B2(n_1572),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1532),
.A2(n_1520),
.B(n_1517),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1531),
.B(n_1544),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1570),
.A2(n_1556),
.B(n_1551),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1507),
.A2(n_1551),
.B(n_1494),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1521),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1507),
.A2(n_1534),
.B(n_1485),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1563),
.A2(n_1501),
.B(n_1571),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1527),
.B(n_1486),
.Y(n_1626)
);

INVx5_ASAP7_75t_SL g1627 ( 
.A(n_1572),
.Y(n_1627)
);

NAND4xp25_ASAP7_75t_L g1628 ( 
.A(n_1493),
.B(n_1503),
.C(n_1559),
.D(n_1550),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1575),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1502),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1486),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1623),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1487),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1610),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1588),
.A2(n_1589),
.B1(n_1591),
.B2(n_1600),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.B(n_1486),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1599),
.A2(n_1534),
.B1(n_1531),
.B2(n_1544),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1590),
.B(n_1486),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1623),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1592),
.B(n_1486),
.Y(n_1640)
);

AND2x2_ASAP7_75t_SL g1641 ( 
.A(n_1592),
.B(n_1534),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1595),
.B(n_1486),
.Y(n_1642)
);

INVx6_ASAP7_75t_L g1643 ( 
.A(n_1573),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1585),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1611),
.A2(n_1489),
.B1(n_1534),
.B2(n_1572),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1579),
.A2(n_1572),
.B1(n_1550),
.B2(n_1557),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1482),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1597),
.Y(n_1648)
);

OR2x6_ASAP7_75t_SL g1649 ( 
.A(n_1618),
.B(n_1505),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_1578),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1619),
.B(n_1482),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1598),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1609),
.A2(n_1572),
.B1(n_1484),
.B2(n_1485),
.Y(n_1653)
);

AND2x4_ASAP7_75t_SL g1654 ( 
.A(n_1586),
.B(n_1514),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1610),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1596),
.A2(n_1572),
.B1(n_1504),
.B2(n_1540),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1651),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1644),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1644),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1635),
.A2(n_1612),
.B1(n_1600),
.B2(n_1587),
.C(n_1613),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1651),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1651),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1624),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1607),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_SL g1667 ( 
.A(n_1650),
.B(n_1574),
.C(n_1581),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1633),
.B(n_1612),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1654),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1633),
.B(n_1576),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1655),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1576),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1656),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1602),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1638),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1645),
.A2(n_1581),
.B1(n_1606),
.B2(n_1582),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1636),
.B(n_1622),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1637),
.A2(n_1583),
.B(n_1604),
.C(n_1614),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1635),
.A2(n_1620),
.B1(n_1574),
.B2(n_1577),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1645),
.A2(n_1601),
.B1(n_1603),
.B2(n_1580),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1637),
.A2(n_1628),
.B1(n_1594),
.B2(n_1608),
.Y(n_1684)
);

INVx5_ASAP7_75t_SL g1685 ( 
.A(n_1630),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1648),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1638),
.A2(n_1604),
.B(n_1617),
.C(n_1584),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1643),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1593),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1639),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1629),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1640),
.B(n_1621),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1639),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1674),
.B(n_1631),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1665),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1658),
.B(n_1671),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1665),
.B(n_1631),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.B(n_1671),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1673),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1673),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1676),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1685),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1682),
.B(n_1650),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1668),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1686),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1658),
.B(n_1640),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1668),
.B(n_1652),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1690),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1659),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1690),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1665),
.B(n_1642),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1685),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1660),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1659),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1693),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1693),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1660),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1661),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1652),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1691),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1691),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1659),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1663),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1663),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1706),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1696),
.B(n_1677),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1696),
.B(n_1681),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1714),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1702),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1696),
.B(n_1681),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1714),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1718),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1706),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1703),
.A2(n_1662),
.B(n_1687),
.C(n_1680),
.Y(n_1741)
);

OAI31xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1698),
.A2(n_1680),
.A3(n_1684),
.B(n_1662),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1718),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1719),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1675),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1698),
.B(n_1692),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1707),
.B(n_1692),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1719),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_1692),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1708),
.B(n_1664),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1697),
.B(n_1675),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1699),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1699),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1700),
.B(n_1701),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1707),
.B(n_1666),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1700),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1695),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1695),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1723),
.Y(n_1762)
);

NAND2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1702),
.B(n_1669),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1715),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1702),
.B(n_1666),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1722),
.B(n_1666),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1701),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1705),
.B(n_1679),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1705),
.B(n_1679),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1695),
.B(n_1679),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1755),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1765),
.B(n_1685),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1755),
.Y(n_1773)
);

NAND2x1_ASAP7_75t_L g1774 ( 
.A(n_1734),
.B(n_1702),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1756),
.Y(n_1775)
);

XOR2xp5_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1682),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1741),
.B(n_1684),
.C(n_1678),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1729),
.B(n_1730),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1729),
.B(n_1713),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1756),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1728),
.B(n_1697),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1728),
.B(n_1713),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1742),
.A2(n_1683),
.B(n_1678),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1739),
.B(n_1697),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1765),
.B(n_1685),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1759),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1712),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1742),
.B(n_1720),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1759),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1729),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1767),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1731),
.B(n_1720),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1667),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1670),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1760),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1732),
.B(n_1747),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1732),
.B(n_1712),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1747),
.B(n_1712),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1763),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1736),
.B(n_1713),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1760),
.B(n_1672),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1767),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1761),
.B(n_1672),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1761),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1736),
.B(n_1722),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1776),
.B(n_1667),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1798),
.B(n_1770),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1783),
.A2(n_1762),
.B(n_1737),
.Y(n_1811)
);

OAI32xp33_ASAP7_75t_L g1812 ( 
.A1(n_1788),
.A2(n_1770),
.A3(n_1763),
.B1(n_1754),
.B2(n_1649),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1777),
.A2(n_1762),
.B(n_1683),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1777),
.A2(n_1687),
.B1(n_1646),
.B2(n_1657),
.C(n_1735),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1797),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1797),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1806),
.B(n_1733),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_SL g1818 ( 
.A(n_1801),
.B(n_1770),
.C(n_1737),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1771),
.B(n_1733),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1781),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1773),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1782),
.A2(n_1649),
.B1(n_1784),
.B2(n_1787),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1794),
.A2(n_1782),
.B1(n_1780),
.B2(n_1804),
.C(n_1791),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1775),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1736),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1790),
.A2(n_1649),
.B1(n_1688),
.B2(n_1753),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1786),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1790),
.A2(n_1653),
.B1(n_1749),
.B2(n_1752),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1789),
.Y(n_1829)
);

AOI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1794),
.A2(n_1765),
.B(n_1735),
.C(n_1734),
.Y(n_1830)
);

OR4x1_ASAP7_75t_L g1831 ( 
.A(n_1774),
.B(n_1746),
.C(n_1745),
.D(n_1738),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1779),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1792),
.B(n_1738),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1820),
.B(n_1793),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1815),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1811),
.B(n_1793),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1809),
.B(n_1779),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1823),
.A2(n_1807),
.B(n_1785),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1816),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_R g1840 ( 
.A(n_1808),
.B(n_1734),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1819),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1813),
.A2(n_1805),
.B(n_1803),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1811),
.A2(n_1823),
.B1(n_1814),
.B2(n_1818),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1832),
.B(n_1779),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1832),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1814),
.A2(n_1802),
.B1(n_1795),
.B2(n_1796),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1828),
.A2(n_1802),
.B1(n_1795),
.B2(n_1772),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1825),
.Y(n_1848)
);

AOI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1812),
.A2(n_1795),
.B1(n_1802),
.B2(n_1751),
.C1(n_1746),
.C2(n_1745),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1822),
.A2(n_1830),
.B(n_1833),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1817),
.A2(n_1734),
.B(n_1735),
.C(n_1751),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1807),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1819),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1843),
.A2(n_1826),
.B1(n_1810),
.B2(n_1831),
.C(n_1833),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1844),
.Y(n_1855)
);

AOI211xp5_ASAP7_75t_L g1856 ( 
.A1(n_1850),
.A2(n_1817),
.B(n_1827),
.C(n_1824),
.Y(n_1856)
);

AOI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1843),
.A2(n_1829),
.B(n_1821),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1848),
.B(n_1749),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1852),
.B(n_1848),
.Y(n_1859)
);

AO22x2_ASAP7_75t_L g1860 ( 
.A1(n_1845),
.A2(n_1735),
.B1(n_1740),
.B2(n_1744),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1845),
.B(n_1749),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1849),
.A2(n_1799),
.B(n_1800),
.C(n_1753),
.Y(n_1862)
);

OAI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1836),
.A2(n_1754),
.B1(n_1769),
.B2(n_1768),
.Y(n_1863)
);

CKINVDCx14_ASAP7_75t_R g1864 ( 
.A(n_1840),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1837),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1859),
.B(n_1835),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1854),
.A2(n_1864),
.B(n_1857),
.C(n_1856),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1855),
.B(n_1839),
.C(n_1838),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1858),
.A2(n_1840),
.B(n_1847),
.Y(n_1869)
);

NAND3x1_ASAP7_75t_L g1870 ( 
.A(n_1861),
.B(n_1834),
.C(n_1841),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1862),
.A2(n_1842),
.B1(n_1846),
.B2(n_1853),
.Y(n_1871)
);

NOR3xp33_ASAP7_75t_L g1872 ( 
.A(n_1865),
.B(n_1851),
.C(n_1765),
.Y(n_1872)
);

NAND4xp25_ASAP7_75t_L g1873 ( 
.A(n_1863),
.B(n_1765),
.C(n_1646),
.D(n_1653),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1860),
.B(n_1743),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1871),
.A2(n_1860),
.B1(n_1740),
.B2(n_1744),
.C(n_1764),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1867),
.A2(n_1769),
.B(n_1768),
.C(n_1764),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1869),
.B(n_1757),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1868),
.A2(n_1766),
.B(n_1758),
.C(n_1752),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1870),
.A2(n_1694),
.B1(n_1743),
.B2(n_1752),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1879),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1877),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1878),
.Y(n_1882)
);

AOI211x1_ASAP7_75t_L g1883 ( 
.A1(n_1876),
.A2(n_1874),
.B(n_1873),
.C(n_1866),
.Y(n_1883)
);

AOI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1875),
.A2(n_1872),
.B(n_1766),
.C(n_1764),
.Y(n_1884)
);

AOI222xp33_ASAP7_75t_L g1885 ( 
.A1(n_1879),
.A2(n_1750),
.B1(n_1758),
.B2(n_1740),
.C1(n_1748),
.C2(n_1744),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1882),
.A2(n_1766),
.B1(n_1750),
.B2(n_1758),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1880),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1881),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1883),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1884),
.Y(n_1890)
);

NAND4xp25_ASAP7_75t_L g1891 ( 
.A(n_1887),
.B(n_1885),
.C(n_1615),
.D(n_1750),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1888),
.Y(n_1892)
);

NOR3x1_ASAP7_75t_L g1893 ( 
.A(n_1889),
.B(n_1757),
.C(n_1723),
.Y(n_1893)
);

AOI211x1_ASAP7_75t_L g1894 ( 
.A1(n_1891),
.A2(n_1890),
.B(n_1886),
.C(n_1743),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1894),
.A2(n_1892),
.B1(n_1893),
.B2(n_1748),
.Y(n_1895)
);

AOI22x1_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1748),
.B1(n_1566),
.B2(n_1724),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1895),
.Y(n_1897)
);

AOI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1724),
.B(n_1715),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1896),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1898),
.A2(n_1724),
.B(n_1715),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1899),
.A2(n_1721),
.B1(n_1627),
.B2(n_1725),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1721),
.B(n_1725),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1900),
.B(n_1725),
.Y(n_1903)
);

OAI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1694),
.B1(n_1726),
.B2(n_1727),
.Y(n_1904)
);

AOI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1716),
.B1(n_1709),
.B2(n_1711),
.C(n_1717),
.Y(n_1905)
);

AOI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1625),
.B(n_1567),
.C(n_1711),
.Y(n_1906)
);


endmodule