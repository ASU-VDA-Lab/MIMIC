module fake_jpeg_28707_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_20),
.B1(n_42),
.B2(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_68),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_57),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_19),
.B1(n_39),
.B2(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_50),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_45),
.B(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_56),
.B1(n_59),
.B2(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_85),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_0),
.Y(n_77)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_2),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_18),
.A3(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_14),
.B1(n_30),
.B2(n_29),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_1),
.B(n_2),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_113),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_16),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_7),
.Y(n_132)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_107),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_24),
.C(n_28),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_130),
.A3(n_134),
.B1(n_125),
.B2(n_126),
.C1(n_127),
.C2(n_129),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_140),
.Y(n_144)
);

AOI221xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_116),
.B1(n_115),
.B2(n_114),
.C(n_106),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_115),
.B1(n_133),
.B2(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_142),
.B1(n_131),
.B2(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_141),
.C(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_11),
.B(n_22),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_25),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_26),
.Y(n_152)
);


endmodule