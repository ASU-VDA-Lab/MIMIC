module fake_jpeg_12257_n_380 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_53),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_62),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_3),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_4),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_5),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_37),
.C(n_40),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_21),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_26),
.C(n_32),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_41),
.B1(n_22),
.B2(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_95),
.B1(n_97),
.B2(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_106),
.C(n_46),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_41),
.B1(n_19),
.B2(n_31),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_19),
.B1(n_31),
.B2(n_33),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_33),
.B1(n_40),
.B2(n_27),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_103),
.B1(n_82),
.B2(n_47),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_33),
.B1(n_38),
.B2(n_23),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_100),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_44),
.A2(n_33),
.B1(n_32),
.B2(n_20),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_54),
.B1(n_70),
.B2(n_55),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_80),
.C(n_71),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_49),
.A2(n_20),
.B1(n_32),
.B2(n_38),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_30),
.B(n_28),
.C(n_27),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_110),
.A2(n_128),
.B(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_69),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_32),
.B1(n_20),
.B2(n_26),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_117),
.B1(n_129),
.B2(n_60),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_32),
.B1(n_20),
.B2(n_7),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_20),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_50),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_144),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_151),
.Y(n_210)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_64),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_142),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_45),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_92),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_167),
.B1(n_122),
.B2(n_87),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_51),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_72),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_42),
.B1(n_65),
.B2(n_43),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_174),
.B(n_150),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_56),
.B1(n_46),
.B2(n_78),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_173),
.B1(n_130),
.B2(n_90),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_102),
.Y(n_157)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_159),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_88),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_161),
.C(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_57),
.C(n_48),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_102),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_9),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_166),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_10),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_101),
.A2(n_10),
.B1(n_11),
.B2(n_118),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_10),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_11),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_120),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_124),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_100),
.A2(n_11),
.B1(n_119),
.B2(n_130),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_90),
.B1(n_108),
.B2(n_83),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_205),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_110),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_180),
.B(n_210),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_121),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_171),
.B1(n_136),
.B2(n_138),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_126),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_115),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_131),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_134),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_83),
.B1(n_87),
.B2(n_122),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_201),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_91),
.B1(n_125),
.B2(n_127),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_91),
.A3(n_115),
.B1(n_126),
.B2(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_147),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_137),
.B1(n_154),
.B2(n_174),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_217),
.A2(n_222),
.B1(n_226),
.B2(n_229),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_164),
.B(n_157),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_177),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_221),
.B(n_244),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_149),
.B1(n_143),
.B2(n_139),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_144),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_172),
.C(n_148),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_240),
.C(n_247),
.Y(n_272)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_135),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_241),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_133),
.B1(n_146),
.B2(n_168),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_156),
.B1(n_158),
.B2(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_232),
.A2(n_242),
.B1(n_217),
.B2(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_171),
.B(n_158),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_249),
.B(n_189),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_183),
.A2(n_156),
.B1(n_176),
.B2(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_216),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_243),
.A2(n_247),
.B(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_210),
.C(n_192),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_198),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_248),
.A2(n_219),
.B(n_246),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_192),
.A2(n_210),
.B(n_178),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_235),
.A2(n_199),
.B1(n_205),
.B2(n_193),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_251),
.A2(n_255),
.B1(n_271),
.B2(n_230),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_197),
.B1(n_190),
.B2(n_185),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_177),
.B(n_185),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_258),
.B(n_248),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_182),
.B(n_212),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_196),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_182),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_194),
.A3(n_203),
.B1(n_212),
.B2(n_202),
.C1(n_204),
.C2(n_189),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_262),
.A2(n_269),
.B(n_278),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_202),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_277),
.C(n_222),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_203),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_226),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_203),
.B1(n_234),
.B2(n_220),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_248),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_220),
.C(n_225),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_219),
.B(n_226),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_288),
.B(n_256),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_224),
.B(n_267),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_272),
.C(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_238),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_293),
.B(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_274),
.B(n_245),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_283),
.B1(n_280),
.B2(n_292),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_259),
.B(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_301),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_261),
.B(n_229),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_268),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_268),
.A2(n_227),
.B1(n_280),
.B2(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_317),
.B(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_251),
.B1(n_255),
.B2(n_271),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_296),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_314),
.C(n_316),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_272),
.C(n_263),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_266),
.C(n_275),
.Y(n_316)
);

AOI22x1_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_253),
.B1(n_258),
.B2(n_264),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_296),
.B1(n_297),
.B2(n_287),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_260),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_291),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_326),
.B(n_328),
.Y(n_343)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_281),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_338),
.B1(n_322),
.B2(n_288),
.Y(n_346)
);

OAI322xp33_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_289),
.A3(n_295),
.B1(n_294),
.B2(n_286),
.C1(n_318),
.C2(n_305),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_332),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_333),
.Y(n_345)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_293),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_299),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_337),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_313),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_284),
.C(n_321),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_313),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_312),
.A2(n_282),
.B1(n_303),
.B2(n_300),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_309),
.B1(n_319),
.B2(n_285),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_317),
.B(n_298),
.Y(n_349)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_318),
.CI(n_307),
.CON(n_341),
.SN(n_341)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_344),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_342),
.A2(n_331),
.B1(n_322),
.B2(n_311),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_346),
.A2(n_340),
.B1(n_285),
.B2(n_325),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_340),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_310),
.C(n_316),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_351),
.C(n_301),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_322),
.C(n_298),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_342),
.A2(n_329),
.B1(n_325),
.B2(n_326),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_355),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_356),
.A2(n_359),
.B1(n_349),
.B2(n_341),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_SL g357 ( 
.A(n_351),
.B(n_333),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_360),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_322),
.C(n_337),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_361),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_327),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_355),
.A2(n_348),
.B1(n_347),
.B2(n_344),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_365),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_364),
.Y(n_372)
);

OAI321xp33_ASAP7_75t_L g366 ( 
.A1(n_354),
.A2(n_348),
.A3(n_352),
.B1(n_302),
.B2(n_341),
.C(n_346),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_366),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_358),
.C(n_345),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_369),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_368),
.A3(n_353),
.B1(n_332),
.B2(n_294),
.C1(n_365),
.C2(n_367),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_373),
.Y(n_377)
);

AOI322xp5_ASAP7_75t_L g374 ( 
.A1(n_372),
.A2(n_367),
.A3(n_359),
.B1(n_270),
.B2(n_265),
.C1(n_345),
.C2(n_276),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_374),
.B(n_371),
.C(n_270),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_375),
.C(n_276),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_378),
.B(n_369),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_377),
.Y(n_380)
);


endmodule