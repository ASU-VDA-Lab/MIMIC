module fake_jpeg_16808_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_17),
.B1(n_27),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_63),
.B1(n_68),
.B2(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_31),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_18),
.B1(n_25),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_33),
.B1(n_35),
.B2(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_64),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_33),
.C(n_19),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_34),
.C(n_23),
.Y(n_90)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_33),
.B1(n_34),
.B2(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_25),
.B1(n_21),
.B2(n_30),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_85),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_24),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_29),
.B(n_64),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_59),
.B1(n_51),
.B2(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_57),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_19),
.C(n_63),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_42),
.B1(n_34),
.B2(n_23),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_63),
.B(n_1),
.Y(n_102)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_100),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_63),
.B(n_48),
.C(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

OR2x4_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_75),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_99),
.B1(n_115),
.B2(n_102),
.Y(n_132)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_32),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_81),
.C(n_85),
.Y(n_146)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_78),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_133),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_142),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22x1_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_77),
.B1(n_91),
.B2(n_32),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_104),
.B1(n_116),
.B2(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_86),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_95),
.B(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_115),
.C(n_96),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_156),
.C(n_166),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_96),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_173),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_171),
.B(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_121),
.C(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_102),
.B1(n_99),
.B2(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_117),
.B1(n_111),
.B2(n_93),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_93),
.B1(n_81),
.B2(n_51),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_103),
.B1(n_106),
.B2(n_114),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_80),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_103),
.C(n_82),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_126),
.C(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_103),
.B1(n_106),
.B2(n_114),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_130),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_109),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_135),
.A3(n_129),
.B1(n_125),
.B2(n_136),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_149),
.B(n_170),
.C(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_183),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_170),
.B(n_165),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_193),
.B(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_124),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_188),
.C(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_143),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_132),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_198),
.B1(n_199),
.B2(n_126),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_153),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_135),
.B(n_142),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_120),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_22),
.C(n_20),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_144),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_179),
.A2(n_158),
.B1(n_157),
.B2(n_160),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_157),
.B1(n_159),
.B2(n_150),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_20),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_137),
.B1(n_120),
.B2(n_166),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_211),
.B1(n_220),
.B2(n_195),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_137),
.B1(n_173),
.B2(n_119),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_65),
.B1(n_46),
.B2(n_119),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_213),
.C(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_82),
.C(n_72),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_72),
.C(n_46),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_97),
.C(n_22),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_221),
.C(n_181),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_97),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_22),
.C(n_20),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_209),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_190),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_189),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_175),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_235),
.B(n_205),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_238),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_182),
.B1(n_176),
.B2(n_10),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_239),
.B1(n_219),
.B2(n_11),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_8),
.B(n_14),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_226),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_202),
.B1(n_209),
.B2(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_226),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_213),
.B1(n_217),
.B2(n_212),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_203),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_236),
.C(n_223),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_239),
.B(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_240),
.B1(n_249),
.B2(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_262),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_242),
.B(n_243),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_223),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_8),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_229),
.C(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_251),
.C(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_260),
.B1(n_256),
.B2(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_273),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_3),
.B(n_5),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_3),
.B(n_6),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_3),
.C(n_7),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_260),
.B1(n_259),
.B2(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_279),
.C(n_9),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_269),
.A3(n_267),
.B1(n_275),
.B2(n_266),
.C1(n_11),
.C2(n_12),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_283),
.B(n_285),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_7),
.B(n_8),
.Y(n_285)
);

AO221x1_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_287),
.B1(n_278),
.B2(n_14),
.C(n_15),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_281),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_282),
.C(n_276),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_288),
.B(n_12),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_15),
.Y(n_293)
);


endmodule