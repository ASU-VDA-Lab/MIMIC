module fake_jpeg_25894_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_0),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_47),
.C(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_63),
.Y(n_68)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_78),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_64),
.B1(n_61),
.B2(n_60),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_84)
);

OA22x2_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_55),
.B1(n_57),
.B2(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_46),
.B1(n_41),
.B2(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_58),
.B1(n_40),
.B2(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_77),
.B1(n_80),
.B2(n_1),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_56),
.B1(n_41),
.B2(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_39),
.B1(n_48),
.B2(n_45),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_0),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_45),
.B1(n_43),
.B2(n_52),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_71),
.A3(n_78),
.B1(n_43),
.B2(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_51),
.B1(n_20),
.B2(n_22),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_24),
.B1(n_36),
.B2(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_103)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_3),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_3),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_4),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_92),
.B1(n_87),
.B2(n_8),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_84),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_110),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_90),
.C(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_108),
.C(n_100),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_91),
.C(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_113),
.B1(n_98),
.B2(n_104),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_112),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

BUFx12f_ASAP7_75t_SL g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_102),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_23),
.B1(n_30),
.B2(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_82),
.C(n_25),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_129),
.C(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_115),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_116),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_127),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_132),
.B(n_126),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_118),
.C(n_17),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_14),
.Y(n_141)
);


endmodule