module fake_ariane_2291_n_1841 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1841);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1841;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_111),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_47),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_109),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_37),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_83),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_8),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_19),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_18),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_74),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_95),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_26),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_36),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_103),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_11),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_4),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_152),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_134),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_67),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_48),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_35),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_71),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_10),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_92),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_106),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_105),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_53),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_48),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_75),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_52),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_14),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_90),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_6),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_18),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_88),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_101),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_46),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_86),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_40),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_156),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_161),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_96),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_139),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_121),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_160),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_21),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_49),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_82),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_108),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_47),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_42),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_54),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_85),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_100),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_84),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_59),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_31),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_33),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_0),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_87),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_45),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_128),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_11),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_118),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_31),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_141),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_44),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_76),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_113),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_43),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_80),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_81),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_72),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_54),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_94),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_41),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_155),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_40),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_52),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_23),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_19),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_51),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_70),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_32),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_55),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_34),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_28),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_56),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

BUFx8_ASAP7_75t_SL g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_271),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_330),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_184),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_227),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_219),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_231),
.B(n_244),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_0),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_224),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_174),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_247),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_252),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_309),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_316),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_208),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_234),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_216),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_303),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_225),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_252),
.B(n_3),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_246),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_315),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_248),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_187),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_189),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_218),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_221),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_254),
.B(n_6),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_250),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_253),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_257),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_317),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_234),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_189),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_269),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_288),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_171),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_270),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_275),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_7),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_234),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_172),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_277),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_288),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_259),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_231),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_172),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_278),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_244),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_259),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_186),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_174),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_186),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_265),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_265),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_245),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_289),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_193),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_289),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_177),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_182),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_185),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_344),
.B(n_199),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_373),
.B(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_345),
.Y(n_433)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_357),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_204),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_366),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_213),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_400),
.B(n_321),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_374),
.B(n_215),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_351),
.B(n_321),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_328),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_385),
.B(n_226),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_376),
.B(n_239),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_372),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_389),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_240),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_342),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_364),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_404),
.B(n_378),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_390),
.B(n_242),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_355),
.B(n_243),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_348),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_363),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_365),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_368),
.A2(n_260),
.B(n_258),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_375),
.B1(n_377),
.B2(n_339),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_434),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_356),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_356),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_453),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_377),
.B1(n_406),
.B2(n_412),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_484),
.B(n_371),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_464),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_413),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_484),
.B(n_379),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_380),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_434),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_SL g510 ( 
.A(n_484),
.B(n_381),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_387),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_391),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_424),
.A2(n_383),
.B1(n_394),
.B2(n_354),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_486),
.A2(n_408),
.B1(n_407),
.B2(n_405),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_478),
.A2(n_318),
.B1(n_402),
.B2(n_396),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_434),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_432),
.B(n_328),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_392),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_486),
.A2(n_212),
.B1(n_301),
.B2(n_329),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_435),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_166),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_464),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

AND3x2_ASAP7_75t_L g538 ( 
.A(n_467),
.B(n_393),
.C(n_180),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g539 ( 
.A(n_480),
.B(n_194),
.C(n_193),
.Y(n_539)
);

AOI21x1_ASAP7_75t_L g540 ( 
.A1(n_414),
.A2(n_191),
.B(n_178),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_434),
.A2(n_202),
.B1(n_200),
.B2(n_196),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_484),
.B(n_166),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_486),
.A2(n_220),
.B1(n_176),
.B2(n_322),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_484),
.B(n_331),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_441),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_434),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_432),
.B(n_167),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_434),
.B(n_334),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_167),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_434),
.A2(n_297),
.B1(n_196),
.B2(n_200),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_336),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_478),
.A2(n_202),
.B1(n_194),
.B2(n_325),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_481),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_484),
.B(n_350),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_442),
.B(n_352),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_480),
.B(n_168),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_484),
.B(n_168),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_444),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_420),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_245),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_484),
.B(n_169),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_485),
.B(n_169),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_485),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_485),
.B(n_170),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_420),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_444),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_421),
.B(n_206),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_445),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_485),
.B(n_170),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_415),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_486),
.A2(n_223),
.B1(n_195),
.B2(n_320),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_417),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_445),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_437),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_437),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_173),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_445),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_415),
.Y(n_584)
);

AND2x2_ASAP7_75t_SL g585 ( 
.A(n_486),
.B(n_178),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_481),
.B(n_410),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_450),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_414),
.B(n_237),
.C(n_205),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_437),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_450),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_481),
.B(n_476),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_452),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_437),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_479),
.A2(n_281),
.B1(n_296),
.B2(n_292),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_452),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_485),
.B(n_173),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_485),
.B(n_175),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_437),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_421),
.B(n_238),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_457),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_485),
.B(n_175),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_437),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_457),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_437),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_437),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_485),
.B(n_179),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_417),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_457),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_466),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_466),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_479),
.A2(n_241),
.B1(n_290),
.B2(n_312),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_439),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_473),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_481),
.B(n_341),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_481),
.B(n_179),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_181),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_469),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_415),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_439),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_463),
.A2(n_393),
.B1(n_327),
.B2(n_326),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_430),
.B(n_332),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_451),
.B(n_245),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_417),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_430),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_468),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_417),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_554),
.B(n_448),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_596),
.B(n_448),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_631),
.B(n_476),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_528),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_567),
.B(n_448),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_536),
.B(n_482),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_514),
.A2(n_448),
.B1(n_483),
.B2(n_476),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_585),
.A2(n_421),
.B1(n_448),
.B2(n_475),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_448),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_617),
.Y(n_649)
);

OAI221xp5_ASAP7_75t_L g650 ( 
.A1(n_601),
.A2(n_474),
.B1(n_463),
.B2(n_483),
.C(n_319),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_483),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_528),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_567),
.B(n_488),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_514),
.A2(n_430),
.B1(n_474),
.B2(n_454),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_494),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_492),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_488),
.B(n_414),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_567),
.B(n_416),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_493),
.B(n_451),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_558),
.B(n_451),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_618),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_618),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_522),
.B(n_458),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_567),
.B(n_416),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_494),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_492),
.B(n_482),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_532),
.B(n_418),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_522),
.B(n_458),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_593),
.B(n_418),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_458),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_522),
.B(n_418),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_507),
.B(n_416),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_507),
.B(n_418),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_520),
.B(n_418),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_520),
.B(n_418),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_598),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_547),
.A2(n_449),
.B1(n_454),
.B2(n_431),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_547),
.B(n_422),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_549),
.B(n_419),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_598),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_535),
.B(n_419),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_548),
.B(n_419),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_550),
.B(n_419),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_519),
.B(n_306),
.C(n_297),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_633),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_624),
.B(n_419),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_585),
.A2(n_421),
.B1(n_475),
.B2(n_456),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_625),
.A2(n_446),
.B1(n_427),
.B2(n_422),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_487),
.B(n_419),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_498),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_523),
.B(n_422),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_556),
.B(n_436),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_482),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_614),
.B(n_436),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_623),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_585),
.A2(n_421),
.B1(n_475),
.B2(n_456),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_584),
.B(n_456),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_495),
.B(n_436),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_627),
.B(n_456),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_627),
.B(n_456),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_634),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_633),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_490),
.B(n_427),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_503),
.B(n_504),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_635),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_523),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_523),
.B(n_427),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_568),
.B(n_433),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_503),
.B(n_436),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_635),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_573),
.A2(n_440),
.B1(n_433),
.B2(n_443),
.Y(n_718)
);

AND2x6_ASAP7_75t_L g719 ( 
.A(n_598),
.B(n_421),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_503),
.B(n_504),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_503),
.B(n_436),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_573),
.A2(n_433),
.B1(n_440),
.B2(n_443),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_634),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_568),
.B(n_440),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_568),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_636),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_504),
.B(n_508),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_499),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_578),
.B(n_443),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_636),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_489),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_489),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_502),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_629),
.A2(n_324),
.B1(n_310),
.B2(n_325),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_497),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_504),
.B(n_436),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_637),
.B(n_438),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_497),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_508),
.B(n_438),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_552),
.B(n_557),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_578),
.B(n_438),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_578),
.B(n_446),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_637),
.B(n_438),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_576),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_490),
.B(n_446),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_490),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_500),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_508),
.B(n_438),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_508),
.B(n_438),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_447),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_637),
.B(n_447),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_588),
.B(n_449),
.C(n_431),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_632),
.B(n_447),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_533),
.A2(n_456),
.B1(n_473),
.B2(n_428),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_563),
.B(n_500),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_509),
.B(n_511),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_539),
.A2(n_455),
.B1(n_203),
.B2(n_299),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_538),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_632),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_347),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_573),
.A2(n_455),
.B1(n_203),
.B2(n_299),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_502),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_543),
.A2(n_473),
.B1(n_426),
.B2(n_428),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_509),
.B(n_455),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_511),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_525),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_629),
.B(n_353),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_505),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_505),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_521),
.Y(n_770)
);

AND2x6_ASAP7_75t_SL g771 ( 
.A(n_606),
.B(n_360),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_525),
.B(n_426),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_630),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_516),
.A2(n_191),
.B1(n_382),
.B2(n_369),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_506),
.B(n_310),
.C(n_327),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_530),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_SL g777 ( 
.A(n_632),
.B(n_306),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_606),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_573),
.A2(n_201),
.B1(n_197),
.B2(n_323),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_530),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_490),
.B(n_439),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_515),
.B(n_362),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_577),
.A2(n_473),
.B1(n_461),
.B2(n_470),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_606),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_531),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_496),
.B(n_473),
.Y(n_786)
);

XOR2xp5_ASAP7_75t_L g787 ( 
.A(n_541),
.B(n_181),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_531),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_590),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_501),
.B(n_439),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_324),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_560),
.B(n_439),
.Y(n_792)
);

AO22x2_ASAP7_75t_L g793 ( 
.A1(n_590),
.A2(n_461),
.B1(n_262),
.B2(n_263),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_521),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_490),
.B(n_439),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_553),
.B(n_326),
.C(n_294),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_560),
.B(n_439),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_541),
.B(n_439),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_529),
.B(n_600),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_529),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_573),
.B(n_473),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_551),
.A2(n_473),
.B1(n_470),
.B2(n_468),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_561),
.B(n_439),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_529),
.B(n_473),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_561),
.B(n_473),
.Y(n_806)
);

AND2x2_ASAP7_75t_SL g807 ( 
.A(n_542),
.B(n_261),
.Y(n_807)
);

AO21x1_ASAP7_75t_L g808 ( 
.A1(n_638),
.A2(n_510),
.B(n_559),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_702),
.B(n_551),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_686),
.A2(n_639),
.B(n_693),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_686),
.A2(n_582),
.B(n_565),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_649),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_656),
.Y(n_813)
);

AND2x6_ASAP7_75t_L g814 ( 
.A(n_802),
.B(n_566),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_661),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_740),
.B(n_708),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_664),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_716),
.A2(n_608),
.B(n_604),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_697),
.B(n_566),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_713),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_677),
.B(n_571),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_721),
.A2(n_613),
.B(n_569),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_736),
.A2(n_575),
.B(n_564),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_739),
.A2(n_603),
.B(n_621),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_579),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_771),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_647),
.A2(n_579),
.B1(n_583),
.B2(n_594),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_800),
.A2(n_594),
.B(n_583),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_792),
.A2(n_540),
.B(n_527),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_657),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_713),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_662),
.B(n_607),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_748),
.A2(n_621),
.B(n_518),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_647),
.A2(n_646),
.B1(n_692),
.B2(n_665),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_713),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_778),
.B(n_545),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_749),
.A2(n_621),
.B(n_518),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_641),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_709),
.A2(n_610),
.B1(n_537),
.B2(n_602),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_712),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_744),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_640),
.B(n_524),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_773),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_641),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_799),
.A2(n_527),
.B(n_524),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_670),
.B(n_512),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_711),
.A2(n_518),
.B(n_512),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_784),
.B(n_529),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_767),
.Y(n_850)
);

AND2x6_ASAP7_75t_L g851 ( 
.A(n_717),
.B(n_534),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_750),
.B(n_534),
.Y(n_852)
);

NOR3xp33_ASAP7_75t_L g853 ( 
.A(n_734),
.B(n_283),
.C(n_279),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_651),
.B(n_537),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_720),
.A2(n_518),
.B(n_512),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_727),
.A2(n_544),
.B(n_512),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_723),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_755),
.B(n_555),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_671),
.Y(n_859)
);

NOR2x1p5_ASAP7_75t_L g860 ( 
.A(n_760),
.B(n_293),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_671),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_672),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_640),
.B(n_555),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_799),
.A2(n_574),
.B(n_572),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_800),
.A2(n_562),
.B(n_544),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_734),
.A2(n_599),
.B1(n_595),
.B2(n_602),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_648),
.B(n_654),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_689),
.A2(n_574),
.B(n_572),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_645),
.B(n_544),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_700),
.B(n_586),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_672),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_673),
.A2(n_586),
.B(n_599),
.C(n_595),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_691),
.A2(n_615),
.B(n_616),
.C(n_589),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_795),
.B(n_529),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_642),
.A2(n_562),
.B(n_597),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_689),
.A2(n_587),
.B(n_589),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_642),
.A2(n_544),
.B(n_597),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_789),
.B(n_562),
.Y(n_878)
);

NOR2x1p5_ASAP7_75t_SL g879 ( 
.A(n_676),
.B(n_587),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_726),
.B(n_615),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_677),
.B(n_562),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_719),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_688),
.A2(n_611),
.B(n_597),
.Y(n_883)
);

INVx11_ASAP7_75t_L g884 ( 
.A(n_719),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_659),
.A2(n_667),
.B(n_658),
.Y(n_885)
);

NAND2x2_ASAP7_75t_L g886 ( 
.A(n_758),
.B(n_706),
.Y(n_886)
);

AO21x1_ASAP7_75t_L g887 ( 
.A1(n_718),
.A2(n_540),
.B(n_616),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_782),
.B(n_597),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_713),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_622),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_650),
.A2(n_626),
.B(n_622),
.C(n_609),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_673),
.B(n_626),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_656),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_659),
.A2(n_667),
.B(n_701),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_669),
.B(n_611),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_722),
.A2(n_611),
.B(n_612),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_801),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_761),
.B(n_600),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_757),
.B(n_611),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_798),
.A2(n_612),
.B(n_526),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_678),
.A2(n_609),
.B(n_605),
.C(n_581),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_804),
.A2(n_526),
.B(n_580),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_756),
.A2(n_682),
.B(n_681),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_690),
.A2(n_581),
.B(n_517),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_704),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_797),
.A2(n_517),
.B(n_609),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_707),
.B(n_612),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_666),
.B(n_612),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_676),
.Y(n_909)
);

NOR2x1_ASAP7_75t_L g910 ( 
.A(n_752),
.B(n_517),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_674),
.B(n_517),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_690),
.A2(n_526),
.B(n_570),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_675),
.B(n_526),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_704),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_704),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_772),
.A2(n_570),
.B(n_580),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_684),
.A2(n_580),
.B1(n_609),
.B2(n_605),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_675),
.B(n_570),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_801),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_787),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_751),
.B(n_570),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_731),
.B(n_580),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_751),
.A2(n_581),
.B(n_605),
.C(n_470),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_764),
.A2(n_605),
.B(n_581),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_699),
.A2(n_268),
.B(n_291),
.C(n_282),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_807),
.A2(n_600),
.B1(n_620),
.B2(n_628),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_698),
.A2(n_272),
.B(n_305),
.C(n_469),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_669),
.B(n_600),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_680),
.A2(n_600),
.B(n_620),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_680),
.A2(n_628),
.B(n_620),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_728),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_781),
.A2(n_628),
.B(n_620),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_732),
.B(n_592),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_694),
.B(n_703),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_699),
.A2(n_471),
.B(n_469),
.C(n_472),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_781),
.A2(n_628),
.B(n_620),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_759),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_779),
.A2(n_741),
.B(n_737),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_725),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_759),
.B(n_643),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_694),
.B(n_703),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_695),
.A2(n_628),
.B(n_620),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_805),
.A2(n_471),
.B(n_472),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_643),
.B(n_592),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_719),
.B(n_592),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_801),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_746),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_733),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_719),
.B(n_592),
.Y(n_950)
);

AO21x2_ASAP7_75t_L g951 ( 
.A1(n_696),
.A2(n_705),
.B(n_790),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_735),
.Y(n_952)
);

CKINVDCx10_ASAP7_75t_R g953 ( 
.A(n_774),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_719),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_653),
.A2(n_628),
.B(n_592),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_737),
.B(n_592),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_777),
.A2(n_653),
.B(n_679),
.C(n_685),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_741),
.A2(n_183),
.B(n_323),
.Y(n_958)
);

CKINVDCx8_ASAP7_75t_R g959 ( 
.A(n_746),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_725),
.B(n_183),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_806),
.A2(n_462),
.B(n_459),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_738),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_807),
.B(n_190),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_747),
.B(n_471),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_743),
.A2(n_714),
.B(n_698),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_746),
.B(n_462),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_743),
.A2(n_796),
.B(n_715),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_765),
.B(n_471),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_746),
.B(n_801),
.Y(n_969)
);

NOR2x1_ASAP7_75t_L g970 ( 
.A(n_714),
.B(n_462),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_791),
.B(n_190),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_786),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_715),
.A2(n_192),
.B(n_197),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_803),
.B(n_462),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_724),
.A2(n_472),
.B(n_459),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_754),
.B(n_192),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_754),
.B(n_201),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_724),
.A2(n_295),
.B(n_298),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_766),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_733),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_803),
.Y(n_981)
);

NAND2x1_ASAP7_75t_L g982 ( 
.A(n_768),
.B(n_462),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_768),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_729),
.A2(n_295),
.B(n_298),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_SL g985 ( 
.A1(n_679),
.A2(n_472),
.B(n_459),
.C(n_462),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_729),
.A2(n_459),
.B(n_304),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_774),
.B(n_793),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_685),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_776),
.B(n_302),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_774),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_742),
.A2(n_302),
.B1(n_304),
.B2(n_314),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_793),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_742),
.A2(n_307),
.B(n_311),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_753),
.B(n_307),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_780),
.A2(n_314),
.B(n_313),
.C(n_311),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_785),
.B(n_313),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_753),
.A2(n_249),
.B(n_209),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_809),
.B(n_788),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_971),
.B(n_775),
.Y(n_999)
);

AOI222xp33_ASAP7_75t_L g1000 ( 
.A1(n_934),
.A2(n_941),
.B1(n_821),
.B2(n_981),
.C1(n_920),
.C2(n_850),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_959),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_853),
.A2(n_793),
.B1(n_790),
.B2(n_745),
.Y(n_1002)
);

BUFx8_ASAP7_75t_L g1003 ( 
.A(n_819),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_835),
.A2(n_763),
.B1(n_783),
.B2(n_644),
.C(n_655),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_931),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_847),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_810),
.A2(n_805),
.B(n_710),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_943),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_811),
.A2(n_652),
.B(n_660),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_812),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_818),
.A2(n_668),
.B(n_683),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_899),
.A2(n_786),
.B1(n_687),
.B2(n_763),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_949),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_897),
.Y(n_1014)
);

BUFx8_ASAP7_75t_SL g1015 ( 
.A(n_844),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_SL g1016 ( 
.A(n_882),
.B(n_762),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_815),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_892),
.A2(n_823),
.B(n_867),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_905),
.B(n_769),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_831),
.B(n_770),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_842),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_993),
.A2(n_794),
.B(n_783),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_827),
.B(n_207),
.Y(n_1023)
);

NOR2xp67_ASAP7_75t_SL g1024 ( 
.A(n_882),
.B(n_210),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_884),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_888),
.B(n_211),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_857),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_938),
.A2(n_465),
.B(n_460),
.C(n_285),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_983),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_835),
.A2(n_255),
.B1(n_217),
.B2(n_284),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_987),
.A2(n_465),
.B1(n_460),
.B2(n_280),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_878),
.A2(n_465),
.B(n_460),
.C(n_276),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_817),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_914),
.B(n_214),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_822),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_843),
.B(n_841),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_882),
.B(n_460),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_961),
.A2(n_460),
.B(n_465),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_952),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_808),
.A2(n_465),
.B(n_15),
.C(n_16),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_940),
.B(n_460),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_816),
.B(n_222),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_944),
.A2(n_460),
.B(n_465),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_925),
.A2(n_465),
.B(n_460),
.C(n_274),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_826),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_886),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_902),
.A2(n_251),
.B(n_229),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_826),
.A2(n_13),
.B(n_17),
.C(n_20),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_860),
.B(n_17),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_839),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_915),
.B(n_20),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_897),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_881),
.B(n_26),
.Y(n_1054)
);

BUFx12f_ASAP7_75t_L g1055 ( 
.A(n_820),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_907),
.A2(n_256),
.B1(n_232),
.B2(n_273),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_892),
.A2(n_460),
.B(n_465),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_962),
.B(n_27),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_979),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_963),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_870),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_992),
.B(n_30),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_882),
.B(n_267),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_921),
.A2(n_465),
.B(n_264),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_820),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_869),
.A2(n_236),
.B(n_235),
.C(n_228),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_863),
.B(n_34),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_948),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_854),
.B(n_35),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_814),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_833),
.B(n_36),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_880),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_880),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_845),
.Y(n_1074)
);

CKINVDCx10_ASAP7_75t_R g1075 ( 
.A(n_953),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_38),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_903),
.A2(n_38),
.B(n_42),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_965),
.A2(n_44),
.B(n_45),
.C(n_49),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_912),
.A2(n_50),
.B(n_53),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_940),
.B(n_55),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_859),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_846),
.A2(n_102),
.B(n_57),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_834),
.A2(n_838),
.B(n_883),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_994),
.B(n_56),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_873),
.A2(n_61),
.B(n_66),
.C(n_68),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_956),
.A2(n_69),
.B(n_78),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_954),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_939),
.A2(n_79),
.B1(n_93),
.B2(n_97),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_904),
.A2(n_99),
.B(n_114),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_990),
.A2(n_117),
.B1(n_120),
.B2(n_126),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_814),
.B(n_131),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_814),
.B(n_140),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_814),
.A2(n_977),
.B1(n_976),
.B2(n_993),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_960),
.A2(n_143),
.B(n_148),
.C(n_150),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_965),
.A2(n_154),
.B(n_162),
.C(n_852),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_820),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_891),
.A2(n_906),
.B(n_957),
.C(n_894),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_830),
.A2(n_829),
.B(n_864),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_885),
.A2(n_972),
.B(n_901),
.C(n_967),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_861),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_937),
.B(n_813),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_937),
.B(n_813),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_904),
.A2(n_848),
.B(n_855),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_989),
.B(n_996),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_856),
.A2(n_916),
.B(n_824),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_928),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_832),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_846),
.A2(n_864),
.B(n_877),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_862),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_871),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_897),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_893),
.B(n_995),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_893),
.B(n_832),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_858),
.B(n_988),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_991),
.B(n_874),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_972),
.A2(n_926),
.B(n_879),
.C(n_986),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_SL g1117 ( 
.A1(n_926),
.A2(n_890),
.B(n_942),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_889),
.B(n_948),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_889),
.B(n_928),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_909),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_832),
.B(n_836),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_919),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_SL g1123 ( 
.A(n_958),
.B(n_984),
.C(n_978),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_923),
.A2(n_840),
.B(n_828),
.C(n_872),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_980),
.B(n_911),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_966),
.B(n_836),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_908),
.A2(n_918),
.B(n_913),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_836),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_828),
.A2(n_922),
.B1(n_840),
.B2(n_895),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_935),
.A2(n_968),
.B(n_964),
.C(n_917),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_825),
.A2(n_875),
.B(n_900),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_922),
.A2(n_895),
.B1(n_968),
.B2(n_964),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_980),
.B(n_851),
.Y(n_1133)
);

INVx5_ASAP7_75t_L g1134 ( 
.A(n_851),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_919),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_974),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_SL g1137 ( 
.A(n_919),
.B(n_947),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_924),
.A2(n_865),
.B(n_876),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_851),
.B(n_866),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_986),
.A2(n_910),
.B(n_927),
.C(n_876),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_982),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_970),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_966),
.B(n_946),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_951),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_917),
.A2(n_868),
.B(n_898),
.C(n_985),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_L g1146 ( 
.A1(n_896),
.A2(n_887),
.B(n_837),
.C(n_945),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_947),
.B(n_950),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_868),
.A2(n_942),
.B(n_929),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_947),
.B(n_973),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_997),
.B(n_933),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_933),
.A2(n_930),
.B(n_936),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_851),
.B(n_951),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1026),
.A2(n_975),
.B(n_955),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1060),
.A2(n_975),
.B1(n_849),
.B2(n_969),
.C(n_932),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1025),
.B(n_1036),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_1148),
.B(n_1097),
.Y(n_1156)
);

AOI221x1_ASAP7_75t_L g1157 ( 
.A1(n_1077),
.A2(n_1030),
.B1(n_1089),
.B2(n_1079),
.C(n_999),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1148),
.A2(n_1151),
.A3(n_1132),
.B(n_1138),
.Y(n_1158)
);

OAI22x1_ASAP7_75t_L g1159 ( 
.A1(n_998),
.A2(n_1084),
.B1(n_1002),
.B2(n_1050),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1001),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1061),
.B(n_1104),
.Y(n_1161)
);

AND2x2_ASAP7_75t_SL g1162 ( 
.A(n_1019),
.B(n_1001),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1003),
.A2(n_1021),
.B1(n_1000),
.B2(n_1006),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1117),
.A2(n_1129),
.B(n_1103),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1015),
.Y(n_1165)
);

BUFx8_ASAP7_75t_SL g1166 ( 
.A(n_1001),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1010),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1027),
.A2(n_1054),
.B1(n_1093),
.B2(n_1071),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1070),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1146),
.A2(n_1140),
.B(n_1018),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1034),
.B(n_1037),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1018),
.A2(n_1067),
.B(n_1127),
.Y(n_1172)
);

INVx8_ASAP7_75t_L g1173 ( 
.A(n_1055),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1078),
.A2(n_1115),
.B(n_1095),
.C(n_1112),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1012),
.A2(n_1088),
.A3(n_1078),
.B1(n_1047),
.B2(n_1056),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1103),
.A2(n_1083),
.B(n_1105),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1072),
.B(n_1073),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_1099),
.A2(n_1094),
.B(n_1066),
.C(n_1069),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1083),
.A2(n_1105),
.B(n_1131),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_1035),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1116),
.A2(n_1102),
.B(n_1101),
.C(n_1149),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1138),
.A2(n_1131),
.B(n_1098),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1064),
.A2(n_1151),
.B(n_1057),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_1076),
.A2(n_1058),
.B(n_1150),
.C(n_1032),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1064),
.A2(n_1057),
.A3(n_1028),
.B(n_1011),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1005),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_1011),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1106),
.Y(n_1189)
);

OAI22x1_ASAP7_75t_L g1190 ( 
.A1(n_1070),
.A2(n_1062),
.B1(n_1080),
.B2(n_1040),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1048),
.A2(n_1007),
.B(n_1009),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1130),
.A2(n_1124),
.B(n_1145),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1126),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1130),
.A2(n_1124),
.B(n_1145),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1007),
.A2(n_1041),
.B(n_1108),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1017),
.B(n_1033),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1060),
.A2(n_1049),
.B(n_1046),
.C(n_1077),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1009),
.A2(n_1045),
.A3(n_1089),
.B(n_1085),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1059),
.B(n_1136),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1008),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1139),
.A2(n_1125),
.B(n_1114),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1013),
.A2(n_1029),
.B1(n_1100),
.B2(n_1074),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1075),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1091),
.A2(n_1092),
.B(n_1113),
.C(n_1063),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1095),
.A2(n_1049),
.B(n_1046),
.C(n_1022),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1079),
.A2(n_1052),
.B(n_1123),
.C(n_1087),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1025),
.B(n_1126),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1023),
.B(n_1090),
.C(n_1086),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1119),
.B1(n_1143),
.B2(n_1043),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1051),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1119),
.B(n_1109),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1096),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1107),
.B(n_1128),
.Y(n_1213)
);

AOI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1086),
.A2(n_1141),
.B1(n_1068),
.B2(n_1142),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1065),
.B(n_1143),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1081),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1134),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1110),
.A2(n_1120),
.A3(n_1133),
.B(n_1048),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1121),
.A2(n_1135),
.B1(n_1068),
.B2(n_1014),
.C(n_1122),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1134),
.A2(n_1004),
.B(n_1082),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1135),
.B(n_1053),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1134),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1014),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1014),
.B(n_1111),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1143),
.A2(n_1042),
.B1(n_1004),
.B2(n_1118),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1042),
.A2(n_1134),
.B1(n_1016),
.B2(n_1082),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1137),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1053),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1053),
.Y(n_1229)
);

AOI221x1_ASAP7_75t_L g1230 ( 
.A1(n_1111),
.A2(n_1122),
.B1(n_1038),
.B2(n_1031),
.C(n_1024),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1111),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1147),
.A2(n_1038),
.A3(n_1042),
.B(n_1122),
.Y(n_1232)
);

AND2x6_ASAP7_75t_L g1233 ( 
.A(n_1042),
.B(n_1136),
.Y(n_1233)
);

AOI31xp67_ASAP7_75t_L g1234 ( 
.A1(n_1042),
.A2(n_1150),
.A3(n_1149),
.B(n_1002),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1010),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1026),
.A2(n_740),
.B(n_554),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1015),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_999),
.A2(n_740),
.B(n_998),
.C(n_554),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_998),
.A2(n_787),
.B1(n_809),
.B2(n_629),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_999),
.B(n_740),
.C(n_557),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1026),
.A2(n_740),
.B(n_554),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_999),
.A2(n_740),
.B(n_998),
.C(n_554),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1070),
.B(n_702),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_998),
.B(n_702),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_999),
.A2(n_740),
.B(n_998),
.C(n_554),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1025),
.B(n_1036),
.Y(n_1248)
);

AOI31xp67_ASAP7_75t_L g1249 ( 
.A1(n_1150),
.A2(n_1149),
.A3(n_1002),
.B(n_1147),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1070),
.B(n_1025),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1010),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1070),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1021),
.B(n_697),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1070),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1005),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1010),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1021),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1005),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_998),
.B(n_702),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1070),
.B(n_1025),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1006),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1010),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1136),
.B(n_1119),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_999),
.A2(n_740),
.B(n_998),
.C(n_554),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_998),
.B(n_702),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1277)
);

OAI22x1_ASAP7_75t_L g1278 ( 
.A1(n_998),
.A2(n_787),
.B1(n_809),
.B2(n_629),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_999),
.A2(n_740),
.B(n_998),
.C(n_554),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_998),
.B(n_702),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_999),
.A2(n_552),
.B(n_557),
.C(n_740),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1003),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1020),
.B(n_697),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1026),
.A2(n_740),
.B(n_554),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1020),
.B(n_697),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_998),
.B(n_702),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1289)
);

BUFx2_ASAP7_75t_R g1290 ( 
.A(n_1015),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_998),
.B(n_702),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1015),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1039),
.A2(n_1098),
.B(n_1044),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_SL g1297 ( 
.A(n_1070),
.B(n_584),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1015),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1000),
.A2(n_767),
.B1(n_774),
.B2(n_782),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1144),
.A2(n_1152),
.A3(n_808),
.B(n_1148),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1015),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1010),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1021),
.B(n_697),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1010),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1148),
.A2(n_810),
.B(n_638),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1015),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_999),
.A2(n_702),
.B1(n_740),
.B2(n_552),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1246),
.B(n_1264),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1173),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1275),
.A2(n_1281),
.B1(n_1291),
.B2(n_1288),
.Y(n_1311)
);

CKINVDCx12_ASAP7_75t_R g1312 ( 
.A(n_1254),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1292),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1298),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1196),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_1242),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1159),
.A2(n_1208),
.B1(n_1168),
.B2(n_1192),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1173),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1167),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1155),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1161),
.B(n_1285),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1162),
.A2(n_1243),
.B1(n_1238),
.B2(n_1286),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1237),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1308),
.A2(n_1247),
.B1(n_1274),
.B2(n_1240),
.Y(n_1324)
);

CKINVDCx6p67_ASAP7_75t_R g1325 ( 
.A(n_1239),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1301),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1194),
.A2(n_1287),
.B1(n_1172),
.B2(n_1271),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1273),
.A2(n_1177),
.B1(n_1220),
.B2(n_1190),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1307),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1223),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1189),
.B(n_1304),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1244),
.A2(n_1280),
.B1(n_1282),
.B2(n_1174),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1273),
.A2(n_1171),
.B1(n_1305),
.B2(n_1303),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1251),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1273),
.A2(n_1233),
.B1(n_1180),
.B2(n_1170),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1205),
.A2(n_1164),
.B1(n_1225),
.B2(n_1197),
.Y(n_1336)
);

BUFx2_ASAP7_75t_SL g1337 ( 
.A(n_1248),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1229),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1176),
.A2(n_1179),
.B(n_1195),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1248),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1261),
.A2(n_1272),
.B1(n_1201),
.B2(n_1216),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1210),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1166),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1203),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1186),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1165),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1245),
.A2(n_1209),
.B1(n_1153),
.B2(n_1226),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1160),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1157),
.A2(n_1212),
.B1(n_1230),
.B2(n_1193),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1233),
.A2(n_1180),
.B1(n_1211),
.B2(n_1175),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1233),
.A2(n_1259),
.B1(n_1263),
.B2(n_1202),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1228),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1193),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1233),
.A2(n_1215),
.B1(n_1213),
.B2(n_1175),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1175),
.A2(n_1297),
.B1(n_1252),
.B2(n_1258),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1169),
.A2(n_1258),
.B1(n_1252),
.B2(n_1187),
.Y(n_1357)
);

OAI22x1_ASAP7_75t_L g1358 ( 
.A1(n_1214),
.A2(n_1227),
.B1(n_1207),
.B2(n_1222),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1169),
.A2(n_1187),
.B1(n_1222),
.B2(n_1217),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1221),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1217),
.A2(n_1269),
.B1(n_1250),
.B2(n_1234),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1231),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1206),
.A2(n_1306),
.B1(n_1302),
.B2(n_1236),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1224),
.A2(n_1154),
.B1(n_1184),
.B2(n_1178),
.Y(n_1364)
);

CKINVDCx8_ASAP7_75t_R g1365 ( 
.A(n_1231),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_SL g1366 ( 
.A(n_1290),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1218),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1219),
.B(n_1232),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1183),
.A2(n_1276),
.B1(n_1267),
.B2(n_1253),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1266),
.A2(n_1270),
.B1(n_1279),
.B2(n_1182),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1182),
.A2(n_1249),
.B1(n_1198),
.B2(n_1188),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1181),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1198),
.A2(n_1284),
.B1(n_1296),
.B2(n_1257),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1232),
.B(n_1156),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1204),
.A2(n_1294),
.B1(n_1268),
.B2(n_1260),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1156),
.Y(n_1376)
);

BUFx4f_ASAP7_75t_L g1377 ( 
.A(n_1255),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1191),
.B(n_1256),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1265),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1198),
.A2(n_1185),
.B1(n_1277),
.B2(n_1289),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1158),
.A2(n_1185),
.B(n_1277),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1158),
.A2(n_1185),
.B1(n_1300),
.B2(n_1293),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1289),
.A2(n_1293),
.B1(n_1295),
.B2(n_1300),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1289),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1158),
.A2(n_1293),
.B1(n_1295),
.B2(n_1300),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1295),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1166),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1262),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1246),
.A2(n_1275),
.B1(n_1281),
.B2(n_1264),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1199),
.Y(n_1390)
);

CKINVDCx14_ASAP7_75t_R g1391 ( 
.A(n_1203),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1173),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1239),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1166),
.Y(n_1397)
);

BUFx10_ASAP7_75t_L g1398 ( 
.A(n_1292),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1254),
.Y(n_1401)
);

BUFx2_ASAP7_75t_R g1402 ( 
.A(n_1166),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1174),
.A2(n_1006),
.B(n_1271),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1199),
.Y(n_1404)
);

BUFx8_ASAP7_75t_L g1405 ( 
.A(n_1283),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1246),
.A2(n_1264),
.B1(n_1281),
.B2(n_1275),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1199),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1408)
);

BUFx8_ASAP7_75t_SL g1409 ( 
.A(n_1203),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1173),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1262),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1189),
.Y(n_1414)
);

BUFx4f_ASAP7_75t_L g1415 ( 
.A(n_1173),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1193),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1193),
.Y(n_1417)
);

CKINVDCx6p67_ASAP7_75t_R g1418 ( 
.A(n_1239),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1223),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1199),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1308),
.A2(n_1282),
.B(n_1242),
.Y(n_1421)
);

INVx6_ASAP7_75t_L g1422 ( 
.A(n_1173),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1189),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1246),
.A2(n_1264),
.B1(n_1281),
.B2(n_1275),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1285),
.B(n_1287),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1199),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1241),
.A2(n_1278),
.B1(n_1299),
.B2(n_774),
.Y(n_1428)
);

OAI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1163),
.A2(n_1308),
.B1(n_702),
.B2(n_787),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1173),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1235),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1199),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1199),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1379),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1311),
.B(n_1406),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1374),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1384),
.Y(n_1437)
);

INVxp33_ASAP7_75t_L g1438 ( 
.A(n_1426),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1315),
.B(n_1321),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1320),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1319),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1363),
.A2(n_1370),
.B(n_1378),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1323),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1334),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1414),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1429),
.A2(n_1389),
.B1(n_1421),
.B2(n_1425),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1327),
.B(n_1385),
.Y(n_1448)
);

CKINVDCx6p67_ASAP7_75t_R g1449 ( 
.A(n_1345),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1381),
.A2(n_1382),
.B(n_1367),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_R g1451 ( 
.A(n_1387),
.B(n_1397),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1409),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1378),
.A2(n_1369),
.B(n_1373),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1423),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1360),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1332),
.A2(n_1324),
.B(n_1358),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1369),
.A2(n_1373),
.B(n_1371),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1309),
.B(n_1338),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1372),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1353),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1371),
.A2(n_1375),
.B(n_1380),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1380),
.A2(n_1339),
.B(n_1376),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1339),
.A2(n_1336),
.B(n_1383),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1327),
.B(n_1368),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1339),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1331),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1383),
.A2(n_1431),
.B(n_1356),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1377),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1317),
.A2(n_1328),
.B(n_1356),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1392),
.A2(n_1393),
.B1(n_1394),
.B2(n_1413),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1348),
.A2(n_1364),
.B(n_1317),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_R g1472 ( 
.A1(n_1366),
.A2(n_1388),
.B(n_1411),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1401),
.B(n_1341),
.Y(n_1473)
);

BUFx4f_ASAP7_75t_SL g1474 ( 
.A(n_1313),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1340),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1322),
.A2(n_1316),
.B1(n_1392),
.B2(n_1408),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1342),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1362),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1343),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1355),
.B(n_1341),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1386),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1403),
.B(n_1337),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1346),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1359),
.A2(n_1328),
.B(n_1357),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1393),
.A2(n_1400),
.B1(n_1413),
.B2(n_1428),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1390),
.B(n_1433),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1404),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1355),
.B(n_1351),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1350),
.A2(n_1432),
.B(n_1420),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1407),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1427),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1365),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1333),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1333),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1422),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1361),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1357),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1330),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1335),
.B(n_1352),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1416),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1359),
.B(n_1419),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1352),
.A2(n_1394),
.B(n_1399),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1399),
.A2(n_1428),
.B(n_1424),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1417),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1417),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1417),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1354),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1354),
.B(n_1424),
.Y(n_1508)
);

OAI31xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1400),
.A2(n_1408),
.A3(n_1412),
.B(n_1366),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.B(n_1412),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1447),
.A2(n_1312),
.B1(n_1349),
.B2(n_1422),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1466),
.B(n_1344),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1454),
.Y(n_1513)
);

OAI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1435),
.A2(n_1344),
.B(n_1347),
.C(n_1410),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1460),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1468),
.B(n_1430),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1455),
.B(n_1405),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1443),
.A2(n_1463),
.B(n_1457),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_SL g1519 ( 
.A1(n_1459),
.A2(n_1410),
.B(n_1318),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1438),
.B(n_1430),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1446),
.B(n_1310),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1446),
.B(n_1310),
.Y(n_1522)
);

CKINVDCx16_ASAP7_75t_R g1523 ( 
.A(n_1451),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1441),
.B(n_1418),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_1396),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1471),
.A2(n_1415),
.B(n_1395),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1459),
.A2(n_1415),
.B1(n_1402),
.B2(n_1325),
.Y(n_1527)
);

INVxp33_ASAP7_75t_L g1528 ( 
.A(n_1458),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1459),
.B(n_1405),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1440),
.B(n_1314),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_SL g1531 ( 
.A1(n_1498),
.A2(n_1495),
.B(n_1472),
.C(n_1476),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1465),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1476),
.A2(n_1313),
.B1(n_1329),
.B2(n_1391),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1440),
.B(n_1326),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1501),
.B(n_1326),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1464),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1473),
.B(n_1398),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1471),
.A2(n_1398),
.B(n_1456),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1459),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_SL g1540 ( 
.A(n_1482),
.B(n_1492),
.Y(n_1540)
);

OAI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1448),
.A2(n_1456),
.B(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1477),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1485),
.A2(n_1502),
.B1(n_1503),
.B2(n_1470),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1482),
.A2(n_1443),
.B(n_1448),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_SL g1545 ( 
.A(n_1482),
.B(n_1492),
.Y(n_1545)
);

A2O1A1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1509),
.A2(n_1488),
.B(n_1499),
.C(n_1480),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1457),
.A2(n_1453),
.B(n_1461),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1478),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1444),
.B(n_1445),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1482),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1475),
.B(n_1481),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1475),
.B(n_1481),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1436),
.B(n_1479),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1442),
.B(n_1436),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1479),
.B(n_1497),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1453),
.A2(n_1461),
.B(n_1462),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1488),
.A2(n_1480),
.B1(n_1469),
.B2(n_1485),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1507),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1469),
.A2(n_1494),
.B1(n_1493),
.B2(n_1496),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1504),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1486),
.A2(n_1489),
.B1(n_1434),
.B2(n_1491),
.C(n_1487),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1442),
.B(n_1500),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1469),
.A2(n_1504),
.B(n_1506),
.C(n_1505),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1483),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1513),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1560),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1563),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1567),
.B(n_1450),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1542),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1519),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1546),
.A2(n_1502),
.B1(n_1508),
.B2(n_1484),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1565),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1518),
.B(n_1556),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1518),
.B(n_1450),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1518),
.B(n_1556),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1566),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1565),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1568),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1587)
);

NOR2x1p5_ASAP7_75t_L g1588 ( 
.A(n_1548),
.B(n_1449),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1450),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1543),
.A2(n_1502),
.B1(n_1508),
.B2(n_1489),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1550),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1550),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1489),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

NAND4xp25_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1533),
.C(n_1531),
.D(n_1538),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1576),
.A2(n_1543),
.B1(n_1559),
.B2(n_1541),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1572),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1570),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1575),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1584),
.B(n_1515),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1544),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1576),
.A2(n_1502),
.B1(n_1510),
.B2(n_1561),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1578),
.B(n_1562),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1584),
.A2(n_1545),
.B(n_1540),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1595),
.B(n_1564),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1581),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1537),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1586),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1562),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1586),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1437),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1583),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1554),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1575),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1585),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1613),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1613),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1618),
.B(n_1575),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1617),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1617),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1601),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1607),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1616),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1607),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1610),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1609),
.B(n_1577),
.Y(n_1645)
);

NAND2x1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.B(n_1571),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1602),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_L g1648 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_R g1653 ( 
.A(n_1601),
.B(n_1452),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1601),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1611),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1596),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1623),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1596),
.B(n_1594),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1599),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1623),
.B(n_1592),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1647),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1622),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1647),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1622),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1626),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1627),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1636),
.B(n_1622),
.Y(n_1669)
);

BUFx2_ASAP7_75t_SL g1670 ( 
.A(n_1637),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1628),
.B(n_1622),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1620),
.Y(n_1672)
);

NAND2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1636),
.B(n_1588),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1627),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1599),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_SL g1679 ( 
.A(n_1653),
.B(n_1523),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1638),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1631),
.B(n_1633),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1641),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1633),
.B(n_1620),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1642),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.Y(n_1687)
);

AOI21xp33_ASAP7_75t_SL g1688 ( 
.A1(n_1637),
.A2(n_1527),
.B(n_1529),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1630),
.B(n_1615),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1654),
.B(n_1588),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1630),
.B(n_1621),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1645),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1474),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1640),
.B(n_1600),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1645),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.B(n_1600),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1656),
.B(n_1624),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1658),
.B(n_1612),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1642),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1634),
.B(n_1618),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1673),
.B(n_1692),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1673),
.B(n_1654),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1679),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1662),
.B(n_1624),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1666),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1664),
.B(n_1639),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1667),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1694),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1667),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1669),
.B(n_1514),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1700),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1449),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1669),
.B(n_1529),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1695),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1668),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1672),
.B(n_1685),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1688),
.B(n_1656),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1657),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1668),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1702),
.B(n_1678),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1678),
.B(n_1661),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1696),
.B(n_1643),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1692),
.B(n_1651),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1670),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1692),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1691),
.B(n_1625),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1694),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1657),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1698),
.B(n_1660),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1674),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1698),
.B(n_1661),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1694),
.B(n_1697),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1674),
.Y(n_1740)
);

OAI32xp33_ASAP7_75t_L g1741 ( 
.A1(n_1724),
.A2(n_1651),
.A3(n_1597),
.B1(n_1697),
.B2(n_1665),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1718),
.B(n_1697),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1733),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1724),
.A2(n_1597),
.B(n_1663),
.C(n_1665),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1733),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1707),
.A2(n_1598),
.B1(n_1604),
.B2(n_1531),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1716),
.A2(n_1671),
.B(n_1663),
.C(n_1646),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1719),
.A2(n_1598),
.B1(n_1604),
.B2(n_1590),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1671),
.C(n_1704),
.D(n_1689),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1727),
.B(n_1693),
.Y(n_1751)
);

O2A1O1Ixp33_ASAP7_75t_SL g1752 ( 
.A1(n_1730),
.A2(n_1646),
.B(n_1659),
.C(n_1512),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1721),
.B(n_1651),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1708),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1660),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1710),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1709),
.B(n_1711),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1712),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1715),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_SL g1761 ( 
.A1(n_1730),
.A2(n_1659),
.B(n_1517),
.C(n_1525),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1720),
.A2(n_1511),
.B1(n_1618),
.B2(n_1651),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1693),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1729),
.B(n_1675),
.Y(n_1764)
);

OAI32xp33_ASAP7_75t_L g1765 ( 
.A1(n_1731),
.A2(n_1704),
.A3(n_1689),
.B1(n_1675),
.B2(n_1684),
.Y(n_1765)
);

AOI32xp33_ASAP7_75t_L g1766 ( 
.A1(n_1705),
.A2(n_1573),
.A3(n_1579),
.B1(n_1699),
.B2(n_1701),
.Y(n_1766)
);

AOI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1741),
.A2(n_1740),
.B1(n_1722),
.B2(n_1726),
.C(n_1737),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1713),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1744),
.B(n_1732),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1763),
.B(n_1706),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1749),
.A2(n_1739),
.B1(n_1546),
.B2(n_1734),
.C(n_1648),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1765),
.A2(n_1735),
.B(n_1734),
.C(n_1736),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1746),
.A2(n_1590),
.B1(n_1618),
.B2(n_1573),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1762),
.A2(n_1618),
.B1(n_1714),
.B2(n_1728),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1753),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1758),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1766),
.A2(n_1648),
.B(n_1706),
.C(n_1717),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1735),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1743),
.B(n_1717),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1753),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1742),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1762),
.A2(n_1757),
.B1(n_1760),
.B2(n_1754),
.C1(n_1759),
.C2(n_1756),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1764),
.Y(n_1784)
);

OAI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1747),
.A2(n_1736),
.B(n_1725),
.C(n_1738),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1783),
.A2(n_1750),
.B1(n_1761),
.B2(n_1755),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1772),
.A2(n_1761),
.B(n_1752),
.C(n_1687),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1782),
.B(n_1699),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_SL g1790 ( 
.A(n_1785),
.B(n_1752),
.C(n_1526),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1776),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1772),
.A2(n_1687),
.B(n_1683),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1777),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1769),
.A2(n_1701),
.B(n_1539),
.Y(n_1794)
);

XNOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1775),
.B(n_1588),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1780),
.B(n_1634),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_L g1797 ( 
.A(n_1770),
.B(n_1676),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1786),
.Y(n_1798)
);

NAND2x1_ASAP7_75t_L g1799 ( 
.A(n_1790),
.B(n_1784),
.Y(n_1799)
);

NOR3xp33_ASAP7_75t_L g1800 ( 
.A(n_1798),
.B(n_1769),
.C(n_1771),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1789),
.Y(n_1801)
);

NAND2xp33_ASAP7_75t_SL g1802 ( 
.A(n_1795),
.B(n_1779),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1791),
.B(n_1768),
.Y(n_1803)
);

OAI321xp33_ASAP7_75t_L g1804 ( 
.A1(n_1787),
.A2(n_1774),
.A3(n_1767),
.B1(n_1773),
.B2(n_1778),
.C(n_1781),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1796),
.B(n_1670),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1794),
.B(n_1625),
.Y(n_1806)
);

NAND5xp2_ASAP7_75t_L g1807 ( 
.A(n_1788),
.B(n_1625),
.C(n_1645),
.D(n_1535),
.E(n_1524),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1793),
.Y(n_1808)
);

NAND2x1_ASAP7_75t_L g1809 ( 
.A(n_1792),
.B(n_1676),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1800),
.B(n_1797),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1799),
.A2(n_1703),
.B1(n_1677),
.B2(n_1680),
.Y(n_1811)
);

NOR4xp25_ASAP7_75t_L g1812 ( 
.A(n_1804),
.B(n_1683),
.C(n_1690),
.D(n_1687),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1809),
.A2(n_1804),
.B(n_1802),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1807),
.A2(n_1690),
.B1(n_1683),
.B2(n_1703),
.C(n_1684),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1812),
.A2(n_1808),
.B1(n_1801),
.B2(n_1803),
.C(n_1805),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1813),
.A2(n_1806),
.B(n_1606),
.C(n_1478),
.Y(n_1816)
);

A2O1A1Ixp33_ASAP7_75t_SL g1817 ( 
.A1(n_1810),
.A2(n_1811),
.B(n_1686),
.C(n_1681),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1677),
.Y(n_1818)
);

NOR2x1_ASAP7_75t_SL g1819 ( 
.A(n_1811),
.B(n_1478),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1813),
.A2(n_1690),
.B(n_1686),
.C(n_1681),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1818),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1815),
.B(n_1680),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1819),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1820),
.B(n_1548),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1816),
.B(n_1524),
.C(n_1619),
.Y(n_1825)
);

OAI321xp33_ASAP7_75t_L g1826 ( 
.A1(n_1823),
.A2(n_1817),
.A3(n_1587),
.B1(n_1579),
.B2(n_1589),
.C(n_1593),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1824),
.B(n_1643),
.Y(n_1827)
);

AOI32xp33_ASAP7_75t_L g1828 ( 
.A1(n_1822),
.A2(n_1652),
.A3(n_1530),
.B1(n_1534),
.B2(n_1520),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1827),
.Y(n_1829)
);

OAI22x1_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1821),
.B1(n_1825),
.B2(n_1826),
.Y(n_1830)
);

XNOR2xp5_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1828),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1830),
.A2(n_1655),
.B1(n_1644),
.B2(n_1649),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1831),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1832),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1833),
.A2(n_1834),
.B1(n_1655),
.B2(n_1644),
.Y(n_1835)
);

AOI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1530),
.B(n_1534),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1835),
.A2(n_1616),
.B(n_1619),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1837),
.B(n_1836),
.Y(n_1838)
);

OR2x6_ASAP7_75t_L g1839 ( 
.A(n_1838),
.B(n_1530),
.Y(n_1839)
);

OAI221xp5_ASAP7_75t_R g1840 ( 
.A1(n_1839),
.A2(n_1534),
.B1(n_1652),
.B2(n_1575),
.C(n_1650),
.Y(n_1840)
);

AOI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1521),
.B(n_1522),
.C(n_1516),
.Y(n_1841)
);


endmodule