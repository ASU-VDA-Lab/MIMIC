module fake_netlist_1_8100_n_6 (n_1, n_0, n_6);
input n_1;
input n_0;
output n_6;
wire n_2;
wire n_4;
wire n_3;
wire n_5;
NAND2xp5_ASAP7_75t_L g2 ( .A(n_1), .B(n_0), .Y(n_2) );
NOR2xp33_ASAP7_75t_SL g3 ( .A(n_0), .B(n_1), .Y(n_3) );
BUFx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
AOI211xp5_ASAP7_75t_SL g5 ( .A1(n_4), .A2(n_3), .B(n_0), .C(n_1), .Y(n_5) );
AOI22xp33_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_3), .B1(n_0), .B2(n_1), .Y(n_6) );
endmodule