module fake_jpeg_11676_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_15),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_49),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_41),
.B1(n_33),
.B2(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_32),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_60),
.B1(n_33),
.B2(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_20),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_29),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_17),
.B1(n_72),
.B2(n_55),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_18),
.C(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_25),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_40),
.C(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_78),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_64),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_116),
.B1(n_72),
.B2(n_87),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_64),
.A3(n_57),
.B1(n_71),
.B2(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_25),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_113),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_67),
.B(n_54),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_112),
.B(n_87),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_66),
.B(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_80),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_19),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_19),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_106),
.C(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_84),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_131),
.B(n_133),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_81),
.C(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_110),
.B1(n_102),
.B2(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_76),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_116),
.B1(n_100),
.B2(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_146),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_101),
.Y(n_147)
);

AOI22x1_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_102),
.B1(n_51),
.B2(n_98),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_149),
.B(n_121),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_95),
.B(n_91),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_56),
.B1(n_85),
.B2(n_75),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_124),
.B1(n_121),
.B2(n_119),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_148),
.B(n_139),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_120),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_149),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_67),
.B(n_54),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_152),
.A3(n_158),
.B1(n_157),
.B2(n_153),
.C1(n_151),
.C2(n_160),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_165),
.B(n_26),
.Y(n_176)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_142),
.B(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_7),
.B(n_8),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_173),
.C(n_17),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_9),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_163),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_24),
.B1(n_12),
.B2(n_13),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_176),
.B(n_26),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_162),
.C(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_134),
.C(n_75),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_56),
.B1(n_26),
.B2(n_27),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_182),
.B1(n_11),
.B2(n_19),
.Y(n_184)
);

NAND4xp25_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_172),
.C(n_13),
.D(n_11),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_184),
.B(n_27),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_188),
.B(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_27),
.B(n_63),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_185),
.Y(n_190)
);


endmodule