module fake_jpeg_26572_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_30),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_46),
.B(n_9),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_22),
.B(n_15),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_21),
.B1(n_11),
.B2(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_13),
.B1(n_17),
.B2(n_6),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_21),
.C(n_10),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_11),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_38),
.B1(n_40),
.B2(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_8),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_57),
.B(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_13),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_54),
.C(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_4),
.B(n_7),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_55),
.C(n_60),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_65),
.B(n_7),
.Y(n_74)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B(n_71),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_70),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_76),
.Y(n_77)
);


endmodule