module fake_netlist_6_4708_n_1335 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1335);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1335;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_474;
wire n_1207;
wire n_527;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_934;
wire n_482;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_814;
wire n_389;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g316 ( 
.A(n_121),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_144),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_132),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_58),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_167),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_49),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_75),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_138),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_72),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_62),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_47),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_101),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_116),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_281),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_44),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_51),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_213),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_192),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_161),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_239),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_277),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_104),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_191),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_81),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_165),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_153),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_47),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_168),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_251),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_238),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_174),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_118),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_236),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_219),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_154),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_137),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_43),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_157),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_228),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_224),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_130),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_308),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_86),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_159),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_145),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_252),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_156),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_49),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_179),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_88),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_68),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_173),
.Y(n_381)
);

BUFx2_ASAP7_75t_SL g382 ( 
.A(n_79),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_65),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_163),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_169),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_148),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_208),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_227),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_56),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_273),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_286),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_13),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_306),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_45),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_287),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_51),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_139),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_262),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_243),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_237),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_304),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_186),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_210),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_108),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_129),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_3),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_162),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_282),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_36),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_22),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_7),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_175),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_310),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_37),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_19),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_12),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_57),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_285),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_1),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_266),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_166),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_66),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_200),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_222),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_126),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_189),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_98),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_55),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_170),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_298),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_172),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_30),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_197),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_209),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_283),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_217),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_73),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_29),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_229),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_16),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_312),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_232),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_315),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_82),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_245),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_225),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_2),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_212),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_119),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_307),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_185),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_178),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_177),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_120),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_270),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_7),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_36),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_176),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_211),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_233),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_297),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_201),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_220),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_50),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_215),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_123),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_147),
.B(n_10),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_265),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_103),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_276),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_184),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_302),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_257),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_155),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_188),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_261),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_246),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_206),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_296),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_196),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_105),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_214),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_59),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_291),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_256),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_136),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_37),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_128),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_80),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_199),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_267),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_260),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_14),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_142),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_25),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_53),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_71),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_11),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_181),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_151),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_33),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_112),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_0),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_15),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_160),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_180),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_4),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_25),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_92),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_131),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_114),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_135),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_223),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_19),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_46),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_309),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_249),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_41),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_27),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_303),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_230),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_280),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_134),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_38),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_23),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_264),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_4),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_269),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_158),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_250),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_203),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_53),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_171),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_48),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_231),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_133),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_125),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_124),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_194),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_95),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_107),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_314),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_328),
.B(n_0),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_419),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_349),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_419),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_349),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_325),
.B(n_1),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_349),
.Y(n_550)
);

INVx6_ASAP7_75t_L g551 ( 
.A(n_542),
.Y(n_551)
);

CKINVDCx6p67_ASAP7_75t_R g552 ( 
.A(n_494),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_542),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_325),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_349),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_352),
.B(n_2),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_525),
.Y(n_560)
);

BUFx12f_ASAP7_75t_L g561 ( 
.A(n_473),
.Y(n_561)
);

AOI22x1_ASAP7_75t_SL g562 ( 
.A1(n_324),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_499),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_525),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_523),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_340),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_523),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_473),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_352),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_370),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_533),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_533),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_370),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_331),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_321),
.B(n_8),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_317),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_321),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_361),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_376),
.Y(n_583)
);

OAI22x1_ASAP7_75t_L g584 ( 
.A1(n_504),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_372),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_414),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_318),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_335),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_356),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_439),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_330),
.B(n_9),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_392),
.Y(n_592)
);

INVx6_ASAP7_75t_L g593 ( 
.A(n_385),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_463),
.B(n_12),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_319),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_516),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_330),
.B(n_13),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_336),
.Y(n_599)
);

BUFx12f_ASAP7_75t_L g600 ( 
.A(n_374),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_377),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_394),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_392),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_387),
.B(n_14),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_406),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_332),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_406),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_387),
.B(n_15),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_334),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_399),
.B(n_405),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_322),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_396),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_316),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_409),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_399),
.A2(n_17),
.B(n_18),
.Y(n_618)
);

BUFx8_ASAP7_75t_SL g619 ( 
.A(n_338),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_405),
.B(n_20),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_495),
.B(n_20),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_323),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_526),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_418),
.B(n_21),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_410),
.Y(n_625)
);

OAI22x1_ASAP7_75t_R g626 ( 
.A1(n_411),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_626)
);

OAI22x1_ASAP7_75t_SL g627 ( 
.A1(n_415),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_339),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_416),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_429),
.B(n_28),
.Y(n_630)
);

AOI22x1_ASAP7_75t_SL g631 ( 
.A1(n_433),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_327),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_326),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_429),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_440),
.B(n_31),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_441),
.Y(n_636)
);

BUFx8_ASAP7_75t_SL g637 ( 
.A(n_362),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_440),
.B(n_32),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_453),
.B(n_32),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_453),
.B(n_33),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_448),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_454),
.B(n_34),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_457),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_337),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_458),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_488),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_343),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_454),
.B(n_35),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_496),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_329),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_455),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_502),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_505),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_320),
.B(n_455),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_347),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_348),
.Y(n_656)
);

INVx6_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_333),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_460),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_460),
.B(n_39),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_487),
.B(n_40),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_515),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_487),
.B(n_42),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_382),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_353),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_357),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_358),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_363),
.B(n_371),
.Y(n_668)
);

BUFx8_ASAP7_75t_SL g669 ( 
.A(n_369),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_373),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_379),
.Y(n_671)
);

OAI22x1_ASAP7_75t_SL g672 ( 
.A1(n_519),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_384),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_520),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_390),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_395),
.B(n_48),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_341),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_402),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_404),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_407),
.B(n_50),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_412),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_413),
.Y(n_684)
);

OAI22x1_ASAP7_75t_SL g685 ( 
.A1(n_375),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_398),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_426),
.A2(n_52),
.B1(n_61),
.B2(n_63),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_417),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_424),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_425),
.B(n_64),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_346),
.B(n_67),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_430),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_342),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_431),
.B(n_69),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_432),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_435),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_437),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_443),
.A2(n_70),
.B(n_74),
.Y(n_698)
);

BUFx12f_ASAP7_75t_L g699 ( 
.A(n_344),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_561),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_607),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_R g703 ( 
.A(n_596),
.B(n_445),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_612),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_553),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_548),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_619),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_R g708 ( 
.A1(n_564),
.A2(n_447),
.B1(n_462),
.B2(n_450),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_637),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_654),
.B(n_367),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_669),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_686),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_693),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_699),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_649),
.B(n_652),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_580),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_614),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_632),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_R g719 ( 
.A(n_628),
.B(n_449),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_550),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_658),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_585),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_588),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_643),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_664),
.B(n_475),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_600),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_593),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_602),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_568),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_560),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_R g733 ( 
.A(n_601),
.B(n_345),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_662),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_565),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_615),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_645),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_593),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_630),
.A2(n_468),
.B(n_480),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_587),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_622),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_622),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_625),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_650),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_650),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_679),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_679),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_679),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_646),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_574),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_664),
.B(n_482),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_629),
.B(n_636),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_674),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_694),
.A2(n_484),
.B(n_483),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_664),
.B(n_486),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_570),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_575),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_581),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_552),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_657),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_657),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_581),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_589),
.B(n_492),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_634),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_571),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_551),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_577),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_R g771 ( 
.A(n_629),
.B(n_472),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_571),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_651),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_651),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_568),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_569),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_554),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_636),
.B(n_350),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_556),
.B(n_500),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_676),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_599),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_676),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_675),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_R g784 ( 
.A(n_691),
.B(n_351),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_571),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_675),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_572),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_568),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_572),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_572),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_624),
.A2(n_471),
.B1(n_490),
.B2(n_464),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_576),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_R g793 ( 
.A(n_545),
.B(n_354),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_576),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_576),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_R g796 ( 
.A(n_547),
.B(n_355),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_688),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_789),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_710),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_710),
.B(n_544),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_759),
.B(n_589),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_763),
.B(n_589),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_775),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_765),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_766),
.B(n_690),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_SL g806 ( 
.A(n_731),
.B(n_559),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_764),
.B(n_559),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_769),
.B(n_690),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_773),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_774),
.B(n_559),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_788),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_715),
.B(n_566),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_739),
.B(n_566),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_702),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_791),
.B(n_638),
.C(n_635),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_770),
.B(n_660),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_776),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_702),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_725),
.A2(n_584),
.B1(n_621),
.B2(n_653),
.C(n_627),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_785),
.B(n_549),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_739),
.B(n_566),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_780),
.B(n_594),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_757),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_SL g826 ( 
.A(n_771),
.B(n_549),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_787),
.B(n_557),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_731),
.Y(n_828)
);

BUFx6f_ASAP7_75t_SL g829 ( 
.A(n_776),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_726),
.B(n_556),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_733),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_797),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_790),
.B(n_792),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_720),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_732),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_784),
.B(n_668),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_794),
.B(n_557),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_751),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_782),
.B(n_605),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_784),
.B(n_668),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_725),
.B(n_605),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_758),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_706),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_723),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_SL g846 ( 
.A(n_753),
.B(n_661),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_740),
.B(n_659),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_730),
.Y(n_848)
);

BUFx8_ASAP7_75t_L g849 ( 
.A(n_705),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_734),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_735),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_772),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_747),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_781),
.B(n_678),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_795),
.B(n_687),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_779),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_777),
.B(n_579),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_741),
.B(n_682),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_742),
.B(n_659),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_768),
.B(n_579),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_744),
.B(n_616),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_734),
.B(n_563),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_745),
.B(n_591),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_716),
.B(n_647),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_733),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_752),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_756),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_750),
.B(n_617),
.C(n_567),
.Y(n_869)
);

BUFx5_ASAP7_75t_L g870 ( 
.A(n_746),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_796),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_778),
.B(n_659),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_717),
.B(n_655),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_778),
.B(n_613),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_718),
.A2(n_698),
.B(n_598),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_703),
.B(n_591),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_721),
.B(n_656),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_748),
.B(n_613),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_793),
.Y(n_879)
);

INVxp33_ASAP7_75t_L g880 ( 
.A(n_719),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_749),
.B(n_666),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_703),
.B(n_598),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_793),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_700),
.B(n_641),
.C(n_531),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_783),
.B(n_670),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_786),
.B(n_671),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_761),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_701),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_820),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_800),
.A2(n_507),
.B1(n_510),
.B2(n_503),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_799),
.B(n_762),
.Y(n_891)
);

BUFx8_ASAP7_75t_L g892 ( 
.A(n_829),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_825),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_888),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_858),
.B(n_604),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_843),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_814),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_831),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_834),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_818),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_854),
.B(n_604),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_867),
.B(n_611),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_866),
.B(n_743),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_835),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_798),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_839),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_863),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_836),
.B(n_713),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_846),
.A2(n_708),
.B1(n_754),
.B2(n_722),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_868),
.B(n_611),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_815),
.A2(n_620),
.B1(n_640),
.B2(n_639),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_874),
.B(n_620),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_875),
.B(n_862),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_856),
.B(n_578),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_836),
.B(n_714),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_640),
.B(n_642),
.C(n_639),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_865),
.B(n_728),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_850),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_837),
.B(n_642),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_887),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_829),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_878),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_815),
.A2(n_648),
.B1(n_663),
.B2(n_618),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_844),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_836),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_873),
.B(n_738),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_819),
.A2(n_648),
.B1(n_663),
.B2(n_618),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_859),
.A2(n_518),
.B(n_521),
.C(n_517),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_871),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_849),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_852),
.B(n_359),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_845),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_848),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_869),
.A2(n_685),
.B1(n_696),
.B2(n_681),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_803),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_811),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_813),
.A2(n_698),
.B(n_530),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_852),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_822),
.B(n_583),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_805),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_808),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_879),
.B(n_724),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_804),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_809),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_877),
.B(n_876),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_832),
.B(n_582),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_841),
.B(n_529),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_883),
.B(n_727),
.Y(n_950)
);

AND3x1_ASAP7_75t_L g951 ( 
.A(n_884),
.B(n_626),
.C(n_562),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_821),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_828),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_872),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_882),
.B(n_729),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_830),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_847),
.B(n_860),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_851),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_812),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_864),
.A2(n_538),
.B1(n_541),
.B2(n_536),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_827),
.B(n_586),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_851),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_851),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_870),
.B(n_823),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_870),
.B(n_543),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_SL g966 ( 
.A(n_816),
.B(n_760),
.C(n_707),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_851),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_842),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_851),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_826),
.A2(n_684),
.B1(n_677),
.B2(n_633),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_838),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_886),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_881),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_870),
.B(n_644),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_857),
.A2(n_824),
.B(n_861),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_810),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_833),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_885),
.A2(n_683),
.B(n_665),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_801),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_855),
.A2(n_684),
.B1(n_677),
.B2(n_697),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_802),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_817),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_830),
.A2(n_695),
.B1(n_680),
.B2(n_364),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_870),
.B(n_680),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_894),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_890),
.A2(n_695),
.B(n_597),
.C(n_590),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_958),
.A2(n_840),
.B(n_807),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_958),
.A2(n_807),
.B(n_880),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_967),
.A2(n_365),
.B(n_360),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_947),
.B(n_704),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_967),
.A2(n_368),
.B(n_366),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_917),
.A2(n_380),
.B(n_378),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_900),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_914),
.A2(n_902),
.B(n_896),
.C(n_920),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_964),
.A2(n_383),
.B(n_381),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_891),
.B(n_899),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_897),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_926),
.B(n_972),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_926),
.B(n_870),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_SL g1000 ( 
.A(n_926),
.B(n_386),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_969),
.A2(n_608),
.B(n_603),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_942),
.B(n_388),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_945),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_943),
.A2(n_673),
.B1(n_689),
.B2(n_667),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_951),
.A2(n_672),
.B1(n_595),
.B2(n_606),
.C(n_609),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_973),
.B(n_709),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_919),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_957),
.B(n_389),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_889),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_982),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_889),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_906),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_974),
.A2(n_393),
.B(n_391),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_928),
.A2(n_673),
.B1(n_689),
.B2(n_667),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_946),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_924),
.A2(n_913),
.B1(n_912),
.B2(n_954),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_912),
.A2(n_400),
.B1(n_401),
.B2(n_397),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_895),
.B(n_711),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_984),
.A2(n_408),
.B(n_403),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_889),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_903),
.B(n_420),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_975),
.A2(n_498),
.B(n_422),
.C(n_423),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_939),
.A2(n_427),
.B(n_421),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_905),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_907),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_893),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_930),
.B(n_712),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_911),
.A2(n_501),
.B1(n_434),
.B2(n_436),
.Y(n_1028)
);

AO22x1_ASAP7_75t_L g1029 ( 
.A1(n_904),
.A2(n_737),
.B1(n_736),
.B2(n_631),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_966),
.B(n_960),
.C(n_922),
.Y(n_1030)
);

OR2x6_ASAP7_75t_SL g1031 ( 
.A(n_931),
.B(n_428),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_956),
.A2(n_442),
.B(n_438),
.Y(n_1032)
);

OAI22x1_ASAP7_75t_L g1033 ( 
.A1(n_935),
.A2(n_493),
.B1(n_446),
.B2(n_451),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_933),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_936),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_949),
.B(n_444),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_959),
.B(n_452),
.Y(n_1038)
);

BUFx10_ASAP7_75t_L g1039 ( 
.A(n_918),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_965),
.A2(n_459),
.B(n_456),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_927),
.B(n_461),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_940),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_466),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_941),
.B(n_467),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_898),
.A2(n_592),
.B(n_610),
.C(n_623),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_961),
.A2(n_513),
.B(n_470),
.C(n_474),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_979),
.A2(n_522),
.B1(n_476),
.B2(n_477),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_893),
.B(n_469),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_935),
.A2(n_512),
.B1(n_479),
.B2(n_481),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_962),
.A2(n_485),
.B(n_478),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_976),
.B(n_489),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_981),
.B(n_491),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_901),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_948),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_963),
.A2(n_953),
.B(n_934),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_915),
.B(n_506),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_983),
.A2(n_540),
.B(n_514),
.C(n_524),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_925),
.A2(n_968),
.B(n_932),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_994),
.A2(n_952),
.B(n_983),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_985),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_997),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1003),
.Y(n_1062)
);

BUFx2_ASAP7_75t_R g1063 ( 
.A(n_1031),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_1009),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_993),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1041),
.A2(n_971),
.B1(n_977),
.B2(n_921),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_996),
.B(n_948),
.Y(n_1067)
);

BUFx4f_ASAP7_75t_SL g1068 ( 
.A(n_1010),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1001),
.A2(n_1055),
.B(n_987),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1015),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1053),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1007),
.B(n_910),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_1011),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_1027),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_1011),
.B(n_977),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_SL g1076 ( 
.A1(n_1058),
.A2(n_978),
.B(n_970),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1024),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1025),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1034),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_1012),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1039),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1020),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_999),
.A2(n_938),
.B(n_937),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1016),
.A2(n_950),
.B(n_938),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_1023),
.A2(n_929),
.B(n_955),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_1020),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1020),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_1022),
.A2(n_916),
.B(n_909),
.Y(n_1089)
);

INVx3_ASAP7_75t_SL g1090 ( 
.A(n_1026),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1008),
.B(n_977),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_1050),
.A2(n_944),
.B(n_937),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_1026),
.B(n_971),
.Y(n_1093)
);

CKINVDCx16_ASAP7_75t_R g1094 ( 
.A(n_1018),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1030),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1014),
.A2(n_980),
.B(n_527),
.Y(n_1096)
);

INVx6_ASAP7_75t_SL g1097 ( 
.A(n_1054),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_990),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_1036),
.B(n_892),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_998),
.Y(n_1100)
);

BUFx2_ASAP7_75t_SL g1101 ( 
.A(n_1042),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_1006),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_1043),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1044),
.B(n_592),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1000),
.B(n_806),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1021),
.A2(n_673),
.B(n_667),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1045),
.Y(n_1107)
);

BUFx2_ASAP7_75t_R g1108 ( 
.A(n_1056),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_689),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_988),
.A2(n_623),
.B(n_76),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_SL g1111 ( 
.A(n_1029),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1038),
.B(n_692),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_992),
.A2(n_692),
.B(n_532),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1051),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_986),
.Y(n_1115)
);

INVx6_ASAP7_75t_L g1116 ( 
.A(n_1033),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1098),
.A2(n_1017),
.B1(n_1052),
.B2(n_1037),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1060),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1060),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1061),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1061),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1062),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1114),
.A2(n_1057),
.B(n_1046),
.C(n_1005),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1068),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1065),
.B(n_1077),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1103),
.B(n_1047),
.Y(n_1126)
);

INVx6_ASAP7_75t_L g1127 ( 
.A(n_1087),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1070),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1059),
.A2(n_995),
.B(n_1013),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1070),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1071),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1071),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1115),
.A2(n_1049),
.B1(n_692),
.B2(n_1004),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1102),
.A2(n_1028),
.B1(n_1048),
.B2(n_511),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1090),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1094),
.A2(n_1032),
.B1(n_989),
.B2(n_991),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1067),
.B(n_534),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1072),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1115),
.A2(n_539),
.B1(n_537),
.B2(n_1019),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1116),
.A2(n_1040),
.B1(n_78),
.B2(n_83),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1080),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1078),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1081),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1066),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1078),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1079),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1079),
.Y(n_1147)
);

BUFx4f_ASAP7_75t_SL g1148 ( 
.A(n_1097),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1091),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1074),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1116),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1082),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1107),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_1153)
);

INVx6_ASAP7_75t_L g1154 ( 
.A(n_1064),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1085),
.A2(n_100),
.B(n_102),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_1064),
.B(n_106),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1107),
.A2(n_1109),
.B(n_1110),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1084),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1069),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1097),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1076),
.A2(n_109),
.B(n_110),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1106),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1138),
.B(n_1095),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1126),
.A2(n_1101),
.B1(n_1108),
.B2(n_1100),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_1104),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1118),
.Y(n_1166)
);

AND2x2_ASAP7_75t_SL g1167 ( 
.A(n_1151),
.B(n_1153),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1150),
.B(n_1063),
.C(n_1111),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1119),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1117),
.A2(n_1112),
.B(n_1089),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1143),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1120),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1120),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1161),
.A2(n_1092),
.B(n_1096),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1125),
.B(n_1075),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1123),
.B(n_1093),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1141),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1135),
.B(n_1073),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1135),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_1124),
.B(n_1099),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1148),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_1144),
.A2(n_1089),
.B(n_1096),
.C(n_1086),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1122),
.B(n_1083),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1128),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1139),
.A2(n_1105),
.B(n_1086),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1130),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_R g1188 ( 
.A(n_1160),
.B(n_111),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1127),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1130),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1154),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1159),
.A2(n_1158),
.B(n_1162),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1132),
.B(n_1083),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1146),
.B(n_1088),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1149),
.A2(n_1113),
.B1(n_1088),
.B2(n_115),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1142),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1127),
.B(n_1156),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1146),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1140),
.B(n_113),
.C(n_117),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1179),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1192),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1167),
.B(n_1147),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1166),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1175),
.B(n_1197),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1166),
.B(n_1131),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1172),
.B(n_1145),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1173),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1165),
.B(n_1152),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1199),
.A2(n_1133),
.B1(n_1153),
.B2(n_1151),
.C(n_1136),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1193),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1193),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1180),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1185),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1187),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1171),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1187),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1169),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1194),
.B(n_1163),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1190),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1190),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1196),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1184),
.B(n_1134),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1198),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1176),
.B(n_1155),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1177),
.B(n_1155),
.Y(n_1225)
);

AOI222xp33_ASAP7_75t_L g1226 ( 
.A1(n_1164),
.A2(n_1158),
.B1(n_1159),
.B2(n_140),
.C1(n_141),
.C2(n_143),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1174),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1186),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1170),
.B(n_1157),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1191),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1178),
.B(n_1129),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1191),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1189),
.B(n_127),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1218),
.B(n_1181),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1231),
.B(n_1168),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1203),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1203),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1213),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1225),
.B(n_1182),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1226),
.B(n_1188),
.C(n_1195),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1213),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1207),
.Y(n_1242)
);

OAI21xp33_ASAP7_75t_L g1243 ( 
.A1(n_1226),
.A2(n_1209),
.B(n_1202),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1209),
.B(n_1183),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1228),
.B(n_146),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1214),
.B(n_149),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1216),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1219),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1220),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1208),
.B(n_152),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1200),
.B(n_164),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1201),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1212),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1212),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1204),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1204),
.B(n_1222),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1223),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1227),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1239),
.B(n_1229),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1242),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1257),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1257),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1239),
.B(n_1224),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1253),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1248),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1249),
.B(n_1221),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1247),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1246),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1256),
.B(n_1210),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1236),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1237),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1238),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1241),
.B(n_1211),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1254),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1252),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1258),
.B(n_1230),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1255),
.B(n_1232),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1259),
.A2(n_1243),
.B(n_1240),
.C(n_1244),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1260),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1275),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1263),
.B(n_1234),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1264),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1263),
.B(n_1235),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1267),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_1269),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1279),
.Y(n_1286)
);

OAI21xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1283),
.A2(n_1268),
.B(n_1270),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1278),
.A2(n_1246),
.B(n_1245),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1285),
.B(n_1277),
.Y(n_1289)
);

OAI221xp5_ASAP7_75t_L g1290 ( 
.A1(n_1282),
.A2(n_1272),
.B1(n_1271),
.B2(n_1251),
.C(n_1274),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1284),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1286),
.B(n_1280),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1289),
.B(n_1281),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1290),
.B(n_1215),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1288),
.A2(n_1287),
.B(n_1291),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1294),
.B(n_1273),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1293),
.B(n_1261),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1295),
.A2(n_1276),
.B(n_1262),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1292),
.B(n_1262),
.Y(n_1299)
);

NAND2x1_ASAP7_75t_L g1300 ( 
.A(n_1299),
.B(n_1265),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1298),
.A2(n_1233),
.B(n_1250),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1301),
.B(n_1266),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1302),
.A2(n_1205),
.B(n_1206),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1300),
.B(n_1217),
.Y(n_1305)
);

NOR4xp25_ASAP7_75t_L g1306 ( 
.A(n_1303),
.B(n_182),
.C(n_183),
.D(n_190),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_L g1307 ( 
.A(n_1305),
.B(n_193),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1304),
.Y(n_1308)
);

NOR3xp33_ASAP7_75t_L g1309 ( 
.A(n_1308),
.B(n_195),
.C(n_198),
.Y(n_1309)
);

NOR2x1_ASAP7_75t_L g1310 ( 
.A(n_1307),
.B(n_202),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1306),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1310),
.Y(n_1312)
);

NAND4xp25_ASAP7_75t_SL g1313 ( 
.A(n_1311),
.B(n_204),
.C(n_205),
.D(n_207),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1309),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1310),
.Y(n_1315)
);

NAND2x1_ASAP7_75t_SL g1316 ( 
.A(n_1315),
.B(n_311),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1314),
.A2(n_216),
.B1(n_221),
.B2(n_226),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1313),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1312),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1316),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1319),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1318),
.A2(n_234),
.B1(n_235),
.B2(n_240),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1317),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1318),
.A2(n_247),
.B1(n_248),
.B2(n_253),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1320),
.A2(n_254),
.B1(n_258),
.B2(n_259),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1321),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1324),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1327),
.A2(n_1323),
.B1(n_1322),
.B2(n_263),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1326),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1329),
.A2(n_1325),
.B(n_271),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1328),
.A2(n_268),
.B(n_272),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1331),
.A2(n_275),
.B1(n_284),
.B2(n_290),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1330),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1333),
.B(n_299),
.Y(n_1334)
);

AOI211xp5_ASAP7_75t_L g1335 ( 
.A1(n_1334),
.A2(n_1332),
.B(n_300),
.C(n_301),
.Y(n_1335)
);


endmodule