module fake_jpeg_8277_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_10),
.Y(n_18)
);

OR2x2_ASAP7_75t_SL g19 ( 
.A(n_6),
.B(n_12),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_6),
.B1(n_12),
.B2(n_7),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

A2O1A1O1Ixp25_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B(n_17),
.C(n_19),
.D(n_15),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_20),
.C(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_14),
.B1(n_16),
.B2(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_32),
.B(n_36),
.Y(n_39)
);


endmodule