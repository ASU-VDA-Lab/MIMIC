module fake_netlist_6_1696_n_1846 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1846);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1846;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_6),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_78),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_14),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_88),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_23),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_67),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_143),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_118),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_70),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_35),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_96),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_126),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_82),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_42),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_13),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_23),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_83),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_155),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_128),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_110),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_39),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_73),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_14),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_93),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_81),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_121),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_98),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_46),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_35),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_37),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_120),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_115),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_47),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_75),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_154),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_38),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_13),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_142),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_107),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_160),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_111),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_127),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_40),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_91),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_79),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_77),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_194),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_36),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_17),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_196),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_173),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_90),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_141),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_85),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_125),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_46),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_11),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_161),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_102),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_119),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_116),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_189),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_8),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_89),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_187),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_198),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_117),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_135),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_137),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_53),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_104),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_183),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_80),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_157),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_29),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_151),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_129),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_10),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_61),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_192),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_59),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_51),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_114),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_108),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_181),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_162),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_65),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_8),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_138),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_32),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_30),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_24),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_174),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_184),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_65),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_71),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_163),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_16),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_16),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_4),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_133),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_167),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_32),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_68),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_57),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_53),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_109),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_105),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_2),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_166),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_169),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_124),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_29),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_10),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_64),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_50),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_55),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_131),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_19),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_63),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_48),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_7),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_175),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_43),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_132),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_177),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_76),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_191),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_11),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_130),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_49),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_24),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_176),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_202),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_147),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_26),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_51),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_182),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_56),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_37),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_139),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_15),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_172),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_149),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_145),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_48),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_61),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_180),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_199),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_36),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_50),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_92),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_9),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_43),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_63),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_6),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_274),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_291),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_239),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_306),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_284),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_284),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_1),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_400),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_239),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_241),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_328),
.B(n_1),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_249),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_229),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_269),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_239),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_239),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_251),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_264),
.B(n_2),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_239),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_242),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_252),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_308),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_223),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_254),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_242),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_229),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_242),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_335),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_256),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_257),
.B(n_3),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_242),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_298),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_352),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_270),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_242),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_273),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_210),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_337),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_206),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_337),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_282),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_210),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_283),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_257),
.B(n_3),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_337),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_290),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_292),
.B(n_4),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_337),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_353),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_337),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_354),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_212),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_216),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_352),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_294),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_354),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_296),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_299),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_233),
.B(n_5),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_317),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_354),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_214),
.B(n_9),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_392),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_333),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_250),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_354),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_399),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_338),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_364),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_364),
.Y(n_477)
);

BUFx2_ASAP7_75t_SL g478 ( 
.A(n_226),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_342),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_343),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_345),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_348),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_350),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_364),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_364),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_261),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_358),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_366),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_212),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_221),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_278),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_243),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_214),
.B(n_12),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_214),
.B(n_12),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_209),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_245),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_293),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_301),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_217),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_217),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_406),
.B(n_226),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_431),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_469),
.B(n_203),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_411),
.B(n_228),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_203),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_236),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_433),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_406),
.B(n_236),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_205),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_331),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_456),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_451),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_331),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_473),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_461),
.B(n_380),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_417),
.B(n_228),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_436),
.B(n_228),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_415),
.B(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_429),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_263),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_437),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_205),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_441),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_478),
.B(n_208),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_404),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_463),
.B(n_208),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_468),
.B(n_211),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_476),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_477),
.A2(n_330),
.B(n_312),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_485),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_419),
.B(n_211),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_501),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_487),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_498),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_419),
.B(n_218),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_443),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_466),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_408),
.B(n_218),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_410),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_412),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_413),
.B(n_380),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_414),
.B(n_204),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_466),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_453),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_445),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_492),
.B(n_219),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_428),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_424),
.B(n_213),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_405),
.B(n_228),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_460),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_416),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_420),
.B(n_312),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_518),
.B(n_448),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_416),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_522),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_567),
.B(n_418),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_573),
.B(n_228),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_567),
.B(n_573),
.Y(n_589)
);

BUFx4f_ASAP7_75t_L g590 ( 
.A(n_573),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_418),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_538),
.B(n_423),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_423),
.Y(n_593)
);

INVxp33_ASAP7_75t_SL g594 ( 
.A(n_535),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_507),
.A2(n_231),
.B1(n_295),
.B2(n_207),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_430),
.C(n_427),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_563),
.B(n_434),
.C(n_407),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_547),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_538),
.B(n_427),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_580),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_518),
.B(n_459),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_550),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_573),
.A2(n_362),
.B1(n_367),
.B2(n_330),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_552),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_567),
.B(n_430),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_567),
.B(n_573),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_362),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_563),
.B(n_435),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_573),
.A2(n_378),
.B1(n_385),
.B2(n_367),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_552),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_559),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_522),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_573),
.B(n_287),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_567),
.B(n_435),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_543),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_573),
.B(n_287),
.Y(n_627)
);

NOR2x1p5_ASAP7_75t_L g628 ( 
.A(n_581),
.B(n_490),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_531),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_502),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_560),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_531),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_546),
.B(n_378),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_579),
.A2(n_497),
.B1(n_493),
.B2(n_482),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_523),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_440),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_510),
.B(n_334),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_551),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_581),
.B(n_385),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_578),
.B(n_287),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_578),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

INVxp33_ASAP7_75t_SL g645 ( 
.A(n_535),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_564),
.B(n_440),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_581),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_522),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_523),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_581),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_576),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_564),
.A2(n_305),
.B1(n_365),
.B2(n_360),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_532),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_536),
.Y(n_655)
);

INVxp33_ASAP7_75t_L g656 ( 
.A(n_535),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_578),
.B(n_287),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_556),
.B(n_562),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_536),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_522),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_579),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_564),
.A2(n_351),
.B1(n_323),
.B2(n_346),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_574),
.B(n_442),
.Y(n_666)
);

AND3x2_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_377),
.C(n_220),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_578),
.B(n_287),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_576),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_577),
.A2(n_442),
.B1(n_489),
.B2(n_488),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_564),
.A2(n_329),
.B1(n_397),
.B2(n_383),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_510),
.B(n_447),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_522),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_532),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_536),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_537),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_532),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_516),
.B(n_447),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_516),
.B(n_449),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_509),
.B(n_449),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_531),
.Y(n_686)
);

INVx6_ASAP7_75t_L g687 ( 
.A(n_571),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_577),
.A2(n_401),
.B1(n_394),
.B2(n_224),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_534),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_533),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_571),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_542),
.B(n_452),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_562),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_542),
.B(n_452),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_533),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_517),
.B(n_462),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_539),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_539),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_572),
.A2(n_491),
.B1(n_489),
.B2(n_488),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_575),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_541),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_574),
.B(n_320),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_521),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_541),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_572),
.A2(n_491),
.B1(n_484),
.B2(n_483),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_509),
.B(n_462),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_537),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_545),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_517),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_531),
.A2(n_332),
.B1(n_324),
.B2(n_321),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_517),
.B(n_464),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_537),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_545),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_540),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_524),
.B(n_464),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_540),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_530),
.A2(n_244),
.B1(n_247),
.B2(n_260),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_534),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_565),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_524),
.B(n_465),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_530),
.B(n_467),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_604),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_621),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_652),
.B(n_467),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_683),
.B(n_524),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_641),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_659),
.B(n_529),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_669),
.B(n_471),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_693),
.B(n_529),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_682),
.B(n_471),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_637),
.B(n_475),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_664),
.A2(n_529),
.B1(n_222),
.B2(n_232),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_724),
.A2(n_571),
.B(n_565),
.C(n_549),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_585),
.B(n_531),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_653),
.A2(n_549),
.B1(n_548),
.B2(n_574),
.C(n_575),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_590),
.A2(n_474),
.B1(n_470),
.B2(n_455),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_587),
.B(n_531),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_617),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_590),
.B(n_571),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_651),
.B(n_571),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_591),
.B(n_531),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_651),
.B(n_593),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_613),
.B(n_548),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_589),
.A2(n_551),
.B(n_570),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_625),
.B(n_504),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_711),
.A2(n_570),
.B(n_566),
.C(n_569),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_631),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_712),
.B(n_551),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_666),
.B(n_475),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_700),
.B(n_480),
.C(n_479),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_643),
.B(n_209),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_646),
.B(n_479),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_692),
.B(n_480),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_592),
.B(n_504),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_695),
.B(n_483),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_615),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_724),
.A2(n_600),
.B1(n_592),
.B2(n_722),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_647),
.B(n_504),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_607),
.A2(n_551),
.B1(n_570),
.B2(n_582),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_643),
.B(n_209),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_701),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_614),
.B(n_694),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_607),
.A2(n_582),
.B1(n_504),
.B2(n_511),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_618),
.A2(n_582),
.B1(n_504),
.B2(n_511),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_643),
.B(n_209),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_694),
.B(n_511),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_694),
.B(n_511),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_633),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_697),
.B(n_307),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_209),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_705),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_618),
.A2(n_653),
.B1(n_671),
.B2(n_665),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_644),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_687),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_660),
.B(n_511),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_644),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_661),
.B(n_514),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_684),
.A2(n_569),
.B(n_568),
.C(n_566),
.Y(n_782)
);

INVx4_ASAP7_75t_SL g783 ( 
.A(n_687),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_680),
.B(n_514),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_713),
.B(n_514),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_665),
.A2(n_514),
.B1(n_393),
.B2(n_361),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_658),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_654),
.B(n_674),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_654),
.B(n_514),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_610),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_687),
.A2(n_267),
.B1(n_315),
.B2(n_395),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_701),
.B(n_674),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_672),
.B(n_219),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_685),
.B(n_503),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_685),
.B(n_209),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_639),
.B(n_503),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_620),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_667),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_606),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_639),
.B(n_505),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_619),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_672),
.B(n_225),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_609),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_715),
.B(n_505),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_681),
.B(n_225),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_715),
.B(n_506),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_690),
.B(n_506),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_696),
.B(n_508),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_671),
.A2(n_720),
.B1(n_712),
.B2(n_588),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_722),
.A2(n_285),
.B1(n_271),
.B2(n_268),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_698),
.B(n_508),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_596),
.B(n_227),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_699),
.B(n_512),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_638),
.A2(n_286),
.B1(n_262),
.B2(n_259),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_620),
.Y(n_815)
);

AO221x1_ASAP7_75t_L g816 ( 
.A1(n_720),
.A2(n_595),
.B1(n_688),
.B2(n_624),
.C(n_626),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_702),
.B(n_706),
.Y(n_817)
);

INVx8_ASAP7_75t_L g818 ( 
.A(n_641),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_689),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_710),
.B(n_512),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_720),
.A2(n_359),
.B1(n_384),
.B2(n_209),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_716),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_628),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_608),
.B(n_209),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_609),
.B(n_681),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_630),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_642),
.B(n_513),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_630),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_642),
.B(n_513),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_718),
.B(n_566),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_718),
.B(n_227),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_657),
.B(n_515),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_608),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_723),
.B(n_566),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_723),
.B(n_234),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_684),
.B(n_234),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_615),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_670),
.B(n_237),
.C(n_235),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_636),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_601),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_636),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_584),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_657),
.B(n_515),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_689),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_608),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_588),
.A2(n_384),
.B1(n_336),
.B2(n_391),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_602),
.B(n_384),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_703),
.B(n_568),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_668),
.B(n_520),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_608),
.B(n_384),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_615),
.B(n_568),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_640),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_668),
.B(n_520),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_634),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_708),
.B(n_235),
.Y(n_855)
);

BUFx6f_ASAP7_75t_SL g856 ( 
.A(n_583),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_708),
.B(n_237),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_601),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_707),
.B(n_568),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_584),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_641),
.B(n_525),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_602),
.B(n_384),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_634),
.A2(n_316),
.B1(n_313),
.B2(n_310),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_602),
.B(n_384),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_635),
.B(n_638),
.C(n_598),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_623),
.B(n_525),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_623),
.B(n_554),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_627),
.B(n_554),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_703),
.B(n_569),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_627),
.B(n_554),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_586),
.B(n_554),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_634),
.B(n_238),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_703),
.A2(n_384),
.B1(n_355),
.B2(n_277),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_586),
.B(n_554),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_586),
.B(n_569),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_602),
.B(n_384),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_622),
.B(n_528),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_649),
.A2(n_558),
.B(n_555),
.C(n_553),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_622),
.B(n_528),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_597),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_691),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_691),
.A2(n_275),
.B1(n_246),
.B2(n_248),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_770),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_771),
.A2(n_675),
.B(n_629),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_765),
.A2(n_622),
.B(n_649),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_748),
.A2(n_745),
.B(n_742),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_746),
.B(n_691),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_773),
.B(n_644),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_856),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_773),
.B(n_644),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_747),
.A2(n_675),
.B(n_662),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_754),
.A2(n_599),
.B(n_597),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_745),
.A2(n_675),
.B(n_629),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_793),
.A2(n_215),
.B(n_265),
.C(n_281),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_790),
.Y(n_895)
);

NOR2x1p5_ASAP7_75t_SL g896 ( 
.A(n_839),
.B(n_655),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_742),
.A2(n_629),
.B(n_612),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_830),
.B(n_648),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_793),
.A2(n_376),
.B(n_656),
.C(n_611),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_834),
.B(n_648),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_801),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_728),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_752),
.B(n_583),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_743),
.A2(n_629),
.B(n_612),
.Y(n_904)
);

O2A1O1Ixp5_ASAP7_75t_L g905 ( 
.A1(n_754),
.A2(n_599),
.B(n_611),
.C(n_605),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_743),
.A2(n_632),
.B(n_612),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_730),
.B(n_648),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_789),
.A2(n_788),
.B(n_796),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_785),
.B(n_648),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_726),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_800),
.A2(n_632),
.B(n_612),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_760),
.B(n_632),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_757),
.B(n_663),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_L g914 ( 
.A1(n_831),
.A2(n_224),
.B(n_221),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_732),
.B(n_663),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_776),
.A2(n_603),
.B1(n_583),
.B2(n_632),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_802),
.A2(n_656),
.B(n_616),
.C(n_605),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_802),
.A2(n_616),
.B(n_719),
.C(n_717),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_736),
.A2(n_662),
.B(n_655),
.Y(n_919)
);

INVx3_ASAP7_75t_SL g920 ( 
.A(n_819),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_603),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_734),
.B(n_663),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_778),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_778),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_797),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_727),
.B(n_603),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_741),
.B(n_594),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_877),
.A2(n_879),
.B(n_874),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_L g929 ( 
.A(n_865),
.B(n_371),
.C(n_240),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_815),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_804),
.A2(n_650),
.B(n_686),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_750),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_734),
.B(n_663),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_806),
.A2(n_650),
.B(n_686),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_755),
.B(n_673),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_763),
.A2(n_677),
.B(n_719),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_803),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_826),
.Y(n_938)
);

AO21x1_ASAP7_75t_L g939 ( 
.A1(n_836),
.A2(n_717),
.B(n_714),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_776),
.B(n_650),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_755),
.B(n_673),
.Y(n_941)
);

AND2x6_ASAP7_75t_L g942 ( 
.A(n_737),
.B(n_673),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_740),
.A2(n_650),
.B(n_686),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_844),
.B(n_594),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_809),
.A2(n_686),
.B1(n_676),
.B2(n_673),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_733),
.B(n_676),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_825),
.B(n_676),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_744),
.A2(n_761),
.B(n_777),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_828),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_733),
.B(n_676),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_777),
.A2(n_679),
.B(n_714),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_762),
.B(n_677),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_777),
.A2(n_709),
.B(n_704),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_777),
.A2(n_780),
.B(n_779),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_762),
.B(n_678),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_756),
.B(n_678),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_780),
.A2(n_679),
.B(n_709),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_756),
.B(n_704),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_780),
.A2(n_527),
.B(n_521),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_841),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_780),
.A2(n_527),
.B(n_521),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_792),
.B(n_766),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_SL g963 ( 
.A(n_805),
.B(n_721),
.C(n_403),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_772),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_731),
.B(n_240),
.C(n_238),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_758),
.B(n_553),
.Y(n_966)
);

AOI33xp33_ASAP7_75t_L g967 ( 
.A1(n_786),
.A2(n_555),
.A3(n_558),
.B1(n_230),
.B2(n_398),
.B3(n_403),
.Y(n_967)
);

CKINVDCx10_ASAP7_75t_R g968 ( 
.A(n_856),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_758),
.B(n_528),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_731),
.B(n_721),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_792),
.B(n_369),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_781),
.A2(n_527),
.B(n_526),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_831),
.B(n_368),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_784),
.A2(n_526),
.B(n_519),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_725),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_809),
.A2(n_369),
.B1(n_396),
.B2(n_390),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_774),
.A2(n_526),
.B(n_519),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_835),
.B(n_764),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_763),
.A2(n_519),
.B(n_540),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_805),
.A2(n_371),
.B1(n_396),
.B2(n_390),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_803),
.B(n_783),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_787),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_766),
.B(n_372),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_822),
.B(n_528),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_848),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_799),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_833),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_833),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_817),
.B(n_528),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_848),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_810),
.B(n_368),
.C(n_402),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_738),
.A2(n_540),
.B(n_557),
.C(n_519),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_835),
.B(n_557),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_836),
.B(n_372),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_855),
.A2(n_557),
.B(n_18),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_855),
.A2(n_645),
.B1(n_253),
.B2(n_255),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_751),
.A2(n_327),
.B(n_266),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_769),
.A2(n_544),
.B(n_339),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_857),
.B(n_258),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_769),
.A2(n_544),
.B(n_340),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_739),
.B(n_373),
.C(n_374),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_857),
.B(n_373),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_794),
.A2(n_544),
.B(n_326),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_767),
.B(n_272),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_881),
.A2(n_544),
.B(n_341),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_767),
.B(n_374),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_859),
.A2(n_881),
.B1(n_751),
.B2(n_821),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_871),
.A2(n_544),
.B(n_325),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_795),
.A2(n_544),
.B(n_347),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_759),
.B(n_645),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_837),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_852),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_795),
.A2(n_311),
.B(n_279),
.C(n_280),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_749),
.A2(n_379),
.B(n_381),
.C(n_387),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_872),
.A2(n_370),
.B(n_402),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_816),
.A2(n_370),
.B1(n_398),
.B2(n_375),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_875),
.A2(n_544),
.B(n_322),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_851),
.B(n_869),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_833),
.A2(n_544),
.B(n_319),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_869),
.B(n_379),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_842),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_867),
.A2(n_318),
.B(n_288),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_838),
.B(n_389),
.C(n_387),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_833),
.A2(n_314),
.B(n_289),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_783),
.B(n_389),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_807),
.B(n_349),
.Y(n_1026)
);

OAI321xp33_ASAP7_75t_L g1027 ( 
.A1(n_814),
.A2(n_388),
.A3(n_386),
.B1(n_382),
.B2(n_375),
.C(n_25),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_827),
.A2(n_309),
.B(n_297),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_861),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_798),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_872),
.A2(n_782),
.B(n_813),
.C(n_820),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_808),
.B(n_357),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_811),
.B(n_304),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_729),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_829),
.A2(n_363),
.B(n_300),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_832),
.A2(n_843),
.B(n_849),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_735),
.B(n_860),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_854),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_783),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_853),
.A2(n_303),
.B(n_302),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_868),
.A2(n_276),
.B(n_381),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_735),
.B(n_386),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_845),
.A2(n_382),
.B(n_74),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_870),
.A2(n_200),
.B(n_186),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_735),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_880),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_845),
.A2(n_185),
.B(n_179),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_178),
.B(n_168),
.Y(n_1048)
);

OAI321xp33_ASAP7_75t_L g1049 ( 
.A1(n_863),
.A2(n_17),
.A3(n_19),
.B1(n_20),
.B2(n_22),
.C(n_25),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_768),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_882),
.B(n_164),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_823),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_753),
.B(n_812),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_840),
.B(n_858),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_846),
.A2(n_156),
.B(n_150),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_729),
.B(n_20),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_775),
.A2(n_122),
.B(n_113),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_847),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_847),
.A2(n_103),
.B(n_101),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_873),
.A2(n_100),
.B1(n_99),
.B2(n_97),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_873),
.B(n_87),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_862),
.A2(n_86),
.B(n_84),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_878),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_929),
.B(n_791),
.C(n_824),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_902),
.B(n_818),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_927),
.A2(n_818),
.B1(n_850),
.B2(n_862),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_978),
.B(n_818),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1034),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_910),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_889),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_978),
.B(n_846),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_981),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_909),
.A2(n_876),
.B(n_864),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_913),
.A2(n_876),
.B(n_864),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_902),
.B(n_22),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_887),
.A2(n_26),
.B(n_27),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_981),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_1034),
.B(n_28),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_920),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_883),
.B(n_28),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_947),
.A2(n_31),
.B(n_34),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_883),
.A2(n_31),
.B(n_41),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_908),
.A2(n_886),
.B(n_891),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_960),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_986),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_952),
.A2(n_66),
.B(n_45),
.Y(n_1086)
);

OAI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_944),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1007),
.A2(n_52),
.B(n_54),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_932),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_923),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_1058),
.B(n_55),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_952),
.A2(n_56),
.B(n_57),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_966),
.B(n_58),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_994),
.A2(n_58),
.B(n_60),
.C(n_62),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_973),
.B(n_66),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_920),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_923),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_923),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_963),
.B(n_991),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1002),
.A2(n_1027),
.B(n_917),
.C(n_899),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_921),
.B(n_926),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1016),
.A2(n_962),
.B1(n_1045),
.B2(n_1055),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1012),
.Y(n_1103)
);

BUFx8_ASAP7_75t_L g1104 ( 
.A(n_903),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_1038),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_964),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_955),
.A2(n_900),
.B(n_898),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_975),
.B(n_1029),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_975),
.B(n_970),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_922),
.A2(n_935),
.B(n_933),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_941),
.A2(n_890),
.B(n_888),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1030),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_996),
.B(n_1010),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1053),
.A2(n_929),
.B1(n_1001),
.B2(n_1018),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1016),
.A2(n_962),
.B1(n_1045),
.B2(n_1061),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_956),
.B(n_958),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_982),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1010),
.B(n_914),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_895),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1001),
.A2(n_965),
.B(n_1023),
.C(n_919),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_901),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_965),
.B(n_1031),
.C(n_894),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1021),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_971),
.A2(n_980),
.B(n_916),
.C(n_976),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_939),
.A2(n_946),
.B(n_950),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_997),
.A2(n_971),
.B(n_1044),
.C(n_1036),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_940),
.A2(n_907),
.B(n_884),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_940),
.A2(n_885),
.B(n_948),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_985),
.B(n_990),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1034),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1034),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_993),
.B(n_1026),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_915),
.A2(n_945),
.B(n_893),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1011),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_968),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_937),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_1020),
.B1(n_937),
.B2(n_1004),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1061),
.A2(n_983),
.B1(n_1006),
.B2(n_1037),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_911),
.A2(n_931),
.B(n_934),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_SL g1141 ( 
.A1(n_1051),
.A2(n_1014),
.B(n_912),
.C(n_969),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_1020),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1038),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1063),
.A2(n_1041),
.B(n_1043),
.C(n_1056),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_989),
.B(n_1046),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_967),
.A2(n_1015),
.B(n_1006),
.C(n_983),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_925),
.B(n_938),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1054),
.A2(n_1052),
.B(n_1022),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_943),
.A2(n_947),
.B(n_897),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_930),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_937),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_923),
.B(n_924),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1025),
.A2(n_937),
.B1(n_924),
.B2(n_1050),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_949),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_924),
.B(n_987),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_987),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1025),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_984),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_924),
.B(n_995),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_904),
.A2(n_906),
.B(n_954),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_918),
.A2(n_1005),
.B(n_928),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_988),
.B(n_942),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_905),
.A2(n_977),
.B(n_972),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1003),
.A2(n_951),
.B(n_957),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1028),
.A2(n_1040),
.B1(n_1035),
.B2(n_1039),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1049),
.A2(n_1060),
.B(n_1013),
.C(n_992),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_953),
.A2(n_1008),
.B(n_998),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1000),
.A2(n_1017),
.B(n_974),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1024),
.B(n_892),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_936),
.B(n_1057),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_979),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_SL g1172 ( 
.A(n_1048),
.B(n_1062),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1009),
.A2(n_1047),
.B(n_1059),
.C(n_1019),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_959),
.B(n_961),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_896),
.B(n_942),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_942),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_942),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_942),
.A2(n_776),
.B1(n_760),
.B2(n_809),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_902),
.B(n_883),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_994),
.A2(n_1002),
.B(n_741),
.C(n_802),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_994),
.A2(n_1002),
.B(n_741),
.C(n_802),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_909),
.A2(n_590),
.B(n_765),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_994),
.A2(n_1002),
.B(n_741),
.C(n_802),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_902),
.B(n_883),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_902),
.B(n_760),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_909),
.A2(n_590),
.B(n_765),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_902),
.B(n_760),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_909),
.A2(n_590),
.B(n_765),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_978),
.A2(n_760),
.B(n_802),
.C(n_793),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_929),
.A2(n_816),
.B1(n_1001),
.B2(n_965),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_970),
.B(n_760),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1016),
.A2(n_776),
.B1(n_760),
.B2(n_809),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_910),
.Y(n_1193)
);

BUFx4f_ASAP7_75t_L g1194 ( 
.A(n_920),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_978),
.B(n_760),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_978),
.B(n_760),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_909),
.A2(n_590),
.B(n_765),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_902),
.B(n_883),
.Y(n_1198)
);

CKINVDCx6p67_ASAP7_75t_R g1199 ( 
.A(n_920),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1034),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1034),
.B(n_981),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_910),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_978),
.A2(n_760),
.B(n_802),
.C(n_793),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_978),
.A2(n_760),
.B(n_802),
.C(n_793),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_975),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_902),
.B(n_883),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1034),
.B(n_729),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_1126),
.B(n_1110),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1189),
.B(n_1204),
.C(n_1203),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1102),
.A2(n_1161),
.A3(n_1139),
.B(n_1128),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1111),
.A2(n_1127),
.B(n_1133),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1132),
.A2(n_1186),
.B(n_1182),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1188),
.A2(n_1197),
.B(n_1134),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1195),
.A2(n_1196),
.B(n_1120),
.C(n_1113),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1141),
.A2(n_1116),
.B(n_1172),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1179),
.A2(n_1198),
.B1(n_1206),
.B2(n_1184),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1192),
.A2(n_1146),
.B(n_1088),
.C(n_1144),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_1192),
.A2(n_1102),
.A3(n_1115),
.B1(n_1178),
.B2(n_1139),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1172),
.A2(n_1119),
.B(n_1107),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1167),
.A2(n_1168),
.B(n_1173),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1163),
.A2(n_1122),
.B(n_1149),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1101),
.B(n_1191),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_1068),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1085),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1160),
.A2(n_1074),
.B(n_1073),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1124),
.A2(n_1180),
.B(n_1181),
.C(n_1183),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1085),
.Y(n_1227)
);

CKINVDCx8_ASAP7_75t_R g1228 ( 
.A(n_1136),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1135),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1089),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1114),
.A2(n_1118),
.B1(n_1190),
.B2(n_1142),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1106),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1194),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1140),
.A2(n_1164),
.B(n_1145),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1175),
.A2(n_1170),
.B(n_1174),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1199),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1093),
.B(n_1108),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1205),
.Y(n_1239)
);

BUFx2_ASAP7_75t_SL g1240 ( 
.A(n_1131),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1100),
.A2(n_1166),
.B(n_1148),
.C(n_1095),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1145),
.A2(n_1171),
.B(n_1071),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1117),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1138),
.A2(n_1125),
.B(n_1169),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1086),
.A2(n_1092),
.A3(n_1176),
.B(n_1080),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1109),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1121),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1125),
.A2(n_1159),
.B(n_1064),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1064),
.A2(n_1157),
.B(n_1075),
.C(n_1094),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1250)
);

BUFx2_ASAP7_75t_R g1251 ( 
.A(n_1079),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1194),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1201),
.B(n_1207),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1070),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1165),
.A2(n_1158),
.B(n_1067),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1087),
.A2(n_1076),
.B(n_1082),
.C(n_1105),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1143),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_SL g1258 ( 
.A1(n_1162),
.A2(n_1147),
.B(n_1155),
.C(n_1066),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1147),
.A2(n_1153),
.B(n_1084),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1065),
.A2(n_1123),
.B(n_1078),
.C(n_1129),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1177),
.A2(n_1072),
.B1(n_1077),
.B2(n_1152),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1103),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1090),
.A2(n_1098),
.B(n_1097),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1104),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1156),
.A2(n_1150),
.B(n_1154),
.C(n_1098),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1090),
.A2(n_1097),
.B(n_1207),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1072),
.B(n_1099),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1091),
.A2(n_1078),
.B1(n_1104),
.B2(n_1207),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1137),
.B(n_1151),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1081),
.A2(n_1078),
.B(n_1112),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1131),
.A2(n_1151),
.B(n_1130),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1091),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1091),
.A2(n_1151),
.A3(n_1130),
.B(n_1068),
.Y(n_1273)
);

AOI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1068),
.A2(n_1130),
.B(n_1200),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1200),
.B(n_902),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1200),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1137),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1205),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1069),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_760),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1126),
.A2(n_939),
.A3(n_1102),
.B(n_1161),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1192),
.A2(n_1088),
.B1(n_1204),
.B2(n_1203),
.C(n_1189),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_SL g1287 ( 
.A(n_1079),
.B(n_1096),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1085),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1069),
.Y(n_1289)
);

BUFx4f_ASAP7_75t_L g1290 ( 
.A(n_1199),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1128),
.A2(n_1083),
.B(n_1126),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1126),
.A2(n_939),
.A3(n_1102),
.B(n_1161),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_1195),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1113),
.A2(n_645),
.B1(n_594),
.B2(n_429),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1189),
.A2(n_760),
.B1(n_1204),
.B2(n_1203),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1137),
.Y(n_1297)
);

NOR4xp25_ASAP7_75t_L g1298 ( 
.A(n_1189),
.B(n_1204),
.C(n_1203),
.D(n_1088),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_1136),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1126),
.A2(n_939),
.A3(n_1102),
.B(n_1161),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1113),
.A2(n_929),
.B1(n_965),
.B2(n_760),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_L g1305 ( 
.A1(n_1189),
.A2(n_1204),
.B1(n_1203),
.B2(n_1088),
.C(n_1192),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1185),
.B(n_902),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1126),
.A2(n_939),
.A3(n_1102),
.B(n_1161),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1185),
.B(n_902),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_760),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1189),
.A2(n_760),
.B1(n_1204),
.B2(n_1203),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1189),
.A2(n_760),
.B1(n_1204),
.B2(n_1203),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1113),
.A2(n_760),
.B1(n_1187),
.B2(n_1185),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1131),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1113),
.A2(n_760),
.B1(n_1187),
.B2(n_1185),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1321)
);

BUFx5_ASAP7_75t_L g1322 ( 
.A(n_1170),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1069),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1185),
.B(n_902),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1069),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1185),
.B(n_902),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1189),
.A2(n_760),
.B1(n_1204),
.B2(n_1203),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1192),
.A2(n_1124),
.B(n_1102),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1128),
.A2(n_1083),
.B(n_1126),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1069),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1137),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1113),
.B(n_760),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1113),
.B(n_429),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_1195),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1069),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_760),
.Y(n_1338)
);

AO22x2_ASAP7_75t_L g1339 ( 
.A1(n_1192),
.A2(n_1102),
.B1(n_1088),
.B2(n_1178),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1140),
.A2(n_1149),
.B(n_1160),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1189),
.A2(n_1204),
.B(n_1203),
.C(n_760),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1192),
.A2(n_1088),
.B1(n_1204),
.B2(n_1203),
.C(n_1189),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1189),
.A2(n_760),
.B1(n_1204),
.B2(n_1203),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1161),
.A2(n_1126),
.B(n_1083),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1083),
.A2(n_590),
.B(n_651),
.Y(n_1348)
);

INVx3_ASAP7_75t_SL g1349 ( 
.A(n_1199),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1229),
.A2(n_1339),
.B1(n_1314),
.B2(n_1295),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1349),
.Y(n_1351)
);

BUFx8_ASAP7_75t_L g1352 ( 
.A(n_1230),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1223),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1290),
.Y(n_1354)
);

CKINVDCx11_ASAP7_75t_R g1355 ( 
.A(n_1228),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1316),
.A2(n_1319),
.B1(n_1333),
.B2(n_1232),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1304),
.A2(n_1319),
.B1(n_1316),
.B2(n_1327),
.Y(n_1357)
);

BUFx8_ASAP7_75t_SL g1358 ( 
.A(n_1252),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1299),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1339),
.A2(n_1282),
.B1(n_1343),
.B2(n_1313),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1223),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1234),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1338),
.A2(n_1209),
.B1(n_1324),
.B2(n_1310),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1223),
.B(n_1318),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1227),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1299),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1233),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1315),
.A2(n_1345),
.B1(n_1335),
.B2(n_1209),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1239),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1278),
.A2(n_1330),
.B1(n_1340),
.B2(n_1328),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1318),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1253),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1306),
.A2(n_1326),
.B1(n_1238),
.B2(n_1222),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1294),
.A2(n_1268),
.B1(n_1267),
.B2(n_1264),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1216),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1246),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1290),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1237),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_1254),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1287),
.B(n_1288),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1246),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1231),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1298),
.A2(n_1305),
.B1(n_1218),
.B2(n_1344),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1243),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1247),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1257),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1255),
.A2(n_1248),
.B1(n_1257),
.B2(n_1279),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1280),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1289),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1276),
.Y(n_1391)
);

INVx4_ASAP7_75t_SL g1392 ( 
.A(n_1273),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1275),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1248),
.A2(n_1259),
.B1(n_1215),
.B2(n_1347),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1347),
.A2(n_1262),
.B1(n_1242),
.B2(n_1219),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1261),
.A2(n_1325),
.B1(n_1331),
.B2(n_1337),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1241),
.A2(n_1249),
.B1(n_1226),
.B2(n_1336),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1277),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1269),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1240),
.Y(n_1400)
);

OAI21xp33_ASAP7_75t_L g1401 ( 
.A1(n_1298),
.A2(n_1214),
.B(n_1293),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1297),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1291),
.A2(n_1329),
.B1(n_1208),
.B2(n_1244),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1285),
.A2(n_1270),
.B1(n_1266),
.B2(n_1213),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1273),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1251),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1291),
.A2(n_1329),
.B1(n_1221),
.B2(n_1322),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1332),
.Y(n_1409)
);

BUFx4f_ASAP7_75t_SL g1410 ( 
.A(n_1332),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1273),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1271),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1221),
.A2(n_1322),
.B1(n_1212),
.B2(n_1211),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1245),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1322),
.A2(n_1211),
.B1(n_1235),
.B2(n_1220),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1322),
.A2(n_1236),
.B1(n_1225),
.B2(n_1218),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1274),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1218),
.A2(n_1217),
.B1(n_1256),
.B2(n_1346),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1322),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1263),
.A2(n_1348),
.B1(n_1341),
.B2(n_1334),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1286),
.A2(n_1307),
.B1(n_1303),
.B2(n_1296),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1265),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1245),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1210),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1260),
.B(n_1210),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1317),
.A2(n_1320),
.B1(n_1210),
.B2(n_1301),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1258),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1284),
.A2(n_1309),
.B1(n_1301),
.B2(n_1292),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1281),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1283),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1284),
.A2(n_1292),
.B1(n_1309),
.B2(n_1301),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1284),
.A2(n_1292),
.B(n_1309),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1342),
.B(n_1300),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1302),
.A2(n_1308),
.B1(n_1311),
.B2(n_1312),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1321),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1224),
.Y(n_1436)
);

BUFx5_ASAP7_75t_L g1437 ( 
.A(n_1272),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1318),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1223),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1250),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1209),
.A2(n_1203),
.B(n_1189),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1229),
.A2(n_1192),
.B1(n_1088),
.B2(n_1339),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1250),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1316),
.A2(n_1319),
.B1(n_760),
.B2(n_1229),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1250),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1290),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1228),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1250),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1316),
.A2(n_1319),
.B(n_760),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1229),
.A2(n_1192),
.B1(n_1088),
.B2(n_1339),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1229),
.A2(n_1192),
.B1(n_1088),
.B2(n_1339),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1229),
.A2(n_1192),
.B1(n_1088),
.B2(n_1339),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_SL g1457 ( 
.A(n_1299),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1250),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1290),
.Y(n_1459)
);

BUFx10_ASAP7_75t_L g1460 ( 
.A(n_1237),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1239),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1223),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1250),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1304),
.B2(n_1113),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1223),
.B(n_1131),
.Y(n_1466)
);

BUFx8_ASAP7_75t_SL g1467 ( 
.A(n_1358),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1419),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1406),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1357),
.A2(n_1456),
.B1(n_1465),
.B2(n_1453),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1411),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1390),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1425),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1425),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1414),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1355),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1350),
.B(n_1443),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1392),
.B(n_1423),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1387),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1463),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1433),
.A2(n_1421),
.B(n_1420),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1428),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1430),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1350),
.B(n_1443),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1433),
.A2(n_1415),
.B(n_1404),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1392),
.B(n_1424),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1383),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1413),
.A2(n_1408),
.B(n_1435),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1442),
.A2(n_1450),
.B1(n_1462),
.B2(n_1368),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1432),
.B(n_1375),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1385),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1452),
.B(n_1454),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1432),
.B(n_1360),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1452),
.B(n_1454),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1384),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1455),
.B(n_1384),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1431),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1386),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1360),
.B(n_1441),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1375),
.Y(n_1500)
);

BUFx2_ASAP7_75t_SL g1501 ( 
.A(n_1457),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1389),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1381),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1370),
.B(n_1368),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1437),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1395),
.A2(n_1394),
.B(n_1422),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1445),
.A2(n_1451),
.B1(n_1356),
.B2(n_1401),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1363),
.B(n_1451),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1373),
.B(n_1363),
.Y(n_1510)
);

BUFx2_ASAP7_75t_SL g1511 ( 
.A(n_1457),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1381),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1437),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1430),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1429),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1367),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1380),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1448),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1405),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1418),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1418),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1416),
.A2(n_1396),
.B(n_1388),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1400),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1373),
.A2(n_1427),
.B1(n_1374),
.B2(n_1412),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1393),
.B(n_1438),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1365),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1436),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1440),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1461),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1444),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1426),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1446),
.B(n_1458),
.Y(n_1532)
);

BUFx2_ASAP7_75t_SL g1533 ( 
.A(n_1399),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1449),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1372),
.B(n_1354),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1426),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1464),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1434),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1434),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1364),
.A2(n_1353),
.B(n_1439),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1466),
.A2(n_1439),
.B(n_1361),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1417),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1391),
.A2(n_1407),
.B1(n_1369),
.B2(n_1409),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1378),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1398),
.Y(n_1545)
);

NAND4xp25_ASAP7_75t_L g1546 ( 
.A(n_1508),
.B(n_1377),
.C(n_1402),
.D(n_1376),
.Y(n_1546)
);

NOR2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1351),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1524),
.A2(n_1459),
.B1(n_1447),
.B2(n_1366),
.C(n_1403),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1508),
.A2(n_1382),
.B(n_1359),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1489),
.A2(n_1362),
.B1(n_1352),
.B2(n_1371),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1527),
.Y(n_1552)
);

NOR2x1_ASAP7_75t_R g1553 ( 
.A(n_1544),
.B(n_1362),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1492),
.A2(n_1410),
.B1(n_1379),
.B2(n_1460),
.C(n_1352),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1499),
.A2(n_1493),
.B(n_1470),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1499),
.A2(n_1542),
.B1(n_1509),
.B2(n_1477),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1490),
.B(n_1526),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1531),
.B(n_1536),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1518),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1478),
.B(n_1486),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1509),
.A2(n_1499),
.B(n_1504),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1536),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1534),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1481),
.A2(n_1485),
.B(n_1488),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1487),
.B(n_1491),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_R g1567 ( 
.A(n_1477),
.B(n_1484),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1506),
.A2(n_1481),
.B(n_1519),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1542),
.A2(n_1484),
.B1(n_1493),
.B2(n_1494),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1493),
.B(n_1503),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1473),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1522),
.C(n_1507),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1498),
.B(n_1502),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1485),
.A2(n_1488),
.B(n_1506),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1512),
.B(n_1532),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1473),
.A2(n_1474),
.B(n_1500),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1514),
.B(n_1483),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1468),
.B(n_1541),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1520),
.C(n_1521),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1500),
.A2(n_1540),
.B(n_1541),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1469),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1469),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1497),
.B(n_1516),
.Y(n_1585)
);

AO32x2_ASAP7_75t_L g1586 ( 
.A1(n_1523),
.A2(n_1480),
.A3(n_1543),
.B1(n_1497),
.B2(n_1482),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1535),
.A2(n_1505),
.B(n_1513),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1517),
.B(n_1472),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1538),
.A2(n_1539),
.B(n_1482),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1557),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1583),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1538),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1580),
.B(n_1514),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1584),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1552),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1539),
.Y(n_1596)
);

NAND2x1_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1468),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1515),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1559),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1580),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1559),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1537),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1566),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1468),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1475),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1588),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1589),
.B(n_1471),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1577),
.B(n_1471),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1572),
.B(n_1520),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1585),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1529),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1563),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1564),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1601),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1609),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1616),
.B(n_1578),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1600),
.Y(n_1621)
);

AND2x2_ASAP7_75t_SL g1622 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1592),
.B(n_1569),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1615),
.B(n_1569),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1596),
.B(n_1576),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1591),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1565),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1555),
.Y(n_1630)
);

INVx5_ASAP7_75t_L g1631 ( 
.A(n_1593),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1617),
.B(n_1574),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1594),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1586),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1614),
.A2(n_1554),
.B(n_1549),
.C(n_1548),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1595),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1605),
.A2(n_1550),
.B1(n_1561),
.B2(n_1581),
.C(n_1546),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1613),
.B(n_1587),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1586),
.Y(n_1642)
);

OAI21xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1603),
.A2(n_1567),
.B(n_1547),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1621),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1629),
.B(n_1604),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1637),
.A2(n_1570),
.B1(n_1556),
.B2(n_1533),
.Y(n_1646)
);

INVx5_ASAP7_75t_L g1647 ( 
.A(n_1630),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1642),
.B(n_1611),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1631),
.B(n_1560),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1627),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1607),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1628),
.B(n_1611),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1625),
.B(n_1618),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1560),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1618),
.B(n_1608),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1623),
.B(n_1612),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1620),
.B(n_1632),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1638),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1633),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1624),
.B(n_1606),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1620),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1560),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1639),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1626),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1648),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1646),
.A2(n_1637),
.B(n_1643),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1665),
.B(n_1622),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1665),
.B(n_1622),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1665),
.B(n_1622),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1622),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1646),
.A2(n_1630),
.B(n_1636),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1660),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1661),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1659),
.B(n_1639),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1631),
.Y(n_1678)
);

INVxp33_ASAP7_75t_L g1679 ( 
.A(n_1654),
.Y(n_1679)
);

OR2x6_ASAP7_75t_SL g1680 ( 
.A(n_1659),
.B(n_1632),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1653),
.B(n_1638),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1663),
.B(n_1639),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1661),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1638),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1621),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1651),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1645),
.A2(n_1635),
.B1(n_1643),
.B2(n_1581),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1666),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1666),
.Y(n_1692)
);

AO22x1_ASAP7_75t_L g1693 ( 
.A1(n_1647),
.A2(n_1621),
.B1(n_1644),
.B2(n_1600),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1655),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1657),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1660),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1660),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1650),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1650),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1650),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1677),
.B(n_1658),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1673),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1650),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1668),
.A2(n_1635),
.B1(n_1630),
.B2(n_1621),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1680),
.B(n_1652),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1670),
.B(n_1650),
.Y(n_1710)
);

NOR3xp33_ASAP7_75t_L g1711 ( 
.A(n_1668),
.B(n_1553),
.C(n_1479),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1656),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1700),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1700),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.B(n_1656),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1672),
.B(n_1656),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1683),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1656),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1675),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1688),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1696),
.B(n_1656),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1677),
.B(n_1686),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1652),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1667),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1693),
.B(n_1644),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1667),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1689),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1656),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1685),
.B(n_1664),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1662),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1685),
.B(n_1664),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1691),
.B(n_1662),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1681),
.B(n_1664),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1689),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1690),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1713),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1733),
.B(n_1681),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1713),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1713),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1715),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1711),
.A2(n_1674),
.B(n_1690),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_L g1746 ( 
.A(n_1722),
.B(n_1674),
.C(n_1693),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1726),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1679),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1708),
.A2(n_1687),
.B1(n_1647),
.B2(n_1682),
.C(n_1684),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1708),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1726),
.B(n_1602),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1722),
.A2(n_1630),
.B1(n_1647),
.B2(n_1697),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1715),
.A2(n_1692),
.B(n_1698),
.C(n_1675),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1715),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1736),
.A2(n_1647),
.B1(n_1630),
.B2(n_1682),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1736),
.B(n_1698),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1728),
.Y(n_1760)
);

OAI31xp33_ASAP7_75t_L g1761 ( 
.A1(n_1717),
.A2(n_1678),
.A3(n_1699),
.B(n_1684),
.Y(n_1761)
);

OAI222xp33_ASAP7_75t_L g1762 ( 
.A1(n_1728),
.A2(n_1647),
.B1(n_1630),
.B2(n_1686),
.C1(n_1694),
.C2(n_1701),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1706),
.Y(n_1763)
);

AOI21xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1728),
.A2(n_1678),
.B(n_1467),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1706),
.Y(n_1765)
);

XNOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1739),
.B(n_1747),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1750),
.A2(n_1678),
.B1(n_1728),
.B2(n_1647),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1751),
.B(n_1602),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1753),
.A2(n_1728),
.B(n_1729),
.C(n_1723),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1745),
.A2(n_1678),
.B(n_1734),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1755),
.B(n_1725),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1743),
.Y(n_1772)
);

OAI222xp33_ASAP7_75t_L g1773 ( 
.A1(n_1749),
.A2(n_1756),
.B1(n_1752),
.B2(n_1748),
.C1(n_1760),
.C2(n_1754),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1734),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1746),
.A2(n_1647),
.B(n_1721),
.C(n_1717),
.Y(n_1775)
);

NAND2x1_ASAP7_75t_L g1776 ( 
.A(n_1741),
.B(n_1733),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1751),
.B(n_1721),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1743),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1761),
.A2(n_1647),
.B1(n_1630),
.B2(n_1702),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1758),
.B(n_1705),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1760),
.B(n_1735),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1764),
.B(n_1476),
.Y(n_1782)
);

NAND2xp33_ASAP7_75t_SL g1783 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1742),
.B(n_1735),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1742),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1756),
.A2(n_1737),
.B1(n_1644),
.B2(n_1707),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1782),
.A2(n_1518),
.B1(n_1511),
.B2(n_1501),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1768),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1771),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1772),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1766),
.A2(n_1762),
.B(n_1744),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1781),
.B(n_1737),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1772),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1781),
.B(n_1784),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1776),
.B(n_1740),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1774),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1778),
.B(n_1703),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.B(n_1767),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1769),
.A2(n_1759),
.B(n_1757),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1789),
.B(n_1770),
.C(n_1775),
.D(n_1779),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1791),
.A2(n_1773),
.B(n_1786),
.C(n_1780),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1794),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1783),
.Y(n_1803)
);

NAND4xp25_ASAP7_75t_L g1804 ( 
.A(n_1796),
.B(n_1765),
.C(n_1763),
.D(n_1707),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1787),
.A2(n_1644),
.B1(n_1710),
.B2(n_1703),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1790),
.B(n_1501),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1792),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_SL g1808 ( 
.A(n_1799),
.B(n_1712),
.C(n_1710),
.Y(n_1808)
);

NOR3x1_ASAP7_75t_L g1809 ( 
.A(n_1793),
.B(n_1729),
.C(n_1723),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1788),
.B(n_1511),
.Y(n_1810)
);

OAI31xp33_ASAP7_75t_L g1811 ( 
.A1(n_1800),
.A2(n_1795),
.A3(n_1798),
.B(n_1792),
.Y(n_1811)
);

AND4x1_ASAP7_75t_L g1812 ( 
.A(n_1801),
.B(n_1798),
.C(n_1797),
.D(n_1795),
.Y(n_1812)
);

AOI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1802),
.A2(n_1797),
.B(n_1712),
.C(n_1716),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1807),
.B(n_1716),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1803),
.B(n_1705),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1808),
.A2(n_1810),
.B1(n_1805),
.B2(n_1804),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1811),
.A2(n_1809),
.B1(n_1731),
.B2(n_1738),
.C(n_1719),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1814),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1816),
.A2(n_1812),
.B(n_1815),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1813),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1814),
.Y(n_1821)
);

XNOR2xp5_ASAP7_75t_L g1822 ( 
.A(n_1812),
.B(n_1806),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1815),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1818),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1819),
.B(n_1822),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1823),
.B(n_1724),
.Y(n_1826)
);

BUFx2_ASAP7_75t_SL g1827 ( 
.A(n_1821),
.Y(n_1827)
);

NOR4xp25_ASAP7_75t_L g1828 ( 
.A(n_1820),
.B(n_1730),
.C(n_1727),
.D(n_1731),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1817),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1825),
.B(n_1824),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1826),
.B(n_1738),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1827),
.B(n_1694),
.Y(n_1832)
);

XNOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1830),
.B(n_1832),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1833),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

XNOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1834),
.B(n_1829),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1835),
.A2(n_1834),
.B1(n_1831),
.B2(n_1828),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1836),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1838),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1837),
.A2(n_1730),
.B(n_1727),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1730),
.B1(n_1727),
.B2(n_1714),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1840),
.B(n_1714),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1842),
.B(n_1718),
.Y(n_1843)
);

OR4x1_ASAP7_75t_L g1844 ( 
.A(n_1843),
.B(n_1841),
.C(n_1718),
.D(n_1720),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_R g1845 ( 
.A1(n_1844),
.A2(n_1720),
.B1(n_1719),
.B2(n_1701),
.C(n_1644),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1545),
.B(n_1724),
.C(n_1732),
.Y(n_1846)
);


endmodule