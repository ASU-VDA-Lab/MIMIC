module fake_netlist_1_12743_n_636 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_636);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_636;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_31), .Y(n_78) );
NOR2xp33_ASAP7_75t_L g79 ( .A(n_58), .B(n_45), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_76), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_3), .Y(n_82) );
BUFx2_ASAP7_75t_SL g83 ( .A(n_54), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_63), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_38), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_72), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_37), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_12), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_47), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_73), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_13), .Y(n_99) );
NOR2xp33_ASAP7_75t_L g100 ( .A(n_51), .B(n_26), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_10), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_49), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_24), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_59), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_77), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_25), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_61), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_34), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_71), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_87), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_86), .B(n_0), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_86), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_80), .B(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
BUFx12f_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_89), .B(n_22), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_89), .B(n_23), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_108), .B(n_2), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_119), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_120), .B(n_78), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_120), .B(n_84), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_130), .B(n_82), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_130), .B(n_96), .Y(n_144) );
AOI22xp5_ASAP7_75t_SL g145 ( .A1(n_120), .A2(n_99), .B1(n_81), .B2(n_106), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_125), .B(n_96), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_128), .B(n_98), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_132), .B(n_95), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_132), .B(n_97), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_125), .B(n_110), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_120), .B(n_90), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_124), .B(n_110), .Y(n_157) );
INVxp33_ASAP7_75t_SL g158 ( .A(n_136), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_124), .A2(n_111), .B1(n_107), .B2(n_90), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_119), .Y(n_160) );
INVxp33_ASAP7_75t_SL g161 ( .A(n_127), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_127), .A2(n_92), .B(n_114), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_161), .B(n_154), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_158), .B(n_124), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_156), .B(n_124), .Y(n_170) );
NOR3xp33_ASAP7_75t_L g171 ( .A(n_141), .B(n_129), .C(n_137), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_147), .B(n_129), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_156), .B(n_137), .C(n_126), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_143), .B(n_126), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_142), .A2(n_126), .B(n_91), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_159), .A2(n_126), .B1(n_109), .B2(n_93), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_148), .B(n_117), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_156), .B(n_134), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_164), .B(n_117), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_164), .B(n_94), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_144), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_156), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_157), .B(n_102), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_159), .B(n_134), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
NOR2xp33_ASAP7_75t_SL g193 ( .A(n_164), .B(n_134), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_164), .B(n_116), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_152), .B(n_103), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
NAND2x1_ASAP7_75t_L g197 ( .A(n_165), .B(n_134), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_153), .B(n_104), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_165), .B(n_134), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_167), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_135), .B1(n_134), .B2(n_93), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_145), .B(n_109), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_163), .B(n_115), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_163), .B(n_91), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_138), .B(n_134), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_138), .B(n_83), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_138), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_200), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_204), .A2(n_135), .B(n_114), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_170), .A2(n_92), .B1(n_112), .B2(n_83), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_183), .A2(n_170), .B(n_193), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_187), .B(n_112), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_180), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_186), .B(n_4), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_186), .B(n_105), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_173), .A2(n_113), .B1(n_118), .B2(n_123), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_176), .B(n_135), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_176), .B(n_135), .Y(n_219) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_203), .A2(n_166), .B(n_160), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_168), .B(n_169), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_173), .A2(n_113), .B(n_118), .C(n_123), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_171), .B(n_135), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_172), .B(n_135), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_191), .A2(n_118), .B(n_123), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_187), .B(n_135), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_200), .B(n_135), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_178), .A2(n_79), .B1(n_100), .B2(n_122), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_177), .A2(n_122), .B(n_131), .C(n_150), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_178), .B(n_4), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_179), .A2(n_122), .B1(n_131), .B2(n_150), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_179), .B(n_5), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_183), .A2(n_166), .B(n_160), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_202), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_195), .B(n_5), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_198), .B(n_6), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_182), .B(n_6), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_202), .B(n_7), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g240 ( .A1(n_188), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_193), .B(n_122), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_221), .A2(n_196), .B(n_189), .C(n_192), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_216), .B(n_174), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_216), .B(n_192), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_228), .A2(n_199), .B(n_185), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_233), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_211), .A2(n_194), .B(n_196), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_208), .A2(n_175), .B1(n_181), .B2(n_174), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_239), .B(n_174), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_219), .A2(n_206), .B(n_175), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_227), .A2(n_184), .B(n_205), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_197), .B(n_201), .Y(n_253) );
NOR2xp67_ASAP7_75t_SL g254 ( .A(n_208), .B(n_175), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_215), .A2(n_190), .B1(n_181), .B2(n_206), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_220), .A2(n_197), .B(n_190), .Y(n_257) );
INVx3_ASAP7_75t_SL g258 ( .A(n_235), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_239), .A2(n_190), .B1(n_181), .B2(n_207), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
AOI221x1_ASAP7_75t_L g261 ( .A1(n_210), .A2(n_122), .B1(n_131), .B2(n_207), .C(n_150), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_231), .B(n_8), .Y(n_262) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_229), .B(n_131), .C(n_160), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_166), .B(n_149), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_215), .A2(n_131), .B1(n_11), .B2(n_12), .Y(n_265) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_264), .A2(n_226), .B(n_230), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_250), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_250), .B(n_255), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_264), .A2(n_241), .B(n_209), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_255), .Y(n_270) );
NAND2x1_ASAP7_75t_L g271 ( .A(n_254), .B(n_225), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_255), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_209), .B(n_234), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_224), .B(n_225), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_257), .A2(n_223), .B(n_217), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_249), .A2(n_238), .B(n_236), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_243), .B(n_210), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_263), .A2(n_222), .B(n_219), .Y(n_278) );
NOR2x1_ASAP7_75t_SL g279 ( .A(n_243), .B(n_244), .Y(n_279) );
BUFx4f_ASAP7_75t_SL g280 ( .A(n_258), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_246), .B(n_237), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_253), .A2(n_217), .B(n_218), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_253), .A2(n_232), .B(n_212), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_149), .B(n_140), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_240), .Y(n_286) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_240), .B(n_131), .C(n_140), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_268), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_268), .B(n_248), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_267), .B(n_258), .Y(n_290) );
NOR2x1_ASAP7_75t_L g291 ( .A(n_272), .B(n_265), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_267), .B(n_256), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_279), .B(n_262), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_279), .B(n_251), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_285), .B(n_245), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_285), .B(n_254), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_266), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
OR2x6_ASAP7_75t_L g304 ( .A(n_271), .B(n_252), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_271), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_277), .B(n_10), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_286), .B(n_11), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_266), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_284), .A2(n_149), .B(n_140), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_266), .Y(n_313) );
AO31x2_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_139), .A3(n_14), .B(n_15), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_284), .A2(n_139), .B(n_48), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
OA21x2_ASAP7_75t_L g319 ( .A1(n_275), .A2(n_139), .B(n_46), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_311), .B(n_275), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_311), .B(n_282), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_308), .A2(n_287), .B1(n_281), .B2(n_276), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_313), .B(n_282), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_303), .B(n_281), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_313), .B(n_282), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_308), .B(n_274), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_302), .B(n_273), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_278), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_305), .B(n_273), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_310), .B(n_316), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_305), .B(n_273), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_310), .B(n_316), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_296), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_298), .B(n_278), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_318), .B(n_283), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_318), .B(n_283), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_299), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_283), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_289), .B(n_278), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_309), .B(n_300), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_317), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_305), .B(n_274), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_312), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_289), .B(n_278), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_312), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_309), .A2(n_269), .B1(n_14), .B2(n_15), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_295), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_314), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_295), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_297), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_300), .B(n_269), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_294), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_325), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_326), .B(n_306), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_326), .B(n_306), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_351), .B(n_297), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_366), .B(n_297), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_352), .B(n_290), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_352), .B(n_307), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_328), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_297), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_351), .B(n_359), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_359), .B(n_297), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_359), .B(n_297), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_329), .B(n_290), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_366), .B(n_304), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_328), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_363), .B(n_292), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_304), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_304), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_366), .B(n_304), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_340), .B(n_304), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_363), .B(n_304), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_328), .B(n_312), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_325), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_365), .B(n_319), .Y(n_398) );
NOR2xp33_ASAP7_75t_R g399 ( .A(n_365), .B(n_307), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_325), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_365), .B(n_319), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_348), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_325), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_365), .B(n_319), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_327), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_337), .B(n_319), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_327), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_370), .B(n_291), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_348), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_370), .B(n_291), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_362), .B(n_13), .Y(n_413) );
NOR2x1p5_ASAP7_75t_SL g414 ( .A(n_344), .B(n_319), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_366), .B(n_315), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_337), .B(n_315), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_337), .B(n_315), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_339), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_339), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_327), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_339), .B(n_269), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_334), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_334), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_344), .B(n_16), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_345), .B(n_16), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_345), .B(n_17), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_341), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_341), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_341), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_362), .B(n_17), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_355), .B(n_18), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_350), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_324), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_350), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_355), .B(n_18), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_324), .B(n_19), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_356), .B(n_20), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_381), .B(n_320), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_381), .B(n_357), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_374), .B(n_320), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_374), .B(n_320), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_386), .B(n_324), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_376), .B(n_369), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_371), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_418), .B(n_321), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_372), .B(n_357), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_371), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_SL g451 ( .A1(n_432), .A2(n_364), .B(n_361), .C(n_324), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_419), .B(n_321), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g453 ( .A(n_386), .B(n_324), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_405), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_373), .B(n_361), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_387), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_387), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_380), .B(n_321), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_380), .B(n_323), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_424), .B(n_364), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_382), .B(n_323), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_375), .B(n_338), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_375), .B(n_338), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_424), .B(n_323), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_382), .B(n_330), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_426), .B(n_330), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_399), .Y(n_469) );
AND3x2_ASAP7_75t_L g470 ( .A(n_426), .B(n_338), .C(n_335), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_386), .B(n_331), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_427), .B(n_436), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_377), .B(n_383), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_383), .B(n_332), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_375), .B(n_335), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_335), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_388), .B(n_335), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_413), .A2(n_322), .B1(n_331), .B2(n_354), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_421), .B(n_338), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_385), .B(n_338), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_421), .B(n_333), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_438), .B(n_369), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_439), .B(n_333), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_400), .Y(n_485) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_434), .B(n_354), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_384), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_406), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_378), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_379), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_429), .B(n_346), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_422), .B(n_353), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_422), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_423), .B(n_346), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_406), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_389), .B(n_390), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_389), .B(n_346), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_423), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_390), .B(n_347), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_430), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_430), .B(n_378), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_397), .B(n_353), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_394), .B(n_347), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_397), .B(n_347), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_394), .B(n_349), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_416), .B(n_349), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_416), .B(n_349), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_417), .B(n_354), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_417), .B(n_354), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_431), .A2(n_322), .B1(n_354), .B2(n_358), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_478), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_445), .B(n_393), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_444), .B(n_434), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_496), .B(n_385), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_471), .A2(n_412), .B1(n_410), .B2(n_391), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_487), .B(n_393), .Y(n_517) );
INVxp33_ASAP7_75t_L g518 ( .A(n_489), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_441), .B(n_403), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_469), .B(n_415), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_501), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_453), .A2(n_437), .B(n_415), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_449), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_469), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_482), .B(n_420), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_490), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_479), .B(n_404), .C(n_401), .D(n_398), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_456), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_449), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_482), .B(n_420), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_473), .B(n_437), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_457), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_496), .B(n_385), .Y(n_534) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_444), .A2(n_396), .B1(n_434), .B2(n_401), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_440), .B(n_391), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_463), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_448), .B(n_391), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_455), .B(n_425), .Y(n_539) );
OAI21xp33_ASAP7_75t_SL g540 ( .A1(n_444), .A2(n_407), .B(n_396), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_451), .A2(n_367), .B(n_360), .C(n_358), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_486), .B(n_409), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_451), .A2(n_409), .B(n_408), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_440), .B(n_408), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
OAI33xp33_ASAP7_75t_L g547 ( .A1(n_472), .A2(n_460), .A3(n_484), .B1(n_468), .B2(n_465), .B3(n_483), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_447), .B(n_428), .Y(n_548) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_481), .B(n_433), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_442), .B(n_435), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_442), .B(n_435), .Y(n_551) );
NAND2x2_ASAP7_75t_L g552 ( .A(n_470), .B(n_414), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_498), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_481), .B(n_367), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_452), .B(n_367), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_494), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_491), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_502), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_492), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_443), .B(n_350), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_547), .A2(n_510), .B1(n_470), .B2(n_508), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_540), .B(n_510), .C(n_450), .Y(n_565) );
AOI31xp33_ASAP7_75t_L g566 ( .A1(n_525), .A2(n_481), .A3(n_464), .B(n_475), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_560), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_558), .B(n_506), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_522), .A2(n_462), .B(n_464), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_549), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_514), .B(n_462), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_559), .B(n_507), .Y(n_573) );
OA22x2_ASAP7_75t_L g574 ( .A1(n_520), .A2(n_464), .B1(n_475), .B2(n_443), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_528), .A2(n_485), .B(n_488), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_507), .Y(n_576) );
AOI21xp33_ASAP7_75t_SL g577 ( .A1(n_518), .A2(n_477), .B(n_480), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_528), .A2(n_458), .B1(n_459), .B2(n_461), .C(n_467), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_562), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g580 ( .A1(n_517), .A2(n_509), .B1(n_458), .B2(n_459), .C1(n_461), .C2(n_467), .Y(n_580) );
AOI322xp5_ASAP7_75t_L g581 ( .A1(n_527), .A2(n_474), .A3(n_505), .B1(n_503), .B2(n_499), .C1(n_497), .C2(n_488), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_523), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_524), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_546), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_511), .A2(n_505), .B1(n_503), .B2(n_499), .C(n_497), .Y(n_585) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_516), .A2(n_495), .B(n_27), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_28), .B(n_29), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_552), .A2(n_32), .B1(n_33), .B2(n_35), .C(n_36), .Y(n_589) );
INVxp33_ASAP7_75t_L g590 ( .A(n_532), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_536), .B(n_41), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_564), .A2(n_538), .B(n_543), .C(n_544), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_566), .A2(n_554), .B1(n_545), .B2(n_531), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_564), .A2(n_555), .B1(n_561), .B2(n_521), .Y(n_595) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_581), .A2(n_531), .B(n_557), .C(n_539), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_574), .A2(n_563), .B1(n_515), .B2(n_534), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_578), .A2(n_513), .B1(n_519), .B2(n_548), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_565), .B(n_541), .C(n_529), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_589), .B(n_542), .C(n_537), .Y(n_600) );
AOI322xp5_ASAP7_75t_L g601 ( .A1(n_585), .A2(n_551), .A3(n_550), .B1(n_533), .B2(n_530), .C1(n_43), .C2(n_44), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_567), .B(n_577), .Y(n_602) );
NOR3x1_ASAP7_75t_L g603 ( .A(n_572), .B(n_50), .C(n_53), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_569), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_579), .B(n_580), .Y(n_605) );
OAI222xp33_ASAP7_75t_L g606 ( .A1(n_575), .A2(n_60), .B1(n_65), .B2(n_66), .C1(n_67), .C2(n_69), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g607 ( .A1(n_570), .A2(n_587), .B(n_591), .C(n_571), .Y(n_607) );
NAND3xp33_ASAP7_75t_SL g608 ( .A(n_576), .B(n_568), .C(n_573), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_570), .A2(n_592), .B(n_584), .C(n_588), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g610 ( .A(n_582), .B(n_586), .C(n_589), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_583), .B(n_590), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_574), .A2(n_540), .B1(n_469), .B2(n_565), .Y(n_612) );
OAI211xp5_ASAP7_75t_SL g613 ( .A1(n_581), .A2(n_564), .B(n_578), .C(n_580), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_564), .A2(n_586), .B(n_540), .C(n_581), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_605), .B(n_598), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_613), .B(n_602), .Y(n_616) );
NAND3x1_ASAP7_75t_L g617 ( .A(n_595), .B(n_600), .C(n_612), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_614), .B(n_603), .C(n_607), .D(n_601), .Y(n_618) );
NAND2xp33_ASAP7_75t_SL g619 ( .A(n_610), .B(n_594), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_598), .B(n_608), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_620), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_619), .B(n_593), .C(n_606), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_617), .Y(n_623) );
INVxp33_ASAP7_75t_SL g624 ( .A(n_616), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_623), .B(n_618), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_621), .B(n_615), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_624), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_625), .B(n_622), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_627), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_629), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_628), .B(n_626), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_630), .Y(n_632) );
INVx4_ASAP7_75t_L g633 ( .A(n_632), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_633), .A2(n_631), .B(n_599), .Y(n_634) );
OAI21x1_ASAP7_75t_SL g635 ( .A1(n_634), .A2(n_604), .B(n_597), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_611), .B1(n_609), .B2(n_596), .Y(n_636) );
endmodule