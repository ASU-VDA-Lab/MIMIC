module fake_jpeg_12421_n_292 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_39),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_1),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_75),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_21),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_29),
.B1(n_22),
.B2(n_35),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_74),
.B1(n_80),
.B2(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_22),
.B1(n_35),
.B2(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_32),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_22),
.B1(n_35),
.B2(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_17),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_86),
.B(n_81),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_38),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_26),
.B1(n_28),
.B2(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_97),
.B1(n_37),
.B2(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_98),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_26),
.B1(n_37),
.B2(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_34),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_100),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_23),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_23),
.B1(n_20),
.B2(n_37),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_3),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_128),
.B1(n_109),
.B2(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_37),
.B1(n_4),
.B2(n_6),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_113),
.B1(n_91),
.B2(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_124),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_131),
.Y(n_150)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_63),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_134),
.B(n_138),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_14),
.B(n_11),
.C(n_13),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_100),
.B(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_81),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_66),
.B(n_81),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_132),
.B(n_127),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_82),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_139),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_88),
.B1(n_82),
.B2(n_87),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_87),
.C(n_102),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_91),
.B1(n_67),
.B2(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_166),
.B1(n_172),
.B2(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_167),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_95),
.B(n_88),
.C(n_70),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_110),
.B(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_84),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_94),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_94),
.C(n_67),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_110),
.C(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_113),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_107),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_134),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_139),
.B1(n_128),
.B2(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_129),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_114),
.B(n_111),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_116),
.A2(n_136),
.B1(n_109),
.B2(n_121),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_199),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_143),
.B1(n_152),
.B2(n_141),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_148),
.B(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_177),
.A2(n_202),
.B(n_174),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_185),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_151),
.B1(n_156),
.B2(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_172),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_166),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_159),
.C(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_163),
.C(n_144),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_158),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_208),
.C(n_197),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_216),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_152),
.B1(n_162),
.B2(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_217),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_188),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_150),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_193),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_202),
.B1(n_182),
.B2(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_175),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_183),
.C(n_202),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_236),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_189),
.B(n_183),
.C(n_182),
.D(n_177),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_244),
.B(n_218),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_199),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_242),
.B(n_210),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_191),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_187),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_254),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_214),
.B1(n_220),
.B2(n_205),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_221),
.B(n_223),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_233),
.B(n_232),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_221),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_215),
.C(n_226),
.Y(n_256)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_220),
.C(n_225),
.D(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_233),
.B1(n_232),
.B2(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_235),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_233),
.B(n_211),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_R g270 ( 
.A(n_266),
.B(n_256),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_249),
.C(n_253),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_267),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_265),
.B(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_277),
.A2(n_213),
.B1(n_247),
.B2(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_259),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_282),
.A2(n_283),
.B(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_259),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_283),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_282),
.C(n_273),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_276),
.C(n_279),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_276),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_255),
.Y(n_292)
);


endmodule