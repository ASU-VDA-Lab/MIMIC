module fake_netlist_6_761_n_2465 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2465);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2465;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_1285;
wire n_383;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_56),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_13),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_36),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_170),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_111),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_152),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_10),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_138),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_190),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_73),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_100),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_126),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_221),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_73),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_142),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_54),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_47),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_116),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_225),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_116),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_46),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_51),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_100),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_196),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_203),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_95),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_153),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_72),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_114),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_4),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_89),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_72),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_148),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_133),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_41),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_111),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_34),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_23),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_28),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_105),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_121),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_238),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_77),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_197),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_181),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_206),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_195),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_87),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_165),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_188),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_41),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_155),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_84),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_149),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_51),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_99),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_78),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_239),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_17),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_182),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_121),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_160),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_159),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_141),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_97),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_18),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_200),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_164),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_90),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_163),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_103),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_110),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_146),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_4),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_216),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_176),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_191),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_233),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_108),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_19),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_76),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_63),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_107),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_6),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_46),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_128),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_20),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_231),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_114),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_60),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_66),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_172),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_19),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_48),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_74),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_180),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_43),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_106),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_22),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_144),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_227),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_236),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_145),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_22),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_143),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_107),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_113),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_11),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_171),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_240),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_79),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_17),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_60),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_104),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_179),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_81),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_25),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_48),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_212),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_109),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_80),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_113),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_150),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_26),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_151),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_10),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_80),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_63),
.Y(n_397)
);

BUFx8_ASAP7_75t_SL g398 ( 
.A(n_42),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_118),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_67),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_79),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_87),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_205),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_67),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_213),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_85),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_94),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_194),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_219),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_93),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_110),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_139),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_68),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_96),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_58),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_37),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_162),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_88),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_90),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_103),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_210),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_136),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_82),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_130),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_76),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_70),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_6),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_36),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_175),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_12),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_12),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_177),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_187),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_15),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_109),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_129),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_102),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_23),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_226),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_106),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_7),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_66),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_25),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_28),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_49),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_122),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_77),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_135),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_83),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_40),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_38),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_108),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_83),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_20),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_94),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_88),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_192),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_31),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_92),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_127),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_44),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_122),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_56),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_211),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_119),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_30),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_168),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_119),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_132),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_13),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_118),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_5),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_198),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_319),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_398),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_398),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_312),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_273),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_387),
.B(n_131),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_352),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_288),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_243),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_401),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_288),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_312),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_276),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_286),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_276),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_319),
.B(n_0),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_247),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_286),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_283),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_352),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_249),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_353),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_353),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_283),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_286),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_250),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_252),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_328),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_0),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_328),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_339),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_255),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_469),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_339),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_469),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_286),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_242),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_253),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_283),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_287),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_387),
.B(n_1),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_460),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_460),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_256),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_286),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_286),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_286),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_470),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_258),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_470),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_470),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_264),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_253),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_268),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_265),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_267),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_271),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_295),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_245),
.B(n_254),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_274),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_295),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_281),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_292),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_303),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_295),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_305),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_306),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_307),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_315),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_316),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_245),
.B(n_2),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_323),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_273),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_326),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_329),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_273),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_330),
.Y(n_569)
);

INVxp33_ASAP7_75t_SL g570 ( 
.A(n_244),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_269),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_333),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_393),
.B(n_2),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_269),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_269),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_334),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_337),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_314),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_279),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_314),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_393),
.B(n_3),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_342),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_343),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_254),
.B(n_3),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_345),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_277),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_314),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_331),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_331),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_359),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_331),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_277),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_374),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_363),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_419),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_393),
.B(n_7),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_419),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_367),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_419),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_368),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_369),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_378),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_379),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_384),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_486),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_477),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_478),
.B(n_287),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_494),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_499),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_504),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_512),
.B(n_277),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_531),
.B(n_388),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_500),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_509),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_503),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_500),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_508),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_510),
.Y(n_622)
);

NOR2x1_ASAP7_75t_L g623 ( 
.A(n_501),
.B(n_336),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_515),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_542),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_564),
.B(n_336),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_586),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_527),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_508),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_519),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_524),
.B(n_474),
.Y(n_632)
);

CKINVDCx6p67_ASAP7_75t_R g633 ( 
.A(n_483),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_519),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_528),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_532),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_535),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_528),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_538),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_498),
.B(n_324),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_539),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_529),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_592),
.B(n_394),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_408),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_487),
.A2(n_424),
.B(n_287),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_540),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_545),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_511),
.B(n_324),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_505),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_530),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_501),
.Y(n_653)
);

AND2x2_ASAP7_75t_SL g654 ( 
.A(n_558),
.B(n_424),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_546),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_479),
.B(n_421),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_501),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_507),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_487),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_506),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_571),
.B(n_336),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_597),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_516),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_507),
.Y(n_665)
);

CKINVDCx6p67_ASAP7_75t_R g666 ( 
.A(n_483),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_507),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_522),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_522),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_481),
.B(n_293),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_512),
.B(n_417),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_522),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_597),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_518),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_571),
.B(n_417),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_547),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_549),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_487),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_503),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_553),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_555),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_525),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_523),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_526),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_562),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_573),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_567),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_569),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_574),
.B(n_417),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_517),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_514),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_573),
.B(n_581),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_576),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_577),
.Y(n_697)
);

CKINVDCx11_ASAP7_75t_R g698 ( 
.A(n_502),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_533),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_582),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_513),
.B(n_396),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_570),
.B(n_396),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_534),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_624),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_605),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_660),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_574),
.Y(n_707)
);

CKINVDCx14_ASAP7_75t_R g708 ( 
.A(n_633),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_605),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_654),
.A2(n_584),
.B1(n_596),
.B2(n_514),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_609),
.B(n_671),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_609),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_660),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_618),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_619),
.B(n_475),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_621),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_626),
.A2(n_495),
.B1(n_485),
.B2(n_596),
.Y(n_720)
);

AO22x2_ASAP7_75t_L g721 ( 
.A1(n_626),
.A2(n_424),
.B1(n_279),
.B2(n_335),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_645),
.B(n_585),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_628),
.B(n_601),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_619),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_689),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_663),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_628),
.B(n_603),
.Y(n_727)
);

INVx6_ASAP7_75t_L g728 ( 
.A(n_671),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_618),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_621),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_631),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_644),
.B(n_604),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_660),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_631),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_644),
.B(n_614),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_618),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_671),
.B(n_534),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_645),
.B(n_478),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_614),
.B(n_543),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_638),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_618),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_638),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_663),
.B(n_674),
.Y(n_743)
);

INVx6_ASAP7_75t_L g744 ( 
.A(n_671),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_641),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_674),
.B(n_502),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_640),
.B(n_552),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_671),
.B(n_374),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_646),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_675),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_657),
.B(n_480),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_654),
.A2(n_581),
.B1(n_497),
.B2(n_489),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_679),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_641),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_689),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_651),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_694),
.B(n_575),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_693),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_657),
.B(n_480),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_679),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_652),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_702),
.B(n_557),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_618),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_613),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_654),
.B(n_482),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_646),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_652),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_613),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_686),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_686),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_699),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_675),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_695),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_699),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_693),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_575),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_662),
.B(n_578),
.Y(n_779)
);

AND3x4_ASAP7_75t_L g780 ( 
.A(n_698),
.B(n_476),
.C(n_251),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_654),
.B(n_482),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_646),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_615),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_640),
.B(n_565),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

AO21x2_ASAP7_75t_L g786 ( 
.A1(n_695),
.A2(n_608),
.B(n_670),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_627),
.B(n_484),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_613),
.B(n_374),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_632),
.A2(n_702),
.B1(n_701),
.B2(n_649),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_615),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_703),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_627),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_607),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_613),
.B(n_484),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_632),
.B(n_572),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_615),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_680),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_656),
.B(n_583),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_662),
.B(n_488),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_623),
.B(n_370),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_680),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_680),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_642),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_662),
.B(n_488),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_649),
.A2(n_594),
.B1(n_598),
.B2(n_590),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_642),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_676),
.B(n_490),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_616),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_676),
.B(n_374),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_676),
.B(n_578),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_692),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_692),
.B(n_490),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_616),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_656),
.B(n_600),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_630),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_630),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_670),
.B(n_521),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_630),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_694),
.B(n_580),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_634),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_694),
.B(n_536),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_634),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_634),
.Y(n_825)
);

AND2x6_ASAP7_75t_L g826 ( 
.A(n_692),
.B(n_374),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_701),
.B(n_491),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_635),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_643),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_643),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_643),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_608),
.A2(n_537),
.B1(n_301),
.B2(n_320),
.C(n_280),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_623),
.B(n_580),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_653),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_658),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_658),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_659),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_611),
.B(n_602),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_659),
.B(n_491),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_665),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_665),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_667),
.B(n_587),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_612),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_667),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_668),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_617),
.B(n_370),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_622),
.B(n_392),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_669),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_669),
.B(n_587),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_625),
.B(n_588),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_629),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_672),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_636),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_672),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_673),
.B(n_374),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_673),
.B(n_588),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_637),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_681),
.B(n_492),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_639),
.B(n_589),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_681),
.B(n_599),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_647),
.B(n_293),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_633),
.B(n_599),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_607),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_735),
.B(n_648),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_789),
.A2(n_655),
.B1(n_678),
.B2(n_677),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_726),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_737),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_775),
.B(n_682),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_767),
.A2(n_781),
.B1(n_792),
.B2(n_711),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_723),
.B(n_683),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_775),
.B(n_257),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_727),
.B(n_688),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_747),
.A2(n_784),
.B1(n_851),
.B2(n_849),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_792),
.B(n_589),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_737),
.Y(n_879)
);

AND2x6_ASAP7_75t_SL g880 ( 
.A(n_799),
.B(n_268),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_750),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_737),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_813),
.B(n_257),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_739),
.A2(n_691),
.B1(n_696),
.B2(n_690),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_732),
.B(n_697),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_704),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_766),
.B(n_770),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_750),
.Y(n_888)
);

OR2x4_ASAP7_75t_L g889 ( 
.A(n_854),
.B(n_280),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_750),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_827),
.A2(n_262),
.B(n_282),
.C(n_261),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_845),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_738),
.B(n_700),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_752),
.B(n_467),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_787),
.B(n_261),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_813),
.A2(n_779),
.B1(n_806),
.B2(n_800),
.Y(n_896)
);

AND2x2_ASAP7_75t_SL g897 ( 
.A(n_788),
.B(n_467),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_760),
.B(n_467),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_722),
.B(n_262),
.Y(n_899)
);

NAND3xp33_ASAP7_75t_SL g900 ( 
.A(n_704),
.B(n_251),
.C(n_248),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_863),
.B(n_633),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_778),
.B(n_591),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_786),
.B(n_282),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_786),
.B(n_285),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_786),
.B(n_285),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_847),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_847),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_728),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_809),
.B(n_308),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_712),
.B(n_467),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_712),
.B(n_467),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_847),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_856),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_845),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_778),
.B(n_591),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_861),
.B(n_595),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_845),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_712),
.B(n_467),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_856),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_814),
.B(n_308),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_796),
.B(n_666),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_794),
.B(n_467),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_724),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_713),
.B(n_313),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_707),
.B(n_595),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_853),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_707),
.B(n_666),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_812),
.B(n_666),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_771),
.B(n_772),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_819),
.A2(n_779),
.B1(n_756),
.B2(n_725),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_773),
.B(n_313),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_853),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_685),
.B(n_593),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_812),
.B(n_541),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_802),
.B(n_392),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_860),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_725),
.B(n_698),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_856),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_684),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_819),
.B(n_684),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_724),
.A2(n_248),
.B1(n_309),
.B2(n_284),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_776),
.B(n_318),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_839),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_776),
.B(n_318),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_759),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_819),
.A2(n_429),
.B1(n_432),
.B2(n_422),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_785),
.B(n_340),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_839),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_860),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_819),
.A2(n_429),
.B1(n_436),
.B2(n_433),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_785),
.B(n_340),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_791),
.B(n_718),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_791),
.B(n_344),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_750),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_719),
.B(n_344),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_860),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_762),
.B(n_371),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_753),
.A2(n_296),
.B(n_320),
.C(n_301),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_842),
.A2(n_685),
.B(n_593),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_779),
.A2(n_448),
.B1(n_457),
.B2(n_439),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_728),
.A2(n_373),
.B1(n_403),
.B2(n_371),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_728),
.A2(n_744),
.B1(n_764),
.B2(n_720),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_802),
.B(n_373),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_728),
.A2(n_405),
.B1(n_409),
.B2(n_403),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_777),
.B(n_687),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_802),
.B(n_405),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_763),
.B(n_409),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_758),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_705),
.A2(n_710),
.B(n_709),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_769),
.B(n_412),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_705),
.B(n_412),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_709),
.B(n_464),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_726),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_750),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_710),
.B(n_730),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_744),
.A2(n_473),
.B1(n_464),
.B2(n_492),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_805),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_758),
.B(n_687),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_717),
.B(n_473),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_SL g981 ( 
.A1(n_730),
.A2(n_493),
.B(n_296),
.C(n_338),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_816),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_716),
.A2(n_309),
.B1(n_332),
.B2(n_284),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_731),
.B(n_493),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_731),
.B(n_503),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_134),
.Y(n_986)
);

INVxp33_ASAP7_75t_L g987 ( 
.A(n_743),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_835),
.B(n_541),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_864),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_734),
.B(n_503),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_734),
.B(n_503),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_862),
.A2(n_593),
.B(n_503),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_740),
.B(n_593),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_840),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_743),
.B(n_335),
.Y(n_995)
);

NOR3x1_ASAP7_75t_L g996 ( 
.A(n_746),
.B(n_338),
.C(n_322),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_768),
.B(n_293),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_740),
.B(n_593),
.Y(n_998)
);

INVx8_ASAP7_75t_L g999 ( 
.A(n_811),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_840),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_742),
.B(n_593),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_768),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_768),
.A2(n_782),
.B(n_803),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_744),
.A2(n_355),
.B1(n_293),
.B2(n_341),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_742),
.B(n_544),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_745),
.B(n_544),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_821),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_821),
.A2(n_341),
.B(n_347),
.C(n_322),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_746),
.B(n_664),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_745),
.B(n_548),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_768),
.B(n_347),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_744),
.A2(n_835),
.B1(n_720),
.B2(n_826),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_755),
.B(n_548),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_864),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_717),
.B(n_835),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_755),
.B(n_550),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_823),
.B(n_550),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_757),
.B(n_551),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_757),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_820),
.B(n_551),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_866),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_720),
.A2(n_355),
.B1(n_293),
.B2(n_354),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_866),
.A2(n_260),
.B1(n_263),
.B2(n_246),
.Y(n_1023)
);

NOR2x2_ASAP7_75t_L g1024 ( 
.A(n_823),
.B(n_332),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_820),
.B(n_554),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_820),
.B(n_554),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_768),
.B(n_556),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_720),
.A2(n_355),
.B1(n_365),
.B2(n_354),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_782),
.B(n_556),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_782),
.B(n_559),
.Y(n_1030)
);

AO22x1_ASAP7_75t_L g1031 ( 
.A1(n_780),
.A2(n_356),
.B1(n_362),
.B2(n_350),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_782),
.B(n_355),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_843),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_865),
.B(n_664),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_782),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_836),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_751),
.B(n_270),
.C(n_266),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_803),
.B(n_559),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_807),
.B(n_661),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_823),
.B(n_560),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_803),
.B(n_560),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_823),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_877),
.A2(n_846),
.B1(n_841),
.B2(n_855),
.Y(n_1043)
);

AND3x1_ASAP7_75t_SL g1044 ( 
.A(n_983),
.B(n_356),
.C(n_350),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_900),
.B(n_808),
.C(n_805),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1030),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_892),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_868),
.B(n_795),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_1030),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_887),
.B(n_885),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_914),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_917),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_SL g1055 ( 
.A1(n_874),
.A2(n_708),
.B1(n_795),
.B2(n_857),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_949),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_876),
.B(n_804),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_949),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1030),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_994),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_873),
.B(n_804),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_899),
.B(n_804),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_978),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_888),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_994),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1011),
.A2(n_826),
.B1(n_811),
.B2(n_721),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_974),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_923),
.B(n_927),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_888),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1000),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_982),
.B(n_893),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1000),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1033),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_988),
.B(n_836),
.Y(n_1074)
);

CKINVDCx6p67_ASAP7_75t_R g1075 ( 
.A(n_978),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_988),
.B(n_837),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1015),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_888),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1033),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_888),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_888),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_975),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_870),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_721),
.B1(n_774),
.B2(n_765),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_959),
.A2(n_834),
.B(n_848),
.C(n_837),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_979),
.B(n_808),
.C(n_275),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_906),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_902),
.B(n_848),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_1015),
.B(n_1042),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_906),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_975),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_SL g1092 ( 
.A(n_928),
.B(n_780),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_926),
.B(n_721),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_870),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_907),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_963),
.A2(n_811),
.B1(n_826),
.B2(n_749),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_907),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_912),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1011),
.A2(n_826),
.B1(n_811),
.B2(n_721),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_902),
.B(n_915),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_893),
.B(n_793),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_915),
.B(n_850),
.Y(n_1102)
);

NAND2x1_ASAP7_75t_L g1103 ( 
.A(n_975),
.B(n_715),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_SL g1104 ( 
.A(n_940),
.B(n_278),
.C(n_272),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_947),
.B(n_650),
.C(n_610),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_912),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_878),
.B(n_850),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_870),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_933),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_975),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_881),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_921),
.B(n_867),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_881),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_959),
.A2(n_765),
.B(n_852),
.C(n_843),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1009),
.B(n_1039),
.C(n_966),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_913),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_884),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_881),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_936),
.A2(n_811),
.B1(n_826),
.B2(n_749),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_886),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_880),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_878),
.B(n_852),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_928),
.B(n_795),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_969),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_955),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_913),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_919),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_919),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_939),
.Y(n_1130)
);

NOR2x1_ASAP7_75t_L g1131 ( 
.A(n_872),
.B(n_715),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1019),
.B(n_765),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_955),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_939),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_926),
.B(n_714),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_935),
.B(n_714),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1021),
.B(n_715),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1036),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_937),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1011),
.A2(n_811),
.B1(n_826),
.B2(n_749),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1011),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_955),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1002),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1002),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1002),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_929),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1035),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_908),
.B(n_729),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_929),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_989),
.B(n_858),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_935),
.B(n_714),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_987),
.B(n_610),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_869),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_950),
.B(n_729),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_908),
.B(n_729),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_957),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1011),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_969),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1011),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_871),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_941),
.B(n_290),
.C(n_289),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1007),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_987),
.B(n_650),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_879),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_882),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_938),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1023),
.B(n_294),
.C(n_291),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1035),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1027),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1042),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_970),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1034),
.B(n_298),
.C(n_297),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1008),
.B(n_300),
.C(n_299),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_999),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_995),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1029),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_995),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_R g1179 ( 
.A(n_901),
.B(n_661),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_924),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1014),
.B(n_736),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1007),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_889),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1008),
.B(n_304),
.C(n_302),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1038),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_890),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1021),
.B(n_736),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_1017),
.B(n_365),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_976),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1005),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_897),
.A2(n_1012),
.B1(n_936),
.B2(n_1017),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_883),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1040),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_908),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1040),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_883),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_875),
.B(n_858),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_953),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1006),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_SL g1201 ( 
.A(n_951),
.B(n_418),
.C(n_411),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_999),
.B(n_736),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1010),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_931),
.B(n_741),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_980),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_930),
.B(n_741),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1028),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_964),
.A2(n_749),
.B1(n_741),
.B2(n_838),
.Y(n_1208)
);

BUFx4f_ASAP7_75t_L g1209 ( 
.A(n_980),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_942),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_986),
.B(n_706),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_897),
.B(n_706),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1013),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_872),
.B(n_311),
.C(n_310),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_889),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_875),
.B(n_733),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_946),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_R g1218 ( 
.A(n_875),
.B(n_317),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1024),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1016),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_875),
.B(n_411),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1018),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_984),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_925),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_916),
.B(n_733),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1041),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1020),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1024),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_895),
.B(n_748),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_961),
.B(n_838),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_943),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_999),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_910),
.B(n_748),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_999),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_964),
.B(n_838),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_910),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_SL g1237 ( 
.A(n_1022),
.B(n_425),
.C(n_418),
.Y(n_1237)
);

AOI31xp67_ASAP7_75t_L g1238 ( 
.A1(n_1170),
.A2(n_898),
.A3(n_894),
.B(n_903),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1061),
.A2(n_905),
.B(n_904),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1148),
.A2(n_1003),
.B(n_918),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1210),
.A2(n_1031),
.B1(n_1037),
.B2(n_459),
.C(n_437),
.Y(n_1241)
);

OAI21xp33_ASAP7_75t_L g1242 ( 
.A1(n_1176),
.A2(n_1004),
.B(n_956),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1141),
.A2(n_922),
.B(n_918),
.Y(n_1243)
);

OAI22x1_ASAP7_75t_L g1244 ( 
.A1(n_1210),
.A2(n_967),
.B1(n_1032),
.B2(n_997),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1050),
.B(n_932),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1103),
.A2(n_911),
.B(n_985),
.Y(n_1246)
);

INVx3_ASAP7_75t_SL g1247 ( 
.A(n_1075),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1172),
.A2(n_1032),
.B(n_997),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1178),
.B(n_996),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1148),
.A2(n_911),
.B(n_967),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1189),
.B(n_1199),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1063),
.B(n_425),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1148),
.A2(n_1026),
.B(n_1025),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1189),
.B(n_958),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1100),
.B(n_909),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1194),
.B(n_920),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1115),
.A2(n_945),
.A3(n_952),
.B(n_948),
.Y(n_1257)
);

AOI221xp5_ASAP7_75t_L g1258 ( 
.A1(n_1221),
.A2(n_437),
.B1(n_459),
.B2(n_430),
.C(n_428),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1087),
.Y(n_1259)
);

AND2x6_ASAP7_75t_L g1260 ( 
.A(n_1234),
.B(n_977),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1156),
.A2(n_922),
.B(n_898),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1067),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1199),
.B(n_968),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1103),
.A2(n_991),
.B(n_990),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1156),
.A2(n_894),
.B(n_993),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1156),
.A2(n_1001),
.B(n_998),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1078),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1071),
.B(n_954),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1146),
.B(n_971),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1087),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1172),
.A2(n_891),
.B(n_972),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1093),
.A2(n_973),
.B(n_965),
.C(n_962),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1084),
.A2(n_934),
.A3(n_810),
.B(n_832),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1078),
.B(n_362),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1113),
.B(n_321),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1046),
.B(n_838),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1095),
.Y(n_1277)
);

AOI221x1_ASAP7_75t_L g1278 ( 
.A1(n_1237),
.A2(n_960),
.B1(n_801),
.B2(n_832),
.C(n_810),
.Y(n_1278)
);

INVx5_ASAP7_75t_L g1279 ( 
.A(n_1078),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1046),
.B(n_1059),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1190),
.B(n_754),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_1108),
.B(n_375),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1190),
.B(n_754),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1170),
.A2(n_833),
.A3(n_801),
.B(n_790),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1230),
.A2(n_833),
.B(n_822),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1204),
.A2(n_824),
.B(n_815),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1146),
.B(n_259),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1235),
.A2(n_992),
.B(n_790),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1207),
.A2(n_440),
.B1(n_377),
.B2(n_259),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1057),
.A2(n_797),
.B(n_783),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1212),
.A2(n_761),
.B(n_749),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1093),
.A2(n_415),
.B(n_375),
.C(n_380),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1203),
.B(n_761),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1079),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1195),
.A2(n_831),
.B(n_830),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1195),
.A2(n_831),
.B(n_830),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1059),
.B(n_838),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1177),
.A2(n_749),
.B(n_783),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1153),
.B(n_1164),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1203),
.B(n_797),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1141),
.A2(n_825),
.B(n_818),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1158),
.A2(n_825),
.B(n_818),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1063),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1177),
.A2(n_828),
.A3(n_829),
.B(n_381),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1158),
.A2(n_829),
.B(n_828),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1136),
.A2(n_817),
.B(n_981),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1195),
.A2(n_831),
.B(n_830),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1213),
.B(n_1220),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1217),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1213),
.B(n_817),
.Y(n_1310)
);

INVx3_ASAP7_75t_SL g1311 ( 
.A(n_1075),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1078),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1160),
.A2(n_817),
.B(n_563),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1079),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1098),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1220),
.B(n_844),
.Y(n_1316)
);

NAND2x1_ASAP7_75t_L g1317 ( 
.A(n_1064),
.B(n_830),
.Y(n_1317)
);

NAND3x1_ASAP7_75t_L g1318 ( 
.A(n_1043),
.B(n_381),
.C(n_380),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1223),
.B(n_844),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1160),
.A2(n_444),
.A3(n_382),
.B(n_390),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1217),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1067),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1223),
.A2(n_1192),
.B(n_1085),
.C(n_1231),
.Y(n_1323)
);

AOI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1101),
.A2(n_981),
.B(n_327),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1186),
.B(n_844),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1159),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1206),
.A2(n_1062),
.B(n_1175),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1236),
.B(n_844),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1175),
.A2(n_831),
.B(n_830),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1233),
.A2(n_563),
.B(n_561),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1152),
.A2(n_1135),
.B(n_1096),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1074),
.A2(n_859),
.B(n_798),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1233),
.A2(n_566),
.B(n_561),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1175),
.B(n_844),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1175),
.A2(n_831),
.B(n_798),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1200),
.B(n_325),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1159),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1226),
.A2(n_423),
.A3(n_390),
.B(n_472),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1053),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1185),
.A2(n_566),
.B(n_395),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1138),
.A2(n_472),
.B(n_454),
.C(n_427),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1200),
.B(n_346),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1222),
.B(n_1224),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1232),
.A2(n_1097),
.B(n_1090),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1232),
.A2(n_395),
.B(n_382),
.Y(n_1345)
);

NOR2xp67_ASAP7_75t_SL g1346 ( 
.A(n_1175),
.B(n_410),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_SL g1347 ( 
.A(n_1179),
.B(n_349),
.C(n_348),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1232),
.A2(n_415),
.B(n_410),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1226),
.A2(n_798),
.B(n_423),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1149),
.B(n_351),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1163),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1078),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1121),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1090),
.A2(n_427),
.B(n_420),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1097),
.A2(n_438),
.B(n_420),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1196),
.A2(n_355),
.B1(n_859),
.B2(n_471),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1117),
.A2(n_444),
.B(n_438),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_357),
.Y(n_1358)
);

NAND3x1_ASAP7_75t_L g1359 ( 
.A(n_1138),
.B(n_454),
.C(n_453),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1149),
.B(n_1116),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1201),
.B(n_358),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1215),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1076),
.A2(n_859),
.B(n_798),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1088),
.A2(n_1102),
.B(n_1209),
.C(n_1123),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1209),
.A2(n_453),
.B(n_407),
.C(n_406),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1089),
.B(n_137),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1089),
.B(n_140),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1227),
.A2(n_859),
.A3(n_9),
.B(n_11),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1064),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1163),
.B(n_259),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1049),
.A2(n_431),
.B1(n_361),
.B2(n_466),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1048),
.B(n_147),
.Y(n_1372)
);

AO21x1_ASAP7_75t_L g1373 ( 
.A1(n_1233),
.A2(n_8),
.B(n_9),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1117),
.A2(n_798),
.B(n_859),
.Y(n_1374)
);

AOI211x1_ASAP7_75t_L g1375 ( 
.A1(n_1165),
.A2(n_259),
.B(n_377),
.C(n_440),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1224),
.B(n_360),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1129),
.A2(n_859),
.B(n_234),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1106),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1227),
.A2(n_157),
.B(n_158),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1129),
.A2(n_224),
.B(n_222),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1125),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1106),
.A2(n_8),
.A3(n_14),
.B(n_15),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1121),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1130),
.A2(n_220),
.B(n_217),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1127),
.A2(n_14),
.A3(n_18),
.B(n_21),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1130),
.A2(n_215),
.B(n_207),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1092),
.A2(n_463),
.B1(n_462),
.B2(n_461),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1105),
.B(n_364),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1089),
.B(n_161),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1209),
.A2(n_458),
.B(n_456),
.C(n_455),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1107),
.B(n_366),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1180),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_SL g1393 ( 
.A(n_1118),
.B(n_259),
.Y(n_1393)
);

OAI22x1_ASAP7_75t_L g1394 ( 
.A1(n_1118),
.A2(n_452),
.B1(n_451),
.B2(n_449),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1127),
.A2(n_447),
.B(n_446),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1142),
.A2(n_202),
.B(n_201),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1182),
.B(n_377),
.Y(n_1397)
);

AOI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1207),
.A2(n_402),
.B1(n_443),
.B2(n_442),
.C(n_441),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1142),
.A2(n_193),
.B(n_189),
.Y(n_1399)
);

BUFx4_ASAP7_75t_SL g1400 ( 
.A(n_1083),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1143),
.A2(n_186),
.B(n_185),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1049),
.A2(n_1229),
.B(n_1208),
.Y(n_1402)
);

AOI211x1_ASAP7_75t_L g1403 ( 
.A1(n_1165),
.A2(n_377),
.B(n_440),
.C(n_435),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1053),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1181),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1308),
.B(n_1205),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1366),
.B(n_1077),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1339),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1344),
.A2(n_1091),
.B(n_1069),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1264),
.A2(n_1091),
.B(n_1069),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1327),
.A2(n_1080),
.B(n_1064),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1290),
.A2(n_1225),
.B(n_1211),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1292),
.A2(n_1099),
.B1(n_1066),
.B2(n_1150),
.C(n_1047),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1275),
.A2(n_1154),
.B1(n_1361),
.B2(n_1318),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1301),
.A2(n_1091),
.B(n_1069),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1321),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1364),
.A2(n_1056),
.B(n_1054),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1339),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1251),
.A2(n_1193),
.B1(n_1197),
.B2(n_1154),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1366),
.B(n_1077),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1404),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1404),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1393),
.B(n_1080),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_SL g1424 ( 
.A(n_1282),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1309),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1248),
.A2(n_1191),
.B(n_1185),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1294),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1369),
.B(n_1080),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1302),
.A2(n_1111),
.B(n_1109),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1313),
.A2(n_1240),
.B(n_1305),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1364),
.A2(n_1056),
.B(n_1054),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1294),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1246),
.A2(n_1111),
.B(n_1109),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1323),
.A2(n_1131),
.B(n_1198),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1275),
.A2(n_1215),
.B1(n_1228),
.B2(n_1219),
.Y(n_1435)
);

INVx6_ASAP7_75t_L g1436 ( 
.A(n_1369),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1245),
.A2(n_1197),
.B1(n_1193),
.B2(n_1236),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1323),
.A2(n_1198),
.B(n_1216),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1285),
.A2(n_1111),
.B(n_1109),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1400),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1309),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1331),
.A2(n_1402),
.B(n_1268),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1254),
.A2(n_1236),
.B1(n_1139),
.B2(n_1157),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1314),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1259),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1266),
.A2(n_1133),
.B(n_1191),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1306),
.A2(n_1255),
.B(n_1261),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1269),
.B(n_1263),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1351),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1289),
.B(n_1168),
.C(n_1086),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1255),
.A2(n_1229),
.B(n_1132),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1351),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1243),
.A2(n_1133),
.B(n_1143),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1337),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1373),
.A2(n_1205),
.B(n_1081),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1253),
.A2(n_1120),
.B(n_1137),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1400),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1361),
.A2(n_1228),
.B1(n_1139),
.B2(n_1157),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1366),
.B(n_1068),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1270),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1243),
.A2(n_1133),
.B(n_1144),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1286),
.A2(n_1147),
.B(n_1144),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1277),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1268),
.A2(n_1216),
.B(n_1150),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1405),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1315),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1405),
.A2(n_1236),
.B1(n_1181),
.B2(n_1161),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_SL g1469 ( 
.A1(n_1250),
.A2(n_1081),
.B(n_1147),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1343),
.B(n_1360),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1369),
.A2(n_1081),
.B(n_1082),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1354),
.A2(n_1151),
.B(n_1134),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1272),
.A2(n_1166),
.B(n_1068),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1279),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1353),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1258),
.A2(n_1188),
.B1(n_1045),
.B2(n_1055),
.C(n_1173),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1272),
.A2(n_1166),
.B(n_1068),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1291),
.A2(n_1052),
.B(n_1051),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1355),
.A2(n_1151),
.B(n_1134),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1357),
.A2(n_1128),
.B(n_1073),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1378),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1299),
.B(n_1180),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1337),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1281),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1256),
.A2(n_1236),
.B1(n_1181),
.B2(n_1161),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1391),
.B(n_1089),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1303),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1367),
.B(n_1171),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1239),
.A2(n_1128),
.B(n_1065),
.Y(n_1489)
);

BUFx2_ASAP7_75t_R g1490 ( 
.A(n_1247),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1265),
.A2(n_1288),
.B(n_1330),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1330),
.A2(n_1073),
.B(n_1058),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1252),
.A2(n_1218),
.B1(n_1108),
.B2(n_1094),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1283),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1333),
.A2(n_1058),
.B(n_1072),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1333),
.A2(n_1060),
.B(n_1065),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1241),
.A2(n_1183),
.B1(n_1110),
.B2(n_1171),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1377),
.A2(n_1060),
.B(n_1072),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1381),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1289),
.B(n_1214),
.C(n_1104),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1278),
.A2(n_1070),
.B(n_1184),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1345),
.A2(n_1070),
.B(n_1174),
.Y(n_1502)
);

AO221x2_ASAP7_75t_L g1503 ( 
.A1(n_1244),
.A2(n_1044),
.B1(n_440),
.B2(n_377),
.C(n_1162),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1380),
.A2(n_1187),
.B(n_1124),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1284),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1367),
.B(n_1155),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1292),
.A2(n_1119),
.A3(n_1169),
.B(n_1094),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1293),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1332),
.A2(n_1211),
.B(n_1155),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1249),
.A2(n_1388),
.B1(n_1324),
.B2(n_1394),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1384),
.A2(n_1140),
.B(n_1169),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1386),
.A2(n_1399),
.B(n_1396),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1284),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1284),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1398),
.B(n_434),
.C(n_376),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1365),
.A2(n_1211),
.B(n_1155),
.C(n_1083),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1401),
.A2(n_1119),
.B(n_1169),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1300),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1348),
.A2(n_1119),
.B(n_1112),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1369),
.A2(n_1234),
.B1(n_1202),
.B2(n_1112),
.Y(n_1520)
);

OAI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1387),
.A2(n_416),
.B1(n_383),
.B2(n_385),
.C(n_386),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1284),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1340),
.A2(n_1112),
.B(n_1114),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1367),
.B(n_1112),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1304),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1336),
.B(n_1183),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1374),
.A2(n_1112),
.B(n_1114),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1365),
.B(n_426),
.C(n_389),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1242),
.A2(n_1234),
.B(n_1114),
.C(n_1126),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1329),
.A2(n_1114),
.B(n_1126),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1389),
.B(n_1183),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1304),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1304),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1389),
.B(n_1114),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1326),
.A2(n_1234),
.B1(n_1202),
.B2(n_1145),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1347),
.A2(n_1167),
.B1(n_1122),
.B2(n_1145),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1280),
.A2(n_1202),
.B(n_400),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1287),
.A2(n_1167),
.B1(n_1122),
.B2(n_1145),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1328),
.A2(n_1202),
.B(n_1145),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1381),
.Y(n_1540)
);

OAI222xp33_ASAP7_75t_L g1541 ( 
.A1(n_1282),
.A2(n_404),
.B1(n_445),
.B2(n_391),
.C1(n_414),
.C2(n_413),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1304),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1389),
.B(n_1126),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1350),
.A2(n_372),
.B1(n_397),
.B2(n_399),
.C(n_1167),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1279),
.B(n_1234),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1383),
.Y(n_1546)
);

AO21x2_ASAP7_75t_L g1547 ( 
.A1(n_1363),
.A2(n_1145),
.B(n_1126),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1342),
.B(n_1126),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1362),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1280),
.A2(n_440),
.B(n_184),
.Y(n_1550)
);

OR2x6_ASAP7_75t_SL g1551 ( 
.A(n_1358),
.B(n_21),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1273),
.B(n_24),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1295),
.A2(n_183),
.B(n_178),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_SL g1554 ( 
.A1(n_1379),
.A2(n_174),
.B(n_169),
.Y(n_1554)
);

INVx4_ASAP7_75t_SL g1555 ( 
.A(n_1260),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1326),
.A2(n_1319),
.B1(n_1316),
.B2(n_1325),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1298),
.A2(n_24),
.B(n_26),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1310),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1257),
.Y(n_1559)
);

AOI21xp33_ASAP7_75t_L g1560 ( 
.A1(n_1376),
.A2(n_27),
.B(n_29),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1257),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1296),
.A2(n_166),
.B(n_29),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1303),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1307),
.A2(n_27),
.B(n_30),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_SL g1565 ( 
.A(n_1279),
.B(n_31),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1312),
.B(n_32),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1262),
.Y(n_1567)
);

BUFx8_ASAP7_75t_SL g1568 ( 
.A(n_1282),
.Y(n_1568)
);

BUFx4f_ASAP7_75t_L g1569 ( 
.A(n_1267),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1370),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1338),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1312),
.B(n_33),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1257),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1335),
.A2(n_35),
.B(n_38),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1338),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_SL g1576 ( 
.A1(n_1395),
.A2(n_39),
.B(n_40),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1273),
.B(n_39),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1262),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1279),
.Y(n_1579)
);

NAND2x1_ASAP7_75t_L g1580 ( 
.A(n_1267),
.B(n_43),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1267),
.B(n_44),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1322),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1257),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1338),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1341),
.A2(n_45),
.B(n_47),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1322),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1328),
.A2(n_45),
.B(n_49),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1334),
.A2(n_50),
.B(n_52),
.Y(n_1588)
);

INVx8_ASAP7_75t_L g1589 ( 
.A(n_1267),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1334),
.A2(n_50),
.B(n_53),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1440),
.B(n_1395),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1423),
.A2(n_1260),
.B1(n_1392),
.B2(n_1397),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1414),
.A2(n_1318),
.B1(n_1247),
.B2(n_1311),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1427),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1455),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1423),
.A2(n_1260),
.B1(n_1371),
.B2(n_1395),
.Y(n_1596)
);

AND2x2_ASAP7_75t_SL g1597 ( 
.A(n_1414),
.B(n_1352),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1512),
.A2(n_1349),
.B(n_1276),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_SL g1599 ( 
.A(n_1451),
.B(n_1390),
.C(n_1341),
.Y(n_1599)
);

AOI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1412),
.A2(n_1346),
.B(n_1271),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1428),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1451),
.A2(n_1372),
.B1(n_1274),
.B2(n_1311),
.Y(n_1602)
);

INVxp33_ASAP7_75t_L g1603 ( 
.A(n_1482),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1559),
.B(n_1273),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1500),
.A2(n_1274),
.B1(n_1260),
.B2(n_1356),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1474),
.B(n_1352),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1461),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1449),
.B(n_1390),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1449),
.B(n_1320),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1428),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1416),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1427),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1557),
.B(n_1352),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1440),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1550),
.A2(n_1442),
.B(n_1477),
.C(n_1473),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1510),
.A2(n_1276),
.B1(n_1297),
.B2(n_1271),
.C(n_1317),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1458),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1450),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1444),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1436),
.Y(n_1620)
);

BUFx12f_ASAP7_75t_L g1621 ( 
.A(n_1458),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1470),
.B(n_1359),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1500),
.B(n_1359),
.C(n_1403),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1444),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1470),
.B(n_1375),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1476),
.A2(n_1297),
.B(n_1320),
.C(n_1385),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1490),
.Y(n_1627)
);

INVx4_ASAP7_75t_L g1628 ( 
.A(n_1436),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1487),
.Y(n_1629)
);

INVx4_ASAP7_75t_L g1630 ( 
.A(n_1436),
.Y(n_1630)
);

OAI222xp33_ASAP7_75t_L g1631 ( 
.A1(n_1570),
.A2(n_1385),
.B1(n_1382),
.B2(n_55),
.C1(n_57),
.C2(n_58),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1448),
.A2(n_1271),
.B(n_1352),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1455),
.Y(n_1633)
);

OR2x6_ASAP7_75t_SL g1634 ( 
.A(n_1528),
.B(n_1486),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1408),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1559),
.B(n_1273),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1484),
.B(n_1338),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1461),
.Y(n_1638)
);

AO31x2_ASAP7_75t_L g1639 ( 
.A1(n_1561),
.A2(n_1573),
.A3(n_1583),
.B(n_1575),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1563),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1408),
.Y(n_1641)
);

CKINVDCx16_ASAP7_75t_R g1642 ( 
.A(n_1455),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1512),
.A2(n_1238),
.B(n_1320),
.Y(n_1643)
);

AND2x4_ASAP7_75t_SL g1644 ( 
.A(n_1407),
.B(n_1260),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1577),
.B(n_1320),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1577),
.B(n_1385),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1515),
.A2(n_1385),
.B1(n_1382),
.B2(n_1368),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1474),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1436),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1450),
.Y(n_1650)
);

BUFx8_ASAP7_75t_L g1651 ( 
.A(n_1531),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1460),
.B(n_1368),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1484),
.B(n_1382),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1526),
.A2(n_1368),
.B1(n_1382),
.B2(n_55),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1418),
.B(n_1368),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_SL g1656 ( 
.A(n_1521),
.B(n_53),
.C(n_54),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1418),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1515),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1503),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1503),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1467),
.Y(n_1661)
);

INVx6_ASAP7_75t_L g1662 ( 
.A(n_1474),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1467),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1503),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_1664)
);

NAND2x1p5_ASAP7_75t_L g1665 ( 
.A(n_1474),
.B(n_1579),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1481),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1421),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1421),
.B(n_69),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1460),
.B(n_70),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1422),
.B(n_71),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1481),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1460),
.B(n_71),
.Y(n_1672)
);

BUFx4f_ASAP7_75t_L g1673 ( 
.A(n_1474),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1422),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1432),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1568),
.Y(n_1676)
);

OAI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1544),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.C(n_81),
.Y(n_1677)
);

BUFx8_ASAP7_75t_SL g1678 ( 
.A(n_1549),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1446),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1516),
.B(n_75),
.C(n_82),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1432),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1579),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1549),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1541),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.C(n_89),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1503),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_R g1686 ( 
.A1(n_1419),
.A2(n_91),
.B(n_93),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_SL g1687 ( 
.A1(n_1529),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_1687)
);

INVx3_ASAP7_75t_SL g1688 ( 
.A(n_1546),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1494),
.B(n_98),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1446),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1534),
.B(n_98),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1528),
.A2(n_124),
.B1(n_101),
.B2(n_102),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1534),
.B(n_99),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1543),
.B(n_101),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1494),
.B(n_104),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1445),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1464),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1491),
.A2(n_105),
.B(n_112),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1445),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1483),
.Y(n_1700)
);

OAI211xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1435),
.A2(n_112),
.B(n_115),
.C(n_117),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1464),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1560),
.A2(n_115),
.B1(n_117),
.B2(n_120),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1425),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1406),
.B(n_1486),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1540),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1483),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1459),
.A2(n_1497),
.B1(n_1538),
.B2(n_1536),
.C(n_1475),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1579),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1453),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1460),
.A2(n_1493),
.B1(n_1506),
.B2(n_1438),
.Y(n_1711)
);

CKINVDCx16_ASAP7_75t_R g1712 ( 
.A(n_1483),
.Y(n_1712)
);

BUFx10_ASAP7_75t_L g1713 ( 
.A(n_1579),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1428),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1525),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1579),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1448),
.A2(n_120),
.B(n_123),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1546),
.A2(n_1407),
.B1(n_1420),
.B2(n_1506),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1582),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1531),
.A2(n_1506),
.B1(n_1488),
.B2(n_1420),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1506),
.A2(n_123),
.B1(n_124),
.B2(n_1488),
.Y(n_1721)
);

INVx4_ASAP7_75t_SL g1722 ( 
.A(n_1507),
.Y(n_1722)
);

INVx4_ASAP7_75t_SL g1723 ( 
.A(n_1507),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1543),
.B(n_1465),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1582),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1578),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1424),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1499),
.Y(n_1728)
);

OR2x4_ASAP7_75t_L g1729 ( 
.A(n_1552),
.B(n_1548),
.Y(n_1729)
);

AO22x2_ASAP7_75t_L g1730 ( 
.A1(n_1561),
.A2(n_1583),
.B1(n_1573),
.B2(n_1555),
.Y(n_1730)
);

OAI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1551),
.A2(n_1406),
.B1(n_1499),
.B2(n_1580),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1578),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1407),
.B(n_1420),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1466),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1542),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1589),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1407),
.A2(n_1420),
.B1(n_1488),
.B2(n_1443),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1488),
.A2(n_1581),
.B1(n_1572),
.B2(n_1566),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1567),
.Y(n_1739)
);

OAI22x1_ASAP7_75t_L g1740 ( 
.A1(n_1585),
.A2(n_1557),
.B1(n_1575),
.B2(n_1571),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1411),
.A2(n_1434),
.B(n_1509),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1581),
.A2(n_1572),
.B1(n_1566),
.B2(n_1565),
.Y(n_1742)
);

BUFx8_ASAP7_75t_SL g1743 ( 
.A(n_1569),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1552),
.B(n_1558),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1508),
.B(n_1518),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1586),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1508),
.B(n_1518),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1564),
.A2(n_1537),
.B1(n_1580),
.B2(n_1441),
.C(n_1452),
.Y(n_1748)
);

CKINVDCx14_ASAP7_75t_R g1749 ( 
.A(n_1424),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1576),
.A2(n_1556),
.B1(n_1413),
.B2(n_1565),
.C(n_1452),
.Y(n_1751)
);

INVx4_ASAP7_75t_SL g1752 ( 
.A(n_1507),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1478),
.A2(n_1485),
.B1(n_1437),
.B2(n_1413),
.C(n_1468),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_L g1754 ( 
.A(n_1545),
.B(n_1520),
.Y(n_1754)
);

CKINVDCx11_ASAP7_75t_R g1755 ( 
.A(n_1551),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1571),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1509),
.A2(n_1471),
.B(n_1489),
.Y(n_1757)
);

AOI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1456),
.A2(n_1501),
.B(n_1426),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1576),
.A2(n_1554),
.B1(n_1456),
.B2(n_1581),
.C(n_1489),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_L g1760 ( 
.A(n_1585),
.B(n_1566),
.C(n_1572),
.Y(n_1760)
);

AOI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1412),
.A2(n_1539),
.B(n_1533),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1524),
.A2(n_1566),
.B1(n_1572),
.B2(n_1581),
.Y(n_1762)
);

AO21x2_ASAP7_75t_L g1763 ( 
.A1(n_1584),
.A2(n_1491),
.B(n_1533),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1589),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1532),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1555),
.B(n_1524),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1589),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1509),
.A2(n_1547),
.B(n_1457),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1505),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1524),
.A2(n_1555),
.B1(n_1557),
.B2(n_1554),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1569),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1555),
.B(n_1507),
.Y(n_1772)
);

AND2x2_ASAP7_75t_SL g1773 ( 
.A(n_1557),
.B(n_1585),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1589),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1569),
.A2(n_1535),
.B1(n_1545),
.B2(n_1417),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1589),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1501),
.A2(n_1426),
.B1(n_1502),
.B2(n_1585),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1507),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1545),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1547),
.A2(n_1457),
.B(n_1517),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1430),
.A2(n_1517),
.B(n_1498),
.Y(n_1781)
);

AO31x2_ASAP7_75t_L g1782 ( 
.A1(n_1513),
.A2(n_1522),
.A3(n_1514),
.B(n_1431),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1426),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1417),
.B(n_1431),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_SL g1785 ( 
.A(n_1547),
.B(n_1457),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1417),
.A2(n_1431),
.B1(n_1501),
.B2(n_1502),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1502),
.A2(n_1501),
.B1(n_1431),
.B2(n_1417),
.C(n_1539),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1502),
.A2(n_1553),
.B1(n_1504),
.B2(n_1562),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1514),
.A2(n_1522),
.B1(n_1469),
.B2(n_1504),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1469),
.A2(n_1587),
.B1(n_1588),
.B2(n_1590),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1587),
.B(n_1447),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1588),
.A2(n_1590),
.B1(n_1562),
.B2(n_1574),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1733),
.B(n_1410),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1677),
.A2(n_1553),
.B1(n_1574),
.B2(n_1519),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1659),
.A2(n_1410),
.B1(n_1447),
.B2(n_1523),
.C(n_1433),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1603),
.A2(n_1519),
.B1(n_1523),
.B2(n_1511),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1688),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1684),
.A2(n_1498),
.B(n_1480),
.C(n_1454),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1656),
.A2(n_1480),
.B1(n_1472),
.B2(n_1479),
.C(n_1492),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1603),
.A2(n_1511),
.B1(n_1530),
.B2(n_1439),
.Y(n_1800)
);

BUFx12f_ASAP7_75t_L g1801 ( 
.A(n_1629),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1708),
.A2(n_1530),
.B1(n_1439),
.B2(n_1495),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1755),
.A2(n_1479),
.B1(n_1472),
.B2(n_1495),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1593),
.A2(n_1496),
.B1(n_1492),
.B2(n_1433),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1592),
.A2(n_1602),
.B1(n_1615),
.B2(n_1688),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1595),
.Y(n_1806)
);

OAI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1660),
.A2(n_1454),
.B(n_1462),
.C(n_1496),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1615),
.A2(n_1462),
.B(n_1430),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1731),
.A2(n_1409),
.B(n_1463),
.C(n_1429),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1755),
.A2(n_1463),
.B1(n_1409),
.B2(n_1429),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1597),
.A2(n_1415),
.B1(n_1527),
.B2(n_1717),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1607),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1638),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1622),
.A2(n_1527),
.B1(n_1742),
.B2(n_1686),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1701),
.A2(n_1680),
.B1(n_1703),
.B2(n_1664),
.C(n_1685),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1658),
.A2(n_1692),
.B1(n_1721),
.B2(n_1608),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_SL g1817 ( 
.A1(n_1597),
.A2(n_1748),
.B1(n_1669),
.B2(n_1672),
.Y(n_1817)
);

OAI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1599),
.A2(n_1623),
.B(n_1605),
.C(n_1687),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1711),
.A2(n_1751),
.B1(n_1741),
.B2(n_1596),
.C(n_1654),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1747),
.B(n_1745),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1749),
.A2(n_1762),
.B1(n_1738),
.B2(n_1642),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1728),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1625),
.A2(n_1669),
.B1(n_1672),
.B2(n_1626),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1620),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1693),
.B(n_1694),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1635),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1669),
.A2(n_1672),
.B1(n_1689),
.B2(n_1695),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1611),
.A2(n_1753),
.B1(n_1739),
.B2(n_1746),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1595),
.Y(n_1830)
);

AO21x2_ASAP7_75t_L g1831 ( 
.A1(n_1788),
.A2(n_1757),
.B(n_1780),
.Y(n_1831)
);

OAI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1634),
.A2(n_1729),
.B1(n_1727),
.B2(n_1712),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1661),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1749),
.A2(n_1627),
.B1(n_1727),
.B2(n_1640),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1663),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1729),
.A2(n_1634),
.B1(n_1720),
.B2(n_1704),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1635),
.Y(n_1837)
);

AOI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1591),
.A2(n_1616),
.B(n_1705),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1694),
.A2(n_1726),
.B1(n_1732),
.B2(n_1609),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1609),
.B(n_1724),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1718),
.A2(n_1629),
.B1(n_1640),
.B2(n_1705),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1676),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1646),
.B(n_1645),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1744),
.B(n_1618),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1772),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1724),
.B(n_1650),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1633),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1627),
.A2(n_1683),
.B1(n_1737),
.B2(n_1760),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1710),
.A2(n_1651),
.B1(n_1670),
.B2(n_1668),
.Y(n_1849)
);

AOI222xp33_ASAP7_75t_L g1850 ( 
.A1(n_1631),
.A2(n_1646),
.B1(n_1645),
.B2(n_1706),
.C1(n_1773),
.C2(n_1747),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1651),
.A2(n_1668),
.B1(n_1670),
.B2(n_1719),
.Y(n_1851)
);

AO31x2_ASAP7_75t_L g1852 ( 
.A1(n_1740),
.A2(n_1786),
.A3(n_1785),
.B(n_1789),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1651),
.A2(n_1725),
.B1(n_1647),
.B2(n_1773),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1614),
.A2(n_1621),
.B1(n_1744),
.B2(n_1750),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1683),
.A2(n_1676),
.B1(n_1617),
.B2(n_1614),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1733),
.B(n_1702),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1641),
.Y(n_1857)
);

OAI211xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1759),
.A2(n_1653),
.B(n_1758),
.C(n_1770),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1733),
.B(n_1633),
.Y(n_1859)
);

OAI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1687),
.A2(n_1792),
.B(n_1790),
.C(n_1777),
.Y(n_1860)
);

AO21x2_ASAP7_75t_L g1861 ( 
.A1(n_1600),
.A2(n_1632),
.B(n_1768),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1700),
.B(n_1707),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1771),
.A2(n_1673),
.B1(n_1617),
.B2(n_1734),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1644),
.A2(n_1613),
.B1(n_1754),
.B2(n_1775),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1621),
.A2(n_1697),
.B1(n_1690),
.B2(n_1679),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1740),
.A2(n_1787),
.B1(n_1778),
.B2(n_1637),
.C(n_1671),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1734),
.A2(n_1666),
.B1(n_1702),
.B2(n_1754),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1700),
.B(n_1707),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1613),
.A2(n_1783),
.B(n_1791),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1641),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1756),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1766),
.A2(n_1644),
.B1(n_1620),
.B2(n_1649),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1652),
.A2(n_1678),
.B1(n_1657),
.B2(n_1667),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1765),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1620),
.A2(n_1628),
.B1(n_1630),
.B2(n_1649),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1657),
.B(n_1667),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1772),
.A2(n_1730),
.B1(n_1649),
.B2(n_1630),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1652),
.A2(n_1678),
.B1(n_1674),
.B2(n_1696),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1673),
.A2(n_1766),
.B1(n_1630),
.B2(n_1628),
.Y(n_1879)
);

NOR2x1_ASAP7_75t_L g1880 ( 
.A(n_1628),
.B(n_1709),
.Y(n_1880)
);

AOI222xp33_ASAP7_75t_L g1881 ( 
.A1(n_1652),
.A2(n_1655),
.B1(n_1674),
.B2(n_1696),
.C1(n_1681),
.C2(n_1699),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1675),
.B(n_1699),
.Y(n_1882)
);

AO21x2_ASAP7_75t_L g1883 ( 
.A1(n_1761),
.A2(n_1781),
.B(n_1643),
.Y(n_1883)
);

OAI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1604),
.A2(n_1636),
.B(n_1698),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1604),
.A2(n_1636),
.B(n_1681),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1743),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1772),
.A2(n_1730),
.B1(n_1673),
.B2(n_1662),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1743),
.Y(n_1888)
);

OAI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1781),
.A2(n_1643),
.B(n_1598),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1662),
.A2(n_1665),
.B1(n_1764),
.B2(n_1736),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1594),
.A2(n_1624),
.B1(n_1619),
.B2(n_1612),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1601),
.B(n_1714),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1601),
.B(n_1714),
.Y(n_1893)
);

NOR3xp33_ASAP7_75t_L g1894 ( 
.A(n_1709),
.B(n_1716),
.C(n_1774),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1730),
.A2(n_1784),
.B(n_1598),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1610),
.A2(n_1662),
.B1(n_1779),
.B2(n_1774),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1655),
.A2(n_1698),
.B1(n_1610),
.B2(n_1736),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1662),
.A2(n_1665),
.B1(n_1767),
.B2(n_1764),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1767),
.A2(n_1776),
.B1(n_1709),
.B2(n_1716),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1774),
.A2(n_1776),
.B1(n_1716),
.B2(n_1610),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1648),
.B(n_1682),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1715),
.A2(n_1735),
.B1(n_1779),
.B2(n_1769),
.Y(n_1902)
);

AOI222xp33_ASAP7_75t_L g1903 ( 
.A1(n_1722),
.A2(n_1723),
.B1(n_1752),
.B2(n_1769),
.C1(n_1715),
.C2(n_1735),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1730),
.A2(n_1648),
.B1(n_1682),
.B2(n_1779),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1648),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1648),
.A2(n_1682),
.B1(n_1784),
.B2(n_1763),
.Y(n_1906)
);

OAI33xp33_ASAP7_75t_L g1907 ( 
.A1(n_1782),
.A2(n_1763),
.A3(n_1722),
.B1(n_1723),
.B2(n_1752),
.B3(n_1713),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1606),
.A2(n_1763),
.B(n_1723),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1722),
.A2(n_1723),
.B(n_1752),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1648),
.A2(n_1682),
.B1(n_1713),
.B2(n_1606),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1682),
.A2(n_1713),
.B1(n_1722),
.B2(n_1752),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1782),
.A2(n_1656),
.B1(n_1755),
.B2(n_1684),
.Y(n_1912)
);

AND2x6_ASAP7_75t_L g1913 ( 
.A(n_1782),
.B(n_1772),
.Y(n_1913)
);

AOI21xp33_ASAP7_75t_L g1914 ( 
.A1(n_1782),
.A2(n_885),
.B(n_784),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1782),
.A2(n_789),
.B1(n_796),
.B2(n_1275),
.C(n_747),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1744),
.B(n_1609),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1744),
.B(n_1609),
.Y(n_1917)
);

AO21x2_ASAP7_75t_L g1918 ( 
.A1(n_1788),
.A2(n_1448),
.B(n_1741),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1615),
.A2(n_1050),
.B(n_1741),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1920)
);

OAI211xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1684),
.A2(n_1116),
.B(n_877),
.C(n_1476),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1615),
.A2(n_1050),
.B(n_1741),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1656),
.A2(n_1755),
.B1(n_1684),
.B2(n_877),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1747),
.B(n_1449),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1603),
.A2(n_877),
.B1(n_1414),
.B2(n_1154),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1677),
.A2(n_921),
.B1(n_885),
.B2(n_1451),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1611),
.Y(n_1928)
);

OAI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1677),
.A2(n_1414),
.B1(n_1393),
.B2(n_1252),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1677),
.A2(n_789),
.B1(n_796),
.B2(n_1275),
.C(n_747),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1744),
.B(n_1609),
.Y(n_1931)
);

NAND2x1_ASAP7_75t_L g1932 ( 
.A(n_1601),
.B(n_1436),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1747),
.B(n_1449),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1677),
.A2(n_877),
.B1(n_747),
.B2(n_784),
.C(n_885),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1656),
.A2(n_1755),
.B1(n_1684),
.B2(n_877),
.Y(n_1935)
);

OAI211xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1684),
.A2(n_1116),
.B(n_877),
.C(n_1476),
.Y(n_1936)
);

AOI222xp33_ASAP7_75t_L g1937 ( 
.A1(n_1684),
.A2(n_1258),
.B1(n_1201),
.B2(n_789),
.C1(n_1237),
.C2(n_1241),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1677),
.A2(n_877),
.B1(n_747),
.B2(n_784),
.C(n_885),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1595),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1656),
.A2(n_885),
.B1(n_877),
.B2(n_796),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1656),
.A2(n_885),
.B1(n_877),
.B2(n_796),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1639),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1733),
.B(n_1772),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1607),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1656),
.A2(n_1755),
.B1(n_1684),
.B2(n_877),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1677),
.A2(n_789),
.B1(n_796),
.B2(n_1275),
.C(n_747),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1677),
.A2(n_789),
.B1(n_796),
.B2(n_1275),
.C(n_747),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1656),
.A2(n_1755),
.B1(n_1684),
.B2(n_877),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1949)
);

AOI321xp33_ASAP7_75t_L g1950 ( 
.A1(n_1677),
.A2(n_789),
.A3(n_1684),
.B1(n_1659),
.B2(n_1664),
.C(n_1660),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1656),
.A2(n_1755),
.B1(n_1684),
.B2(n_877),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_SL g1952 ( 
.A1(n_1677),
.A2(n_921),
.B1(n_885),
.B2(n_1451),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1677),
.A2(n_789),
.B1(n_796),
.B2(n_1275),
.C(n_747),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1956)
);

OAI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1684),
.A2(n_1289),
.B(n_877),
.C(n_983),
.Y(n_1957)
);

NAND2xp33_ASAP7_75t_R g1958 ( 
.A(n_1599),
.B(n_1179),
.Y(n_1958)
);

AOI322xp5_ASAP7_75t_L g1959 ( 
.A1(n_1684),
.A2(n_1289),
.A3(n_983),
.B1(n_942),
.B2(n_1659),
.C1(n_1664),
.C2(n_1660),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1960)
);

BUFx10_ASAP7_75t_L g1961 ( 
.A(n_1627),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1889),
.A2(n_1808),
.B(n_1895),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1871),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1847),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1821),
.B(n_1870),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1843),
.B(n_1840),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1908),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1843),
.B(n_1918),
.Y(n_1968)
);

NOR2x1_ASAP7_75t_L g1969 ( 
.A(n_1832),
.B(n_1875),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1874),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1852),
.B(n_1918),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1913),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1852),
.B(n_1916),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1847),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1844),
.B(n_1917),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1939),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1931),
.B(n_1812),
.Y(n_1977)
);

OR2x2_ASAP7_75t_SL g1978 ( 
.A(n_1823),
.B(n_1856),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1908),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1913),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1942),
.B(n_1906),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1813),
.Y(n_1982)
);

CKINVDCx11_ASAP7_75t_R g1983 ( 
.A(n_1842),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1852),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1906),
.B(n_1845),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1852),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1913),
.B(n_1909),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1833),
.B(n_1835),
.Y(n_1988)
);

INVxp67_ASAP7_75t_L g1989 ( 
.A(n_1846),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1939),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1827),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1827),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1909),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1913),
.B(n_1831),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1831),
.B(n_1793),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1837),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1793),
.Y(n_1997)
);

AO21x2_ASAP7_75t_L g1998 ( 
.A1(n_1919),
.A2(n_1922),
.B(n_1914),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1846),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1793),
.B(n_1866),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1883),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1882),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1944),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1889),
.Y(n_2004)
);

AND2x4_ASAP7_75t_SL g2005 ( 
.A(n_1943),
.B(n_1892),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1876),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1904),
.B(n_1861),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1861),
.B(n_1883),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1857),
.B(n_1885),
.Y(n_2009)
);

BUFx6f_ASAP7_75t_L g2010 ( 
.A(n_1892),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1869),
.B(n_1836),
.Y(n_2011)
);

OAI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1930),
.A2(n_1955),
.B1(n_1947),
.B2(n_1946),
.C(n_1934),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1884),
.Y(n_2013)
);

AO21x2_ASAP7_75t_L g2014 ( 
.A1(n_1804),
.A2(n_1860),
.B(n_1838),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1800),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1902),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1829),
.B(n_1867),
.Y(n_2017)
);

OAI222xp33_ASAP7_75t_L g2018 ( 
.A1(n_1912),
.A2(n_1820),
.B1(n_1923),
.B2(n_1945),
.C1(n_1951),
.C2(n_1948),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1796),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1839),
.B(n_1924),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1893),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1902),
.Y(n_2022)
);

INVxp67_ASAP7_75t_SL g2023 ( 
.A(n_1809),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1943),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1887),
.B(n_1877),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1943),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1896),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1839),
.B(n_1933),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1897),
.B(n_1810),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1915),
.B(n_1940),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1858),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1891),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1897),
.B(n_1864),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1881),
.B(n_1853),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1891),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1853),
.B(n_1819),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1905),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1826),
.B(n_1920),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1926),
.B(n_1949),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1953),
.B(n_1954),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1829),
.B(n_1867),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1956),
.B(n_1960),
.Y(n_2042)
);

AND2x4_ASAP7_75t_SL g2043 ( 
.A(n_1825),
.B(n_1872),
.Y(n_2043)
);

INVx4_ASAP7_75t_L g2044 ( 
.A(n_1825),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_1802),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1794),
.A2(n_1807),
.B(n_1798),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1903),
.B(n_1803),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1901),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1803),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1850),
.B(n_1824),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2003),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2003),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1963),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2012),
.A2(n_1941),
.B1(n_1952),
.B2(n_1927),
.C(n_1951),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1964),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_R g2056 ( 
.A(n_1983),
.B(n_1842),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2012),
.A2(n_1923),
.B1(n_1948),
.B2(n_1945),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1991),
.Y(n_2058)
);

OAI33xp33_ASAP7_75t_L g2059 ( 
.A1(n_2031),
.A2(n_1929),
.A3(n_1925),
.B1(n_1936),
.B2(n_1921),
.B3(n_1928),
.Y(n_2059)
);

AOI221xp5_ASAP7_75t_L g2060 ( 
.A1(n_2018),
.A2(n_1938),
.B1(n_1935),
.B2(n_1957),
.C(n_1912),
.Y(n_2060)
);

OAI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2030),
.A2(n_1935),
.B1(n_1950),
.B2(n_1958),
.C(n_1937),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1989),
.B(n_1797),
.Y(n_2062)
);

OA21x2_ASAP7_75t_L g2063 ( 
.A1(n_1962),
.A2(n_1795),
.B(n_1810),
.Y(n_2063)
);

NAND3xp33_ASAP7_75t_L g2064 ( 
.A(n_2030),
.B(n_1958),
.C(n_1959),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1983),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1991),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1968),
.B(n_1966),
.Y(n_2067)
);

INVx2_ASAP7_75t_SL g2068 ( 
.A(n_2005),
.Y(n_2068)
);

AOI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2018),
.A2(n_1818),
.B1(n_1805),
.B2(n_1815),
.C(n_1848),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1962),
.A2(n_1799),
.B(n_1814),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2031),
.A2(n_1816),
.B1(n_1865),
.B2(n_1824),
.C(n_1828),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_1998),
.A2(n_1900),
.B(n_1863),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_L g2073 ( 
.A(n_2014),
.B(n_1969),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2050),
.A2(n_1817),
.B1(n_1816),
.B2(n_1822),
.Y(n_2074)
);

NAND4xp25_ASAP7_75t_SL g2075 ( 
.A(n_2050),
.B(n_1841),
.C(n_1854),
.D(n_1849),
.Y(n_2075)
);

NOR3xp33_ASAP7_75t_L g2076 ( 
.A(n_2023),
.B(n_1879),
.C(n_1855),
.Y(n_2076)
);

AND2x6_ASAP7_75t_SL g2077 ( 
.A(n_2025),
.B(n_1801),
.Y(n_2077)
);

OAI221xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2023),
.A2(n_1828),
.B1(n_1849),
.B2(n_1854),
.C(n_1851),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1992),
.Y(n_2079)
);

AO21x2_ASAP7_75t_L g2080 ( 
.A1(n_1998),
.A2(n_1894),
.B(n_1899),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1963),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_SL g2082 ( 
.A1(n_2011),
.A2(n_1932),
.B1(n_1898),
.B2(n_1890),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1989),
.B(n_1865),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1992),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2017),
.A2(n_1851),
.B1(n_1878),
.B2(n_1873),
.Y(n_2085)
);

OR2x2_ASAP7_75t_SL g2086 ( 
.A(n_2011),
.B(n_1905),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1970),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1968),
.B(n_1873),
.Y(n_2088)
);

OAI211xp5_ASAP7_75t_L g2089 ( 
.A1(n_2017),
.A2(n_1878),
.B(n_1811),
.C(n_1910),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1970),
.Y(n_2090)
);

NAND3xp33_ASAP7_75t_L g2091 ( 
.A(n_2013),
.B(n_1880),
.C(n_1806),
.Y(n_2091)
);

OAI322xp33_ASAP7_75t_L g2092 ( 
.A1(n_2041),
.A2(n_1834),
.A3(n_1886),
.B1(n_1806),
.B2(n_1830),
.C1(n_1888),
.C2(n_1862),
.Y(n_2092)
);

AOI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_2049),
.A2(n_1907),
.B1(n_1859),
.B2(n_1830),
.C(n_1868),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1982),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1999),
.B(n_1911),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1982),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1997),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1992),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1999),
.B(n_1825),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2034),
.A2(n_1801),
.B1(n_1888),
.B2(n_1961),
.Y(n_2100)
);

AOI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_2049),
.A2(n_1961),
.B1(n_2041),
.B2(n_2013),
.C(n_2019),
.Y(n_2101)
);

AOI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2019),
.A2(n_1961),
.B1(n_2015),
.B2(n_2034),
.C(n_2033),
.Y(n_2102)
);

OAI221xp5_ASAP7_75t_L g2103 ( 
.A1(n_1969),
.A2(n_2011),
.B1(n_2015),
.B2(n_2045),
.C(n_2033),
.Y(n_2103)
);

AO21x2_ASAP7_75t_L g2104 ( 
.A1(n_1998),
.A2(n_1962),
.B(n_2046),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_2034),
.A2(n_2033),
.B1(n_2045),
.B2(n_2029),
.C(n_2014),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1968),
.B(n_1966),
.Y(n_2106)
);

OA21x2_ASAP7_75t_L g2107 ( 
.A1(n_2001),
.A2(n_2008),
.B(n_1971),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_2004),
.A2(n_2008),
.B(n_1971),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1975),
.B(n_2038),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1965),
.B(n_1975),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_1973),
.B(n_1978),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1966),
.B(n_2024),
.Y(n_2112)
);

NAND4xp25_ASAP7_75t_L g2113 ( 
.A(n_2000),
.B(n_2022),
.C(n_2016),
.D(n_2032),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_2010),
.Y(n_2114)
);

NAND3xp33_ASAP7_75t_L g2115 ( 
.A(n_2032),
.B(n_2035),
.C(n_2016),
.Y(n_2115)
);

AOI31xp33_ASAP7_75t_L g2116 ( 
.A1(n_2025),
.A2(n_2036),
.A3(n_2000),
.B(n_2047),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2014),
.A2(n_2047),
.B1(n_2025),
.B2(n_2036),
.Y(n_2117)
);

OAI211xp5_ASAP7_75t_L g2118 ( 
.A1(n_2047),
.A2(n_2007),
.B(n_2000),
.C(n_2027),
.Y(n_2118)
);

HB1xp67_ASAP7_75t_L g2119 ( 
.A(n_2009),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1964),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1996),
.Y(n_2121)
);

OAI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_2020),
.A2(n_2028),
.B1(n_2027),
.B2(n_1972),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2009),
.Y(n_2123)
);

NOR4xp25_ASAP7_75t_SL g2124 ( 
.A(n_1980),
.B(n_2027),
.C(n_1972),
.D(n_2001),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_SL g2125 ( 
.A1(n_1971),
.A2(n_2007),
.B1(n_2020),
.B2(n_2028),
.C(n_2036),
.Y(n_2125)
);

NOR4xp25_ASAP7_75t_SL g2126 ( 
.A(n_1980),
.B(n_2001),
.C(n_2026),
.D(n_2035),
.Y(n_2126)
);

NAND3xp33_ASAP7_75t_L g2127 ( 
.A(n_2022),
.B(n_1984),
.C(n_1986),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_2010),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_2014),
.A2(n_2029),
.B1(n_1998),
.B2(n_2046),
.Y(n_2129)
);

NOR2xp67_ASAP7_75t_L g2130 ( 
.A(n_2118),
.B(n_1997),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2119),
.B(n_1973),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2058),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2053),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2067),
.B(n_1995),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2067),
.B(n_1995),
.Y(n_2135)
);

NAND4xp25_ASAP7_75t_L g2136 ( 
.A(n_2064),
.B(n_2007),
.C(n_2029),
.D(n_2028),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2106),
.B(n_1995),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2123),
.B(n_2009),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2111),
.B(n_1973),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2051),
.B(n_2048),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2051),
.B(n_2048),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2066),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2053),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2081),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2081),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2066),
.Y(n_2146)
);

NAND5xp2_ASAP7_75t_L g2147 ( 
.A(n_2069),
.B(n_1987),
.C(n_1994),
.D(n_1980),
.E(n_2014),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_2097),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2052),
.B(n_2006),
.Y(n_2149)
);

OR2x6_ASAP7_75t_L g2150 ( 
.A(n_2073),
.B(n_1987),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2086),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2111),
.B(n_1978),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2106),
.B(n_1978),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2114),
.B(n_1967),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2112),
.B(n_1994),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2112),
.B(n_1994),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2052),
.B(n_2006),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2087),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2087),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2090),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2097),
.B(n_1985),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2090),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2110),
.B(n_2002),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_2055),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2065),
.B(n_2038),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2117),
.B(n_2109),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2088),
.B(n_1985),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2079),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2088),
.B(n_1985),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2107),
.B(n_1984),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2114),
.B(n_1987),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2114),
.B(n_1997),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2128),
.B(n_1997),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2094),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2079),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_2128),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2094),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2084),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2107),
.B(n_1986),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_2073),
.B(n_1993),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2128),
.B(n_1997),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_2108),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2108),
.B(n_2029),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2096),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2117),
.B(n_2002),
.Y(n_2185)
);

AND2x4_ASAP7_75t_SL g2186 ( 
.A(n_2068),
.B(n_2044),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2086),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2107),
.B(n_2029),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2098),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2098),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2121),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2107),
.B(n_1981),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2129),
.B(n_1981),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2068),
.B(n_1967),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_2125),
.B(n_2008),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2139),
.B(n_2127),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2130),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2133),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_SL g2200 ( 
.A(n_2130),
.B(n_2065),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2166),
.B(n_2105),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2151),
.B(n_2124),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2133),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2143),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2166),
.B(n_2116),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2163),
.B(n_2167),
.Y(n_2206)
);

NAND2xp33_ASAP7_75t_SL g2207 ( 
.A(n_2151),
.B(n_2056),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2143),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2187),
.B(n_2167),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2187),
.B(n_2072),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2139),
.B(n_2115),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_2185),
.Y(n_2212)
);

INVxp67_ASAP7_75t_SL g2213 ( 
.A(n_2152),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2170),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2163),
.B(n_2101),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2144),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2144),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2167),
.B(n_2072),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2169),
.B(n_2072),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2170),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2169),
.B(n_2024),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2165),
.B(n_2100),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2185),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2131),
.B(n_2122),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2136),
.A2(n_2103),
.B(n_2061),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2145),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_2164),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2145),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2158),
.Y(n_2229)
);

INVxp67_ASAP7_75t_L g2230 ( 
.A(n_2149),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_2154),
.B(n_1993),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2169),
.B(n_2024),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2131),
.B(n_2083),
.Y(n_2233)
);

NAND2x1_ASAP7_75t_SL g2234 ( 
.A(n_2188),
.B(n_2100),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2136),
.B(n_2102),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2195),
.B(n_2113),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2147),
.B(n_2054),
.C(n_2057),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_2154),
.B(n_1993),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2147),
.A2(n_2060),
.B1(n_2075),
.B2(n_2076),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2170),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2149),
.B(n_2157),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2195),
.B(n_2121),
.Y(n_2242)
);

NOR2xp67_ASAP7_75t_L g2243 ( 
.A(n_2152),
.B(n_2091),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2179),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2157),
.B(n_2062),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2193),
.B(n_2093),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2158),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2159),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2179),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2215),
.B(n_2201),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2199),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2214),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2211),
.B(n_2195),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2209),
.Y(n_2254)
);

OAI31xp33_ASAP7_75t_L g2255 ( 
.A1(n_2207),
.A2(n_2193),
.A3(n_2089),
.B(n_2078),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2235),
.B(n_2212),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2227),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2199),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2211),
.B(n_2138),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2203),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2223),
.B(n_2193),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2203),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2204),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_SL g2264 ( 
.A1(n_2225),
.A2(n_2085),
.B1(n_2188),
.B2(n_2082),
.Y(n_2264)
);

NAND2x1_ASAP7_75t_SL g2265 ( 
.A(n_2197),
.B(n_2188),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2204),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2205),
.B(n_2161),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2208),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2208),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2196),
.B(n_2138),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2234),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2214),
.Y(n_2272)
);

NAND2x1p5_ASAP7_75t_L g2273 ( 
.A(n_2243),
.B(n_2164),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2216),
.Y(n_2274)
);

NAND2xp33_ASAP7_75t_SL g2275 ( 
.A(n_2234),
.B(n_2126),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_SL g2276 ( 
.A(n_2239),
.B(n_2077),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2230),
.B(n_2161),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2214),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2196),
.B(n_2153),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2237),
.A2(n_2070),
.B(n_2074),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2216),
.Y(n_2281)
);

NAND3x1_ASAP7_75t_SL g2282 ( 
.A(n_2202),
.B(n_2071),
.C(n_2077),
.Y(n_2282)
);

NAND2xp33_ASAP7_75t_SL g2283 ( 
.A(n_2236),
.B(n_2153),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2246),
.B(n_2161),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2220),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2217),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2198),
.Y(n_2287)
);

NOR4xp25_ASAP7_75t_SL g2288 ( 
.A(n_2213),
.B(n_2026),
.C(n_2177),
.D(n_2162),
.Y(n_2288)
);

AOI221xp5_ASAP7_75t_SL g2289 ( 
.A1(n_2236),
.A2(n_2192),
.B1(n_2183),
.B2(n_2092),
.C(n_2082),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2217),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2245),
.B(n_2155),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2242),
.B(n_2150),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_SL g2293 ( 
.A(n_2200),
.B(n_2092),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2241),
.B(n_2155),
.Y(n_2294)
);

NOR2xp67_ASAP7_75t_L g2295 ( 
.A(n_2243),
.B(n_2148),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2209),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2226),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2220),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2222),
.B(n_2206),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2221),
.B(n_2155),
.Y(n_2300)
);

INVx1_ASAP7_75t_SL g2301 ( 
.A(n_2257),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2251),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2258),
.Y(n_2303)
);

OAI321xp33_ASAP7_75t_L g2304 ( 
.A1(n_2273),
.A2(n_2202),
.A3(n_2210),
.B1(n_2218),
.B2(n_2219),
.C(n_2150),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2299),
.B(n_2210),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2260),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_2250),
.B(n_2233),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2276),
.A2(n_2293),
.B1(n_2264),
.B2(n_2289),
.Y(n_2308)
);

AOI211xp5_ASAP7_75t_L g2309 ( 
.A1(n_2276),
.A2(n_2218),
.B(n_2219),
.C(n_2059),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2253),
.B(n_2233),
.Y(n_2310)
);

AOI322xp5_ASAP7_75t_L g2311 ( 
.A1(n_2256),
.A2(n_2299),
.A3(n_2283),
.B1(n_2275),
.B2(n_2284),
.C1(n_2261),
.C2(n_2192),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_2280),
.A2(n_2070),
.B(n_2150),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2273),
.B(n_2192),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2262),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2263),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2266),
.Y(n_2316)
);

AOI21x1_ASAP7_75t_SL g2317 ( 
.A1(n_2267),
.A2(n_2154),
.B(n_2194),
.Y(n_2317)
);

AOI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2283),
.A2(n_2183),
.B1(n_2182),
.B2(n_2240),
.C(n_2249),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2271),
.B(n_2231),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2255),
.B(n_2221),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2296),
.B(n_2232),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2254),
.B(n_2232),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2271),
.B(n_2224),
.Y(n_2323)
);

OAI322xp33_ASAP7_75t_L g2324 ( 
.A1(n_2253),
.A2(n_2242),
.A3(n_2224),
.B1(n_2179),
.B2(n_2249),
.C1(n_2240),
.C2(n_2220),
.Y(n_2324)
);

OAI332xp33_ASAP7_75t_L g2325 ( 
.A1(n_2279),
.A2(n_2249),
.A3(n_2240),
.B1(n_2244),
.B2(n_2095),
.B3(n_2148),
.C1(n_2226),
.C2(n_2248),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2279),
.B(n_2038),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2275),
.A2(n_2150),
.B1(n_2180),
.B2(n_2198),
.C(n_2183),
.Y(n_2327)
);

AOI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2295),
.A2(n_2150),
.B(n_2180),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2270),
.B(n_2244),
.Y(n_2329)
);

NOR4xp25_ASAP7_75t_L g2330 ( 
.A(n_2282),
.B(n_2198),
.C(n_2244),
.D(n_2247),
.Y(n_2330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2331 ( 
.A1(n_2282),
.A2(n_2248),
.B(n_2247),
.C(n_2228),
.D(n_2229),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2277),
.B(n_2039),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2288),
.A2(n_2150),
.B1(n_2180),
.B2(n_2020),
.Y(n_2333)
);

AOI221xp5_ASAP7_75t_SL g2334 ( 
.A1(n_2292),
.A2(n_2182),
.B1(n_2229),
.B2(n_2228),
.C(n_2198),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2270),
.A2(n_2080),
.B1(n_2046),
.B2(n_1998),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2268),
.Y(n_2336)
);

AOI221x1_ASAP7_75t_L g2337 ( 
.A1(n_2287),
.A2(n_2141),
.B1(n_2140),
.B2(n_2099),
.C(n_2177),
.Y(n_2337)
);

OA21x2_ASAP7_75t_L g2338 ( 
.A1(n_2265),
.A2(n_2238),
.B(n_2231),
.Y(n_2338)
);

OAI21xp33_ASAP7_75t_L g2339 ( 
.A1(n_2265),
.A2(n_2180),
.B(n_1977),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2291),
.B(n_2039),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2269),
.Y(n_2341)
);

NAND2x1_ASAP7_75t_L g2342 ( 
.A(n_2338),
.B(n_2287),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2301),
.Y(n_2343)
);

OAI21xp33_ASAP7_75t_L g2344 ( 
.A1(n_2308),
.A2(n_2259),
.B(n_2292),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2302),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2307),
.B(n_2259),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2303),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2325),
.B(n_2294),
.Y(n_2348)
);

OAI33xp33_ASAP7_75t_L g2349 ( 
.A1(n_2333),
.A2(n_2281),
.A3(n_2274),
.B1(n_2286),
.B2(n_2297),
.B3(n_2290),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2307),
.B(n_2300),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2310),
.B(n_2252),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_L g2352 ( 
.A(n_2320),
.B(n_2287),
.Y(n_2352)
);

A2O1A1Ixp33_ASAP7_75t_L g2353 ( 
.A1(n_2311),
.A2(n_2182),
.B(n_2164),
.C(n_2043),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2306),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2314),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2338),
.Y(n_2356)
);

AOI21xp33_ASAP7_75t_L g2357 ( 
.A1(n_2323),
.A2(n_2312),
.B(n_2304),
.Y(n_2357)
);

NAND2xp33_ASAP7_75t_SL g2358 ( 
.A(n_2331),
.B(n_2148),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2323),
.B(n_2039),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2319),
.B(n_2313),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2309),
.B(n_2040),
.Y(n_2361)
);

NAND3xp33_ASAP7_75t_SL g2362 ( 
.A(n_2330),
.B(n_2298),
.C(n_2285),
.Y(n_2362)
);

AOI221xp5_ASAP7_75t_L g2363 ( 
.A1(n_2324),
.A2(n_2182),
.B1(n_2278),
.B2(n_2272),
.C(n_2298),
.Y(n_2363)
);

NOR2x1_ASAP7_75t_L g2364 ( 
.A(n_2310),
.B(n_2252),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2327),
.B(n_2285),
.C(n_2278),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2315),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2316),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2326),
.B(n_2272),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2336),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2338),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2341),
.Y(n_2371)
);

OAI22xp33_ASAP7_75t_L g2372 ( 
.A1(n_2305),
.A2(n_2180),
.B1(n_2182),
.B2(n_2063),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2364),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_2343),
.B(n_2339),
.Y(n_2374)
);

INVxp67_ASAP7_75t_L g2375 ( 
.A(n_2352),
.Y(n_2375)
);

OR2x2_ASAP7_75t_L g2376 ( 
.A(n_2361),
.B(n_2321),
.Y(n_2376)
);

AND3x1_ASAP7_75t_L g2377 ( 
.A(n_2353),
.B(n_2318),
.C(n_2313),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2360),
.B(n_2319),
.Y(n_2378)
);

AOI322xp5_ASAP7_75t_L g2379 ( 
.A1(n_2348),
.A2(n_2334),
.A3(n_2335),
.B1(n_2322),
.B2(n_2332),
.C1(n_2340),
.C2(n_2337),
.Y(n_2379)
);

NOR4xp25_ASAP7_75t_SL g2380 ( 
.A(n_2358),
.B(n_2337),
.C(n_2317),
.D(n_2328),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2348),
.B(n_2329),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2344),
.B(n_2329),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2358),
.B(n_2182),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2345),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2347),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2346),
.B(n_2040),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2354),
.Y(n_2387)
);

XNOR2xp5_ASAP7_75t_L g2388 ( 
.A(n_2350),
.B(n_2043),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2349),
.B(n_2140),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2342),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2362),
.A2(n_2104),
.B1(n_2180),
.B2(n_2046),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2359),
.B(n_2040),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2356),
.Y(n_2393)
);

OAI22xp33_ASAP7_75t_L g2394 ( 
.A1(n_2357),
.A2(n_2120),
.B1(n_2055),
.B2(n_1967),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2352),
.B(n_2141),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2355),
.Y(n_2396)
);

NOR2x1_ASAP7_75t_L g2397 ( 
.A(n_2356),
.B(n_2231),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2390),
.Y(n_2398)
);

OAI321xp33_ASAP7_75t_L g2399 ( 
.A1(n_2381),
.A2(n_2383),
.A3(n_2394),
.B1(n_2391),
.B2(n_2382),
.C(n_2353),
.Y(n_2399)
);

OAI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2383),
.A2(n_2370),
.B1(n_2363),
.B2(n_2372),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2393),
.B(n_2370),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2378),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2378),
.B(n_2366),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2377),
.B(n_2365),
.Y(n_2404)
);

OAI221xp5_ASAP7_75t_L g2405 ( 
.A1(n_2389),
.A2(n_2367),
.B1(n_2369),
.B2(n_2371),
.C(n_2351),
.Y(n_2405)
);

NOR4xp25_ASAP7_75t_L g2406 ( 
.A(n_2375),
.B(n_2372),
.C(n_2368),
.D(n_2176),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2374),
.B(n_2231),
.Y(n_2407)
);

AOI322xp5_ASAP7_75t_L g2408 ( 
.A1(n_2389),
.A2(n_2374),
.A3(n_2373),
.B1(n_2395),
.B2(n_2384),
.C1(n_2396),
.C2(n_2385),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2379),
.A2(n_2238),
.B(n_2194),
.Y(n_2409)
);

AND4x1_ASAP7_75t_L g2410 ( 
.A(n_2397),
.B(n_2171),
.C(n_2135),
.D(n_2137),
.Y(n_2410)
);

NOR4xp25_ASAP7_75t_L g2411 ( 
.A(n_2387),
.B(n_2390),
.C(n_2395),
.D(n_2376),
.Y(n_2411)
);

NAND4xp25_ASAP7_75t_L g2412 ( 
.A(n_2386),
.B(n_2194),
.C(n_2238),
.D(n_2120),
.Y(n_2412)
);

AOI211xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2399),
.A2(n_2380),
.B(n_2392),
.C(n_2388),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_L g2414 ( 
.A1(n_2411),
.A2(n_2104),
.B1(n_2046),
.B2(n_2238),
.C(n_2080),
.Y(n_2414)
);

O2A1O1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2404),
.A2(n_2104),
.B(n_2080),
.C(n_2176),
.Y(n_2415)
);

OAI211xp5_ASAP7_75t_L g2416 ( 
.A1(n_2408),
.A2(n_2063),
.B(n_2171),
.C(n_2176),
.Y(n_2416)
);

AOI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2400),
.A2(n_2194),
.B1(n_2159),
.B2(n_2160),
.C(n_2162),
.Y(n_2417)
);

OAI211xp5_ASAP7_75t_SL g2418 ( 
.A1(n_2405),
.A2(n_2160),
.B(n_2174),
.C(n_2184),
.Y(n_2418)
);

NOR3xp33_ASAP7_75t_L g2419 ( 
.A(n_2403),
.B(n_2044),
.C(n_1977),
.Y(n_2419)
);

NAND2xp33_ASAP7_75t_SL g2420 ( 
.A(n_2402),
.B(n_2042),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2400),
.B(n_2194),
.Y(n_2421)
);

AOI221xp5_ASAP7_75t_L g2422 ( 
.A1(n_2406),
.A2(n_2409),
.B1(n_2407),
.B2(n_2398),
.C(n_2412),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2401),
.A2(n_2186),
.B1(n_2154),
.B2(n_2171),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2410),
.A2(n_2186),
.B1(n_2154),
.B2(n_2043),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_2420),
.Y(n_2425)
);

AOI211xp5_ASAP7_75t_L g2426 ( 
.A1(n_2421),
.A2(n_2172),
.B(n_2173),
.C(n_2181),
.Y(n_2426)
);

NAND2xp33_ASAP7_75t_SL g2427 ( 
.A(n_2413),
.B(n_2042),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2422),
.Y(n_2428)
);

OAI322xp33_ASAP7_75t_L g2429 ( 
.A1(n_2423),
.A2(n_2174),
.A3(n_2184),
.B1(n_2135),
.B2(n_2134),
.C1(n_2137),
.C2(n_2156),
.Y(n_2429)
);

AOI222xp33_ASAP7_75t_L g2430 ( 
.A1(n_2417),
.A2(n_2042),
.B1(n_2135),
.B2(n_2134),
.C1(n_2137),
.C2(n_2156),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2419),
.B(n_2172),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2416),
.A2(n_2186),
.B1(n_2172),
.B2(n_2173),
.Y(n_2432)
);

NAND3xp33_ASAP7_75t_L g2433 ( 
.A(n_2428),
.B(n_2414),
.C(n_2418),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_R g2434 ( 
.A(n_2425),
.B(n_1964),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2427),
.Y(n_2435)
);

CKINVDCx20_ASAP7_75t_R g2436 ( 
.A(n_2432),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2426),
.B(n_2424),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2429),
.Y(n_2438)
);

OAI21xp33_ASAP7_75t_L g2439 ( 
.A1(n_2431),
.A2(n_2430),
.B(n_2415),
.Y(n_2439)
);

NAND4xp25_ASAP7_75t_L g2440 ( 
.A(n_2431),
.B(n_1976),
.C(n_1990),
.D(n_1974),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2434),
.Y(n_2441)
);

NOR4xp25_ASAP7_75t_L g2442 ( 
.A(n_2435),
.B(n_2134),
.C(n_2173),
.D(n_2181),
.Y(n_2442)
);

NOR3xp33_ASAP7_75t_L g2443 ( 
.A(n_2433),
.B(n_2439),
.C(n_2438),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2437),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_SL g2445 ( 
.A(n_2436),
.B(n_2044),
.C(n_2181),
.Y(n_2445)
);

OAI322xp33_ASAP7_75t_L g2446 ( 
.A1(n_2440),
.A2(n_2191),
.A3(n_2142),
.B1(n_2132),
.B2(n_2168),
.C1(n_2189),
.C2(n_2175),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2435),
.Y(n_2447)
);

NOR3xp33_ASAP7_75t_SL g2448 ( 
.A(n_2445),
.B(n_1965),
.C(n_1988),
.Y(n_2448)
);

AOI211xp5_ASAP7_75t_L g2449 ( 
.A1(n_2443),
.A2(n_2156),
.B(n_1967),
.C(n_1979),
.Y(n_2449)
);

CKINVDCx20_ASAP7_75t_R g2450 ( 
.A(n_2447),
.Y(n_2450)
);

OAI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2444),
.A2(n_2191),
.B1(n_2142),
.B2(n_2168),
.Y(n_2451)
);

HB1xp67_ASAP7_75t_L g2452 ( 
.A(n_2450),
.Y(n_2452)
);

OR5x1_ASAP7_75t_L g2453 ( 
.A(n_2449),
.B(n_2441),
.C(n_2442),
.D(n_2446),
.E(n_2037),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2452),
.A2(n_2448),
.B1(n_2451),
.B2(n_2453),
.Y(n_2454)
);

AOI221xp5_ASAP7_75t_L g2455 ( 
.A1(n_2452),
.A2(n_2191),
.B1(n_2142),
.B2(n_2132),
.C(n_2168),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2454),
.B(n_1974),
.Y(n_2456)
);

NAND3x2_ASAP7_75t_L g2457 ( 
.A(n_2455),
.B(n_2026),
.C(n_2021),
.Y(n_2457)
);

HB1xp67_ASAP7_75t_L g2458 ( 
.A(n_2454),
.Y(n_2458)
);

OA21x2_ASAP7_75t_L g2459 ( 
.A1(n_2458),
.A2(n_2175),
.B(n_2189),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2456),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2460),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2459),
.A2(n_2456),
.B1(n_2457),
.B2(n_1967),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2461),
.A2(n_2459),
.B1(n_2146),
.B2(n_2190),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2463),
.A2(n_2462),
.B1(n_2459),
.B2(n_2178),
.Y(n_2464)
);

AOI211xp5_ASAP7_75t_L g2465 ( 
.A1(n_2464),
.A2(n_1976),
.B(n_1990),
.C(n_1974),
.Y(n_2465)
);


endmodule