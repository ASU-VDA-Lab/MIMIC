module fake_jpeg_21429_n_261 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_1),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_24),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_48),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_23),
.B1(n_44),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_31),
.B1(n_17),
.B2(n_27),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_26),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_19),
.B1(n_25),
.B2(n_21),
.Y(n_59)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_45),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_69),
.B1(n_82),
.B2(n_100),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_44),
.B1(n_40),
.B2(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_70),
.B(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_101),
.B1(n_62),
.B2(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_44),
.B1(n_32),
.B2(n_29),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_41),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_67),
.B(n_22),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_16),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_89),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_30),
.B(n_34),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_65),
.C(n_41),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_2),
.B(n_3),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_2),
.B(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_16),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_36),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_83),
.B1(n_77),
.B2(n_100),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_109),
.B1(n_121),
.B2(n_127),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_61),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_119),
.B(n_122),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_34),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_117),
.Y(n_146)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_87),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_36),
.B1(n_28),
.B2(n_67),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_72),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_80),
.A3(n_70),
.B1(n_79),
.B2(n_84),
.C1(n_8),
.C2(n_9),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_143),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_140),
.Y(n_168)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_110),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_103),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_94),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_105),
.B1(n_119),
.B2(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_155),
.B1(n_106),
.B2(n_93),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_90),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_81),
.B1(n_90),
.B2(n_99),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_71),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_113),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_71),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_127),
.B(n_121),
.C(n_117),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_4),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_122),
.C(n_119),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_148),
.C(n_139),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_123),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_179),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_123),
.B1(n_122),
.B2(n_126),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_175),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_116),
.A3(n_126),
.B1(n_120),
.B2(n_102),
.C1(n_113),
.C2(n_22),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_120),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_135),
.B1(n_140),
.B2(n_97),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_131),
.B1(n_91),
.B2(n_28),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_4),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_98),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_191),
.C(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_162),
.B1(n_161),
.B2(n_158),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_139),
.C(n_133),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_150),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_198),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_137),
.C(n_86),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_150),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_91),
.C(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_198),
.C(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_5),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_213),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_177),
.A3(n_171),
.B1(n_173),
.B2(n_175),
.C(n_161),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_200),
.B(n_192),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_177),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_216),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_158),
.A3(n_161),
.B1(n_171),
.B2(n_164),
.C1(n_175),
.C2(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_163),
.B1(n_159),
.B2(n_7),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_159),
.B1(n_184),
.B2(n_7),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_200),
.B(n_182),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_229),
.B(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_201),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_202),
.B(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_220),
.B(n_218),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_229),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_187),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_210),
.B1(n_211),
.B2(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_5),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_211),
.B1(n_203),
.B2(n_7),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_234),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_15),
.B1(n_6),
.B2(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_222),
.B(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_227),
.C(n_8),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_237),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_239),
.B(n_235),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_249),
.B(n_250),
.Y(n_252)
);

AOI31xp33_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_231),
.A3(n_234),
.B(n_10),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_244),
.C(n_245),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_242),
.B(n_241),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_6),
.C(n_9),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_10),
.B(n_11),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_14),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_252),
.C(n_13),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_11),
.Y(n_261)
);


endmodule