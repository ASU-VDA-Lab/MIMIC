module fake_jpeg_30928_n_516 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g115 ( 
.A(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_58),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_15),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_78),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_26),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_75),
.Y(n_118)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_1),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_90),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_14),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_19),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_77),
.Y(n_111)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_102),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_13),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_100),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_105),
.B(n_119),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_144),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_37),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_142),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_127),
.B(n_137),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_65),
.B(n_37),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_61),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_30),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_64),
.A2(n_32),
.B1(n_36),
.B2(n_24),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_32),
.B1(n_51),
.B2(n_36),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_72),
.B(n_27),
.C(n_36),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_62),
.Y(n_167)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_161),
.Y(n_217)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_113),
.B(n_25),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_163),
.B(n_171),
.Y(n_227)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_180),
.Y(n_226)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_208),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_48),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_182),
.B1(n_189),
.B2(n_193),
.Y(n_230)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_173),
.Y(n_241)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_130),
.Y(n_175)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_75),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_181),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_123),
.A2(n_48),
.B1(n_27),
.B2(n_53),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_84),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_184),
.B(n_192),
.Y(n_256)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_196),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_123),
.A2(n_48),
.B1(n_27),
.B2(n_52),
.Y(n_189)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_56),
.B1(n_95),
.B2(n_36),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_139),
.A2(n_101),
.B1(n_99),
.B2(n_98),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_130),
.A2(n_54),
.B(n_83),
.C(n_30),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_194),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_32),
.B1(n_51),
.B2(n_39),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_199),
.B1(n_213),
.B2(n_201),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_120),
.B(n_38),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_206),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_143),
.A2(n_96),
.B1(n_92),
.B2(n_88),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_114),
.B(n_38),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_200),
.Y(n_253)
);

CKINVDCx9p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_116),
.B(n_54),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_43),
.C(n_23),
.Y(n_239)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_136),
.B(n_47),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_108),
.B(n_33),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_47),
.Y(n_209)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_212),
.B(n_109),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_154),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_79),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_131),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_157),
.B1(n_125),
.B2(n_129),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_218),
.A2(n_243),
.B1(n_133),
.B2(n_183),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_135),
.B1(n_157),
.B2(n_125),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_161),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_184),
.A2(n_135),
.B1(n_118),
.B2(n_129),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_224),
.A2(n_258),
.B(n_226),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_115),
.B1(n_153),
.B2(n_156),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_246),
.B1(n_261),
.B2(n_164),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_262),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_117),
.B1(n_158),
.B2(n_145),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_185),
.A2(n_115),
.B1(n_153),
.B2(n_138),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_117),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_249),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_138),
.C(n_74),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_187),
.C(n_207),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_174),
.B(n_145),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_188),
.A2(n_79),
.A3(n_34),
.B1(n_46),
.B2(n_33),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_194),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_167),
.B(n_158),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_180),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_180),
.A2(n_33),
.B(n_43),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_186),
.A2(n_109),
.B1(n_133),
.B2(n_122),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_237),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_208),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_225),
.B1(n_222),
.B2(n_231),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_204),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_276),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_165),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_268),
.B(n_278),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_275),
.B1(n_277),
.B2(n_288),
.Y(n_305)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_255),
.A2(n_184),
.B1(n_80),
.B2(n_82),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_226),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_67),
.B1(n_85),
.B2(n_193),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_197),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_281),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_219),
.A2(n_164),
.B1(n_214),
.B2(n_215),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_280),
.A2(n_284),
.B1(n_217),
.B2(n_210),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_283),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_179),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_219),
.A2(n_196),
.B1(n_177),
.B2(n_212),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_234),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_289),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_236),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_287),
.B(n_296),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_199),
.B1(n_176),
.B2(n_168),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_162),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_191),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_227),
.B(n_181),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_294),
.A2(n_301),
.B(n_239),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_109),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_260),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_231),
.B1(n_242),
.B2(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_227),
.B(n_13),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_298),
.B(n_299),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_248),
.B(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

NAND2x1_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_224),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_34),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_302),
.B(n_303),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_259),
.B(n_34),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_286),
.C(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_314),
.C(n_320),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_308),
.A2(n_315),
.B1(n_317),
.B2(n_324),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_313),
.B(n_274),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_235),
.B(n_262),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_229),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_229),
.B1(n_170),
.B2(n_242),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_251),
.B1(n_220),
.B2(n_228),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_336),
.B1(n_288),
.B2(n_275),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_251),
.C(n_232),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_269),
.A2(n_232),
.B1(n_240),
.B2(n_217),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_321),
.A2(n_325),
.B1(n_296),
.B2(n_285),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_245),
.C(n_220),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_326),
.C(n_300),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_39),
.B1(n_21),
.B2(n_23),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_277),
.A2(n_217),
.B1(n_245),
.B2(n_228),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_272),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_252),
.B1(n_190),
.B2(n_241),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_148),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_340),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_196),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_268),
.Y(n_342)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_327),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_347),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_318),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_360),
.Y(n_392)
);

CKINVDCx10_ASAP7_75t_R g350 ( 
.A(n_306),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_307),
.A2(n_270),
.B(n_274),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_353),
.Y(n_388)
);

OAI21xp33_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_357),
.B(n_313),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_283),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_309),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_365),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_362),
.B1(n_368),
.B2(n_373),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_358),
.B(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_310),
.B(n_264),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_305),
.A2(n_323),
.B1(n_321),
.B2(n_316),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_319),
.B1(n_333),
.B2(n_328),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_301),
.B1(n_267),
.B2(n_279),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_364),
.A2(n_371),
.B1(n_42),
.B2(n_31),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_263),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_369),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_302),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_265),
.B1(n_303),
.B2(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_21),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_340),
.A2(n_298),
.B1(n_292),
.B2(n_271),
.Y(n_371)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_173),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_329),
.A2(n_292),
.B1(n_23),
.B2(n_43),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_320),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_386),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_376),
.B1(n_395),
.B2(n_366),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_363),
.A2(n_314),
.B1(n_326),
.B2(n_338),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_378),
.A2(n_355),
.B(n_349),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_342),
.B(n_339),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_380),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_360),
.B(n_330),
.Y(n_380)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

A2O1A1O1Ixp25_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_330),
.B(n_311),
.C(n_322),
.D(n_328),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_241),
.Y(n_389)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_352),
.A2(n_271),
.B(n_325),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_3),
.B(n_4),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_346),
.A2(n_252),
.B1(n_39),
.B2(n_35),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_35),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_396),
.Y(n_412)
);

OA21x2_ASAP7_75t_SL g397 ( 
.A1(n_351),
.A2(n_21),
.B(n_42),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_3),
.Y(n_427)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_367),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_399),
.B(n_350),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_2),
.Y(n_401)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_403),
.A2(n_346),
.B1(n_349),
.B2(n_369),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_404),
.A2(n_407),
.B1(n_409),
.B2(n_411),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_364),
.B1(n_348),
.B2(n_356),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_403),
.A2(n_396),
.B1(n_385),
.B2(n_384),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_402),
.A2(n_361),
.B1(n_370),
.B2(n_355),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_348),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_415),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_359),
.Y(n_414)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_414),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_417),
.A2(n_419),
.B1(n_387),
.B2(n_380),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_392),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_377),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_392),
.A2(n_372),
.B(n_341),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_42),
.C(n_31),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_376),
.C(n_396),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_31),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_428),
.Y(n_432)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_395),
.Y(n_444)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_426),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_427),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_374),
.B(n_3),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_433),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_384),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_414),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_437),
.A2(n_444),
.B1(n_447),
.B2(n_448),
.Y(n_452)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_439),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_422),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_441),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_406),
.C(n_428),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_445),
.C(n_446),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_391),
.C(n_385),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_391),
.C(n_377),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_388),
.B1(n_381),
.B2(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_404),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_436),
.A2(n_416),
.B(n_408),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_454),
.B(n_435),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_453),
.B(n_455),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_445),
.A2(n_394),
.B(n_412),
.Y(n_454)
);

XOR2x2_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_386),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_434),
.B(n_421),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_460),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_442),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_459),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_409),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_429),
.A2(n_405),
.B1(n_412),
.B2(n_387),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_420),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_463),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_425),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_393),
.C(n_382),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_443),
.C(n_438),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_459),
.B(n_461),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_472),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_462),
.A2(n_444),
.B1(n_443),
.B2(n_432),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_479),
.Y(n_492)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_393),
.B(n_432),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_456),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_4),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_465),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_464),
.B(n_4),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_480),
.B(n_6),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_456),
.B(n_5),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_481),
.Y(n_489)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_487),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_471),
.A2(n_465),
.B1(n_458),
.B2(n_8),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_491),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_493),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_6),
.C(n_7),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_6),
.C(n_8),
.Y(n_493)
);

MAJx2_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_473),
.C(n_475),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_496),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_469),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_499),
.A2(n_491),
.B(n_493),
.Y(n_503)
);

AOI31xp67_ASAP7_75t_L g500 ( 
.A1(n_487),
.A2(n_477),
.A3(n_469),
.B(n_478),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_500),
.B(n_501),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_475),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_497),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_505),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_488),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_489),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_509),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_506),
.C(n_494),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_495),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_510),
.Y(n_513)
);

AOI21xp33_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_492),
.B(n_486),
.Y(n_514)
);

O2A1O1Ixp33_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_515)
);

OAI211xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_11),
.B(n_414),
.C(n_510),
.Y(n_516)
);


endmodule