module fake_jpeg_9872_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_14),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_22),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_26),
.B1(n_28),
.B2(n_13),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_28),
.B1(n_20),
.B2(n_19),
.Y(n_79)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_43),
.C(n_29),
.Y(n_87)
);

NAND2x1_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_21),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_60),
.B(n_51),
.C(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_21),
.C(n_39),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.C(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_21),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_44),
.C(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_25),
.B1(n_19),
.B2(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_86),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_50),
.B1(n_49),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_94),
.B1(n_98),
.B2(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_64),
.B1(n_71),
.B2(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_25),
.B1(n_53),
.B2(n_15),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_41),
.B1(n_18),
.B2(n_17),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_61),
.B1(n_73),
.B2(n_65),
.Y(n_102)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_111),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_97),
.C(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_117),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_112),
.B1(n_99),
.B2(n_85),
.Y(n_131)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_65),
.B1(n_70),
.B2(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_118),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_96),
.B(n_102),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_128),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_116),
.C(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_109),
.C(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_135),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_101),
.B(n_98),
.C(n_100),
.D(n_38),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_68),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_59),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_143),
.Y(n_157)
);

NAND4xp25_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_59),
.C(n_104),
.D(n_68),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_153),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_129),
.B1(n_133),
.B2(n_122),
.Y(n_156)
);

AOI31xp67_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_109),
.A3(n_113),
.B(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_59),
.B1(n_38),
.B2(n_6),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_122),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_166),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_142),
.C(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_138),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_146),
.C(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_164),
.C(n_163),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_170),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_142),
.C(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_143),
.C(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_165),
.B1(n_159),
.B2(n_160),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_38),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_12),
.C(n_11),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_178),
.B1(n_174),
.B2(n_175),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_183),
.B1(n_8),
.B2(n_9),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_185),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_185),
.Y(n_187)
);


endmodule