module fake_netlist_6_2563_n_1827 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1827);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1827;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_82),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_39),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_72),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_9),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_35),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_12),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_121),
.Y(n_193)
);

INVx4_ASAP7_75t_R g194 ( 
.A(n_111),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_102),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_21),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_80),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_56),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_41),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_52),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_132),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_37),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_24),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_87),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_42),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_75),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_159),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_45),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_143),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_137),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_36),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_15),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

INVxp33_ASAP7_75t_R g237 ( 
.A(n_152),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_68),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_81),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_20),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_9),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_113),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_25),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_119),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_44),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_28),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_30),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_167),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_115),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_53),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_41),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_36),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_30),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_11),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_0),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_99),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_27),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_142),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_164),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_26),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_61),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_88),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_61),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_91),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_57),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_23),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_79),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_28),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_53),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_110),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_34),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_156),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_94),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_124),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_58),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_78),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_116),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_144),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_40),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_48),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_147),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_27),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_23),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_73),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_52),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_0),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_2),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_22),
.Y(n_312)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_146),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_108),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_109),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_39),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_59),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_57),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_6),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_45),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_130),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_14),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_85),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_46),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_24),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_154),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_157),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_140),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_55),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_20),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_112),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g333 ( 
.A(n_29),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_17),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_258),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_221),
.B(n_1),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_209),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_229),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_187),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_258),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_168),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_230),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_189),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_170),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_172),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_258),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_195),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_195),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_216),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_181),
.B(n_199),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_216),
.B(n_1),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_221),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_174),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_187),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_199),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_232),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_244),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_245),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_179),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_245),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_246),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_288),
.B(n_4),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_246),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_182),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_251),
.B(n_5),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_251),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_230),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_177),
.B(n_6),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_284),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_262),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_262),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_263),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_263),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_265),
.B(n_8),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_302),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_214),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_302),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_295),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_295),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_265),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_196),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_R g399 ( 
.A(n_306),
.B(n_114),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_266),
.B(n_8),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_198),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_202),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_205),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_215),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_267),
.B(n_10),
.Y(n_405)
);

BUFx6f_ASAP7_75t_SL g406 ( 
.A(n_252),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_267),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_173),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_270),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_270),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_217),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_223),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_227),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_228),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_238),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_239),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_335),
.A2(n_185),
.B(n_178),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_177),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_210),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_392),
.B(n_252),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_345),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_340),
.B(n_214),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_341),
.B(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_250),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_210),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_349),
.B(n_219),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_340),
.B(n_358),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_388),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_340),
.B(n_219),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_360),
.B(n_193),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_396),
.A2(n_207),
.B(n_171),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_366),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_352),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_353),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_353),
.B(n_290),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_343),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_367),
.B(n_240),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_342),
.B(n_296),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_367),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_378),
.B(n_290),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_368),
.B(n_242),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_368),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_370),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_371),
.B(n_243),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_378),
.B(n_171),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

BUFx8_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_387),
.B(n_207),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_384),
.B(n_247),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_343),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_387),
.B(n_178),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_336),
.B(n_282),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_385),
.B(n_185),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_385),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_347),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_348),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_426),
.B(n_491),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_372),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_483),
.B(n_338),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_424),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_350),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_361),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_490),
.A2(n_484),
.B1(n_477),
.B2(n_489),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_426),
.B(n_491),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_392),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_490),
.A2(n_484),
.B1(n_477),
.B2(n_489),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_454),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_483),
.B(n_369),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_377),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_425),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_483),
.B(n_398),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_418),
.B(n_401),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_425),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_418),
.B(n_402),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_470),
.B(n_490),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

AND3x2_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_354),
.C(n_346),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_441),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_470),
.B(n_404),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_490),
.A2(n_400),
.B1(n_405),
.B2(n_372),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_427),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_490),
.A2(n_400),
.B1(n_405),
.B2(n_357),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_470),
.B(n_411),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_394),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_419),
.B(n_412),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_426),
.B(n_491),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_419),
.B(n_413),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_487),
.B(n_414),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_429),
.A2(n_394),
.B1(n_373),
.B2(n_204),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_441),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_477),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_415),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_467),
.B(n_416),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_463),
.B(n_374),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_489),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_471),
.B(n_403),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_490),
.A2(n_357),
.B1(n_406),
.B2(n_283),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_420),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_490),
.B(n_399),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_429),
.B(n_339),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_439),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_471),
.B(n_391),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_439),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_475),
.A2(n_241),
.B1(n_276),
.B2(n_274),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_406),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_440),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_490),
.B(n_257),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_489),
.B(n_282),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_449),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_449),
.B(n_254),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_463),
.B(n_440),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_463),
.B(n_386),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_356),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_432),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_486),
.B(n_252),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_436),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_282),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_477),
.B(n_252),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_477),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_437),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_484),
.A2(n_406),
.B1(n_278),
.B2(n_283),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_437),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_488),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_453),
.B(n_255),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_488),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_439),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_473),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_473),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_484),
.A2(n_278),
.B1(n_332),
.B2(n_329),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_473),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_445),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_453),
.B(n_237),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_439),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_484),
.A2(n_286),
.B1(n_303),
.B2(n_304),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_427),
.B(n_269),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_445),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_488),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_473),
.B(n_282),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_444),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_433),
.B(n_272),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_433),
.A2(n_286),
.B1(n_332),
.B2(n_329),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_433),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_473),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_476),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_476),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_433),
.A2(n_188),
.B1(n_273),
.B2(n_331),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_433),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_457),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_417),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_457),
.B(n_356),
.Y(n_628)
);

CKINVDCx16_ASAP7_75t_R g629 ( 
.A(n_446),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_447),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_447),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_444),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_444),
.B(n_282),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_448),
.B(n_180),
.C(n_175),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_448),
.B(n_183),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_456),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_456),
.B(n_184),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_476),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_476),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_444),
.B(n_277),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_500),
.B(n_282),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_458),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_495),
.B(n_444),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_513),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_512),
.B(n_191),
.C(n_186),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_505),
.B(n_444),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_568),
.B(n_203),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_551),
.B(n_444),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_625),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_594),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_537),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_498),
.B(n_279),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_526),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_551),
.B(n_452),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_500),
.B(n_218),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_618),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_590),
.B(n_452),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_572),
.B(n_206),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_580),
.B(n_208),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_522),
.B(n_452),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_545),
.B(n_452),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_527),
.A2(n_451),
.B(n_435),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_494),
.B(n_458),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_580),
.B(n_552),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_503),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_452),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_508),
.A2(n_260),
.B1(n_190),
.B2(n_192),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_496),
.B(n_459),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_591),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_577),
.B(n_452),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_526),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_547),
.B(n_606),
.C(n_570),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_602),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_597),
.B(n_212),
.C(n_211),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_629),
.B(n_459),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_555),
.B(n_479),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_558),
.B(n_213),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_535),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_496),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_509),
.B(n_479),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_624),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_544),
.B(n_479),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_479),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_605),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_637),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_504),
.B(n_479),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

OAI221xp5_ASAP7_75t_L g699 ( 
.A1(n_603),
.A2(n_304),
.B1(n_303),
.B2(n_482),
.C(n_481),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_504),
.B(n_507),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_642),
.A2(n_451),
.B(n_435),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_556),
.B(n_469),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_525),
.B(n_220),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_611),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_507),
.B(n_479),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_517),
.B(n_479),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_517),
.B(n_518),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_520),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_579),
.B(n_469),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_510),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_518),
.B(n_451),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_556),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_542),
.B(n_506),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_515),
.B(n_222),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_630),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_533),
.B(n_224),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_511),
.B(n_571),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_231),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_631),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_637),
.B(n_235),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_637),
.B(n_236),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_536),
.A2(n_259),
.B1(n_190),
.B2(n_192),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_596),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_596),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_598),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_500),
.B(n_218),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_524),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_540),
.B(n_451),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_579),
.B(n_478),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_564),
.B(n_574),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_627),
.A2(n_417),
.B1(n_455),
.B2(n_200),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_583),
.B(n_248),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_540),
.B(n_460),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_546),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_553),
.B(n_460),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_554),
.B(n_563),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_627),
.A2(n_417),
.B1(n_455),
.B2(n_200),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_624),
.B(n_478),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_557),
.B(n_218),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_510),
.B(n_480),
.Y(n_742)
);

NOR2x1p5_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_249),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_608),
.A2(n_417),
.B1(n_455),
.B2(n_271),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_546),
.B(n_326),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_554),
.B(n_460),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_497),
.B(n_253),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_563),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_578),
.B(n_460),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_612),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_597),
.A2(n_297),
.B1(n_285),
.B2(n_292),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_612),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_546),
.B(n_480),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_578),
.B(n_581),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_541),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_581),
.B(n_417),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_550),
.B(n_261),
.C(n_334),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_619),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_497),
.B(n_264),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_619),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_557),
.B(n_559),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_636),
.B(n_481),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_557),
.B(n_218),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_497),
.B(n_176),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_585),
.B(n_586),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_529),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_585),
.B(n_472),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_586),
.B(n_472),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_530),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_589),
.B(n_268),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_592),
.B(n_472),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_592),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_523),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_623),
.A2(n_233),
.B1(n_321),
.B2(n_314),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_538),
.B(n_218),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_493),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_574),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_576),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_632),
.B(n_474),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_523),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_528),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_548),
.A2(n_233),
.B1(n_321),
.B2(n_314),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_575),
.B(n_482),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_514),
.B(n_176),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_528),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_543),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_616),
.B(n_197),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_576),
.B(n_485),
.Y(n_789)
);

AND2x2_ASAP7_75t_SL g790 ( 
.A(n_593),
.B(n_201),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_638),
.B(n_201),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_543),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_499),
.B(n_225),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_560),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_573),
.A2(n_465),
.B(n_464),
.Y(n_795)
);

OR2x2_ASAP7_75t_SL g796 ( 
.A(n_635),
.B(n_225),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_493),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_560),
.Y(n_798)
);

AO221x1_ASAP7_75t_L g799 ( 
.A1(n_499),
.A2(n_234),
.B1(n_226),
.B2(n_259),
.C(n_271),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_566),
.B(n_485),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_499),
.B(n_226),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_521),
.B(n_492),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_595),
.B(n_313),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_595),
.B(n_313),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_574),
.A2(n_328),
.B1(n_327),
.B2(n_323),
.Y(n_805)
);

INVxp33_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_501),
.B(n_516),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_531),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_501),
.B(n_234),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_501),
.B(n_516),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_671),
.A2(n_307),
.B(n_280),
.Y(n_811)
);

BUFx12f_ASAP7_75t_L g812 ( 
.A(n_654),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_516),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_740),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_667),
.A2(n_588),
.B(n_534),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_740),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_652),
.B(n_519),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_668),
.A2(n_588),
.B(n_534),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_652),
.B(n_519),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_647),
.A2(n_588),
.B(n_534),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_662),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_762),
.B(n_519),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_717),
.A2(n_275),
.B1(n_280),
.B2(n_287),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_670),
.B(n_531),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_681),
.B(n_531),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_686),
.A2(n_275),
.B(n_298),
.C(n_287),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_708),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_686),
.A2(n_307),
.B(n_298),
.C(n_293),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_651),
.A2(n_567),
.B(n_582),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_791),
.A2(n_726),
.B(n_661),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_674),
.A2(n_567),
.B(n_582),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_679),
.A2(n_567),
.B(n_582),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_492),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_806),
.A2(n_293),
.B1(n_599),
.B2(n_569),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_689),
.B(n_569),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_712),
.B(n_531),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_689),
.B(n_569),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_690),
.B(n_599),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_661),
.A2(n_640),
.B(n_621),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_690),
.B(n_599),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_685),
.A2(n_660),
.B(n_653),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_713),
.B(n_502),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_713),
.B(n_502),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_696),
.B(n_532),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_756),
.A2(n_621),
.B(n_640),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_567),
.B(n_532),
.Y(n_847)
);

AND3x2_ASAP7_75t_L g848 ( 
.A(n_745),
.B(n_397),
.C(n_409),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_669),
.A2(n_693),
.B(n_691),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_740),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_729),
.B(n_622),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_696),
.B(n_532),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_700),
.A2(n_567),
.B(n_532),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_727),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_707),
.A2(n_532),
.B(n_561),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_662),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_680),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_806),
.B(n_622),
.Y(n_858)
);

AOI21xp33_ASAP7_75t_L g859 ( 
.A1(n_703),
.A2(n_281),
.B(n_289),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_787),
.B(n_626),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_769),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_787),
.B(n_626),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_676),
.A2(n_613),
.B(n_565),
.C(n_584),
.Y(n_863)
);

OAI21xp33_ASAP7_75t_SL g864 ( 
.A1(n_761),
.A2(n_775),
.B(n_739),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_684),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_677),
.B(n_561),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_677),
.B(n_561),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_607),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_738),
.B(n_607),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_680),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_692),
.B(n_607),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_666),
.B(n_386),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_666),
.B(n_395),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_644),
.A2(n_641),
.B(n_639),
.Y(n_874)
);

NOR2x1_ASAP7_75t_R g875 ( 
.A(n_710),
.B(n_291),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_714),
.A2(n_574),
.B1(n_587),
.B2(n_634),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_687),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_703),
.A2(n_641),
.B(n_639),
.C(n_634),
.Y(n_878)
);

AO21x1_ASAP7_75t_L g879 ( 
.A1(n_726),
.A2(n_613),
.B(n_620),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_644),
.A2(n_601),
.B(n_620),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_730),
.A2(n_607),
.B(n_615),
.Y(n_881)
);

AOI21xp33_ASAP7_75t_L g882 ( 
.A1(n_733),
.A2(n_317),
.B(n_316),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_694),
.A2(n_604),
.B(n_600),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_692),
.B(n_607),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_688),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_754),
.B(n_615),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_765),
.B(n_714),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_716),
.B(n_718),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_753),
.B(n_395),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_716),
.A2(n_574),
.B1(n_587),
.B2(n_614),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_687),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_718),
.B(n_615),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_755),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_761),
.A2(n_615),
.B(n_601),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_735),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_779),
.A2(n_600),
.B(n_614),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_692),
.A2(n_604),
.B(n_562),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_692),
.B(n_574),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_789),
.B(n_299),
.Y(n_899)
);

CKINVDCx11_ASAP7_75t_R g900 ( 
.A(n_784),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_665),
.B(n_397),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_662),
.B(n_562),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_770),
.A2(n_584),
.B(n_565),
.C(n_315),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_770),
.A2(n_294),
.B(n_461),
.C(n_465),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_643),
.B(n_313),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_665),
.B(n_300),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_643),
.B(n_313),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_731),
.A2(n_587),
.B(n_633),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_SL g909 ( 
.A1(n_775),
.A2(n_410),
.B(n_407),
.C(n_409),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_657),
.B(n_407),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_672),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_733),
.A2(n_461),
.B(n_462),
.C(n_465),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_736),
.B(n_587),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_697),
.A2(n_464),
.B(n_462),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_705),
.A2(n_464),
.B(n_462),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_777),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_777),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_706),
.A2(n_461),
.B(n_587),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_711),
.A2(n_808),
.B(n_807),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_777),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_720),
.A2(n_319),
.B(n_305),
.C(n_308),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_808),
.A2(n_587),
.B(n_194),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_810),
.A2(n_633),
.B(n_410),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_748),
.Y(n_924)
);

CKINVDCx6p67_ASAP7_75t_R g925 ( 
.A(n_784),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_783),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_720),
.B(n_326),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_672),
.B(n_648),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_731),
.A2(n_633),
.B(n_330),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_721),
.B(n_326),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_748),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_772),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_742),
.B(n_301),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_739),
.A2(n_633),
.B(n_325),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_790),
.A2(n_313),
.B1(n_326),
.B2(n_633),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_645),
.B(n_309),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_772),
.B(n_633),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_709),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_741),
.A2(n_324),
.B(n_322),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_709),
.B(n_320),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_649),
.A2(n_318),
.B1(n_311),
.B2(n_310),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_701),
.A2(n_63),
.B(n_158),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_657),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_782),
.A2(n_11),
.B(n_13),
.C(n_16),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_795),
.A2(n_746),
.B(n_749),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_673),
.B(n_13),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_778),
.B(n_802),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_SL g948 ( 
.A(n_658),
.B(n_66),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_741),
.A2(n_74),
.B(n_155),
.Y(n_949)
);

OAI321xp33_ASAP7_75t_L g950 ( 
.A1(n_782),
.A2(n_17),
.A3(n_18),
.B1(n_26),
.B2(n_29),
.C(n_31),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_763),
.A2(n_77),
.B(n_139),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_723),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_722),
.A2(n_18),
.B(n_31),
.C(n_32),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_675),
.B(n_678),
.Y(n_954)
);

AND2x6_ASAP7_75t_L g955 ( 
.A(n_800),
.B(n_656),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_790),
.B(n_89),
.Y(n_956)
);

INVx11_ASAP7_75t_L g957 ( 
.A(n_796),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_721),
.B(n_90),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_763),
.A2(n_162),
.B(n_133),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_682),
.B(n_32),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_774),
.A2(n_33),
.B(n_35),
.C(n_38),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_728),
.A2(n_95),
.B(n_128),
.Y(n_962)
);

AO21x1_ASAP7_75t_L g963 ( 
.A1(n_774),
.A2(n_42),
.B(n_44),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_747),
.B(n_98),
.Y(n_964)
);

BUFx4f_ASAP7_75t_L g965 ( 
.A(n_657),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_734),
.A2(n_100),
.B(n_127),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_695),
.B(n_47),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_698),
.A2(n_131),
.B1(n_126),
.B2(n_125),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_646),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_704),
.B(n_47),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_715),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_737),
.A2(n_123),
.B(n_122),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_767),
.A2(n_106),
.B(n_103),
.Y(n_973)
);

O2A1O1Ixp5_ASAP7_75t_L g974 ( 
.A1(n_788),
.A2(n_50),
.B(n_51),
.C(n_54),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_719),
.B(n_51),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_699),
.A2(n_54),
.B(n_55),
.C(n_58),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_747),
.B(n_759),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_768),
.A2(n_59),
.B(n_60),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_724),
.B(n_60),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_725),
.B(n_62),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_771),
.A2(n_655),
.B(n_646),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_655),
.B(n_62),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_732),
.B(n_758),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_750),
.A2(n_760),
.B(n_752),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_776),
.A2(n_797),
.B(n_798),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_759),
.B(n_773),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_776),
.A2(n_797),
.B(n_786),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_780),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_781),
.B(n_785),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_744),
.A2(n_764),
.B1(n_784),
.B2(n_650),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_792),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_794),
.A2(n_804),
.B(n_803),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_803),
.A2(n_804),
.B(n_744),
.Y(n_994)
);

NOR2x1_ASAP7_75t_R g995 ( 
.A(n_861),
.B(n_766),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_823),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_891),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_924),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_888),
.A2(n_683),
.B(n_764),
.C(n_757),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_857),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_812),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_977),
.B(n_743),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_887),
.B(n_751),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_938),
.B(n_805),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_826),
.A2(n_799),
.B(n_846),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_872),
.B(n_873),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_817),
.A2(n_814),
.B1(n_816),
.B2(n_850),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_901),
.B(n_889),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_906),
.B(n_859),
.C(n_882),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_SL g1010 ( 
.A1(n_956),
.A2(n_908),
.B(n_986),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_817),
.A2(n_956),
.B1(n_868),
.B2(n_822),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_892),
.A2(n_849),
.B(n_842),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_895),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_906),
.B(n_947),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_938),
.B(n_954),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_911),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_864),
.A2(n_819),
.B(n_992),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_926),
.B(n_865),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_990),
.A2(n_986),
.B1(n_865),
.B2(n_930),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_931),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_899),
.A2(n_885),
.B1(n_971),
.B2(n_854),
.Y(n_1021)
);

INVx3_ASAP7_75t_SL g1022 ( 
.A(n_925),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_858),
.A2(n_899),
.B(n_942),
.C(n_933),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_954),
.B(n_926),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_858),
.B(n_813),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_916),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_936),
.B(n_933),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_869),
.A2(n_886),
.B(n_844),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_SL g1029 ( 
.A1(n_927),
.A2(n_958),
.B(n_824),
.C(n_964),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_870),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_SL g1031 ( 
.A1(n_945),
.A2(n_936),
.B(n_836),
.C(n_841),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_828),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_828),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_854),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_877),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_910),
.B(n_971),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_994),
.A2(n_984),
.B(n_958),
.C(n_921),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_910),
.B(n_821),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_988),
.B(n_843),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_916),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_811),
.A2(n_831),
.B(n_879),
.C(n_840),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_952),
.B(n_851),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_893),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_834),
.B(n_893),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_815),
.A2(n_818),
.B(n_820),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_940),
.B(n_957),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_875),
.B(n_941),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_881),
.A2(n_894),
.B(n_830),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_900),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_832),
.A2(n_833),
.B(n_855),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_910),
.B(n_943),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_946),
.A2(n_960),
.B(n_967),
.C(n_970),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_916),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_827),
.A2(n_829),
.B(n_982),
.C(n_950),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_969),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_983),
.B(n_860),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_989),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_862),
.B(n_911),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_991),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_916),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_948),
.A2(n_955),
.B1(n_867),
.B2(n_866),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_991),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_838),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_982),
.A2(n_845),
.B1(n_852),
.B2(n_928),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_917),
.B(n_920),
.Y(n_1067)
);

OAI22x1_ASAP7_75t_L g1068 ( 
.A1(n_928),
.A2(n_963),
.B1(n_848),
.B2(n_837),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_856),
.B(n_836),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_839),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_943),
.B(n_965),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_L g1072 ( 
.A1(n_848),
.A2(n_944),
.B1(n_979),
.B2(n_980),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_841),
.A2(n_993),
.B(n_904),
.C(n_903),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_835),
.B(n_905),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_909),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_985),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_953),
.A2(n_929),
.B(n_934),
.C(n_976),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_917),
.B(n_920),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_974),
.A2(n_961),
.B(n_912),
.C(n_978),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_965),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_917),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_853),
.A2(n_919),
.B(n_883),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_987),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_917),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_955),
.B(n_981),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_955),
.B(n_935),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_939),
.B(n_935),
.C(n_974),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_920),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_905),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_878),
.A2(n_907),
.B(n_968),
.C(n_825),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_876),
.B(n_890),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_907),
.B(n_913),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_902),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_847),
.A2(n_898),
.B(n_896),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_884),
.B(n_871),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_884),
.A2(n_863),
.B(n_897),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_937),
.B(n_918),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_902),
.B(n_914),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_922),
.A2(n_915),
.B(n_923),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_874),
.B(n_880),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_973),
.A2(n_972),
.B(n_966),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_902),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_902),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_902),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_949),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_962),
.A2(n_951),
.B(n_959),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_888),
.B(n_671),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_828),
.Y(n_1109)
);

CKINVDCx8_ASAP7_75t_R g1110 ( 
.A(n_861),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_885),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_892),
.A2(n_500),
.B(n_888),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_889),
.B(n_671),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_888),
.B(n_671),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_888),
.B(n_671),
.C(n_686),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_888),
.B(n_671),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_888),
.A2(n_671),
.B(n_906),
.C(n_652),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_892),
.A2(n_500),
.B(n_888),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_888),
.A2(n_958),
.B(n_829),
.C(n_827),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_881),
.A2(n_894),
.B(n_830),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_888),
.B(n_671),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_888),
.B(n_671),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_892),
.A2(n_500),
.B(n_888),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_888),
.A2(n_671),
.B(n_887),
.C(n_824),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_888),
.B(n_671),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_916),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_888),
.B(n_671),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_888),
.B(n_671),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_812),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_821),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_916),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_888),
.B(n_671),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_888),
.A2(n_671),
.B1(n_887),
.B2(n_717),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_888),
.A2(n_671),
.B(n_906),
.C(n_652),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_889),
.B(n_671),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_888),
.B(n_671),
.Y(n_1136)
);

NOR2x1p5_ASAP7_75t_L g1137 ( 
.A(n_861),
.B(n_769),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_888),
.B(n_671),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_828),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_888),
.B(n_671),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_888),
.A2(n_671),
.B(n_887),
.C(n_824),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_SL g1142 ( 
.A(n_1110),
.B(n_995),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1026),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1034),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_997),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1038),
.B(n_1015),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_1016),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_1047),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_1082),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_1082),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1117),
.A2(n_1134),
.B(n_1140),
.C(n_1023),
.Y(n_1154)
);

OAI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1006),
.A2(n_1125),
.B1(n_1128),
.B2(n_1108),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1032),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1011),
.A2(n_1077),
.A3(n_1037),
.B(n_1073),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1116),
.B(n_1121),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1009),
.A2(n_1141),
.B(n_1124),
.C(n_1115),
.Y(n_1159)
);

NAND3x1_ASAP7_75t_L g1160 ( 
.A(n_1048),
.B(n_1009),
.C(n_1052),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1138),
.B(n_1113),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1124),
.A2(n_1141),
.B(n_1003),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_998),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_1041),
.A2(n_1028),
.B(n_1097),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1008),
.B(n_1033),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1135),
.B(n_1114),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1122),
.B(n_1136),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1112),
.A2(n_1118),
.B(n_1123),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1111),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1133),
.B(n_1059),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1115),
.A2(n_1053),
.B(n_1025),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1013),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1041),
.A2(n_1028),
.B(n_1097),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1109),
.B(n_1139),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_1045),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1001),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1020),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1112),
.A2(n_1118),
.B(n_1123),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_999),
.B(n_1019),
.C(n_1002),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1046),
.A2(n_1031),
.B(n_1102),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1058),
.B(n_1042),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1029),
.A2(n_1010),
.B(n_1093),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1102),
.A2(n_1051),
.B(n_1119),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1039),
.A2(n_1057),
.B1(n_1021),
.B2(n_1086),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1044),
.Y(n_1186)
);

AOI221x1_ASAP7_75t_L g1187 ( 
.A1(n_1072),
.A2(n_1088),
.B1(n_1068),
.B2(n_1107),
.C(n_1100),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1043),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1016),
.A2(n_1063),
.B1(n_1074),
.B2(n_1060),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1129),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1018),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1109),
.B(n_1139),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_1080),
.B(n_1024),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1070),
.B(n_1065),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1107),
.A2(n_1098),
.B(n_1085),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_999),
.B(n_1055),
.C(n_1079),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1050),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1092),
.A2(n_1091),
.B(n_1083),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_996),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1015),
.A2(n_1076),
.B1(n_1061),
.B2(n_1064),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1091),
.A2(n_1099),
.B(n_1004),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1101),
.A2(n_1066),
.A3(n_1007),
.B(n_1106),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1005),
.A2(n_1069),
.B(n_1075),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1137),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1088),
.A2(n_1070),
.B1(n_1090),
.B2(n_1000),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1079),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1096),
.A2(n_1106),
.B1(n_1093),
.B2(n_1036),
.C(n_1038),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1036),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1055),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1071),
.B(n_1094),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_1081),
.B(n_1126),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1103),
.A2(n_1090),
.B1(n_1130),
.B2(n_1030),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1035),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_L g1215 ( 
.A(n_1131),
.B(n_1084),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1022),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1089),
.B(n_1126),
.Y(n_1217)
);

AOI221x1_ASAP7_75t_L g1218 ( 
.A1(n_1026),
.A2(n_1040),
.B1(n_1054),
.B2(n_1062),
.C(n_1084),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1022),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1040),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1131),
.A2(n_1054),
.B(n_1062),
.Y(n_1221)
);

INVx3_ASAP7_75t_SL g1222 ( 
.A(n_1054),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1062),
.A2(n_1084),
.B(n_1131),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1087),
.B(n_1127),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1023),
.A2(n_811),
.A3(n_1017),
.B(n_1012),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1009),
.B(n_1117),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1230)
);

BUFx2_ASAP7_75t_R g1231 ( 
.A(n_1110),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1033),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1094),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1023),
.A2(n_811),
.A3(n_1017),
.B(n_1012),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1110),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1117),
.A2(n_1134),
.B(n_1027),
.C(n_1023),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1032),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1023),
.A2(n_811),
.A3(n_1017),
.B(n_1012),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1032),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1117),
.A2(n_1134),
.B(n_1023),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1117),
.A2(n_782),
.B1(n_1134),
.B2(n_1027),
.C(n_774),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1034),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1009),
.A2(n_1027),
.B1(n_686),
.B2(n_1014),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1113),
.B(n_1135),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_L g1254 ( 
.A(n_1137),
.B(n_696),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1027),
.B(n_1127),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1034),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1056),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1027),
.B(n_1127),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1041),
.A2(n_1017),
.B(n_1082),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1117),
.A2(n_1134),
.B(n_1027),
.C(n_1132),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1113),
.B(n_1135),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1113),
.B(n_1135),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1117),
.A2(n_1134),
.B(n_1023),
.C(n_888),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1034),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_997),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1047),
.B(n_708),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1056),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1041),
.A2(n_1017),
.B(n_1082),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1027),
.A2(n_671),
.B1(n_380),
.B2(n_388),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1045),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1032),
.Y(n_1279)
);

OAI21xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1006),
.A2(n_956),
.B(n_888),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1095),
.A2(n_1120),
.B(n_1049),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1026),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1056),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1056),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1001),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1009),
.A2(n_1027),
.B1(n_686),
.B2(n_1014),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1012),
.A2(n_1017),
.B(n_888),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1009),
.A2(n_1127),
.B1(n_1140),
.B2(n_1132),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1146),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1170),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1235),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1257),
.A2(n_1260),
.B1(n_1291),
.B2(n_1247),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1274),
.A2(n_1257),
.B1(n_1260),
.B2(n_1196),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1173),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1291),
.A2(n_1289),
.B1(n_1226),
.B2(n_1285),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1177),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1164),
.Y(n_1300)
);

BUFx4f_ASAP7_75t_SL g1301 ( 
.A(n_1288),
.Y(n_1301)
);

INVx8_ASAP7_75t_L g1302 ( 
.A(n_1143),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_1230),
.B1(n_1276),
.B2(n_1283),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1178),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1186),
.Y(n_1305)
);

BUFx2_ASAP7_75t_SL g1306 ( 
.A(n_1237),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_SL g1307 ( 
.A(n_1222),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1226),
.A2(n_1228),
.B1(n_1145),
.B2(n_1242),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1246),
.B(n_1250),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1253),
.B(n_1256),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1180),
.A2(n_1162),
.B1(n_1284),
.B2(n_1172),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1155),
.A2(n_1171),
.B1(n_1280),
.B2(n_1167),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_SL g1313 ( 
.A(n_1222),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1217),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1197),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1149),
.A2(n_1182),
.B1(n_1248),
.B2(n_1264),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1156),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1143),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1175),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1204),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1155),
.A2(n_1168),
.B1(n_1158),
.B2(n_1198),
.Y(n_1321)
);

OAI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1161),
.A2(n_1166),
.B1(n_1149),
.B2(n_1224),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1245),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1231),
.Y(n_1324)
);

CKINVDCx14_ASAP7_75t_R g1325 ( 
.A(n_1268),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1198),
.A2(n_1265),
.B1(n_1201),
.B2(n_1185),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1183),
.A2(n_1142),
.B1(n_1189),
.B2(n_1201),
.Y(n_1327)
);

INVx8_ASAP7_75t_L g1328 ( 
.A(n_1220),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1176),
.B1(n_1275),
.B2(n_1191),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1220),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1220),
.Y(n_1331)
);

CKINVDCx6p67_ASAP7_75t_R g1332 ( 
.A(n_1219),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1217),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1279),
.Y(n_1334)
);

INVx3_ASAP7_75t_SL g1335 ( 
.A(n_1144),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1220),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1160),
.A2(n_1270),
.B1(n_1258),
.B2(n_1193),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1216),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1232),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1269),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1259),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1263),
.A2(n_1154),
.B1(n_1176),
.B2(n_1275),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1148),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1232),
.A2(n_1194),
.B1(n_1199),
.B2(n_1188),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1150),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_1159),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1150),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1261),
.A2(n_1273),
.B1(n_1184),
.B2(n_1236),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1272),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1190),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1236),
.A2(n_1205),
.B1(n_1192),
.B2(n_1175),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1205),
.A2(n_1287),
.B1(n_1286),
.B2(n_1192),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1207),
.A2(n_1187),
.B1(n_1200),
.B2(n_1240),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1261),
.A2(n_1273),
.B1(n_1184),
.B2(n_1267),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1148),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_SL g1357 ( 
.A(n_1282),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1282),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1244),
.A2(n_1174),
.B1(n_1165),
.B2(n_1262),
.Y(n_1359)
);

BUFx10_ASAP7_75t_L g1360 ( 
.A(n_1282),
.Y(n_1360)
);

BUFx4f_ASAP7_75t_SL g1361 ( 
.A(n_1214),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1210),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1254),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1229),
.A2(n_1290),
.B1(n_1277),
.B2(n_1252),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1163),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_1214),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1212),
.A2(n_1215),
.B1(n_1211),
.B2(n_1233),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1163),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1229),
.A2(n_1277),
.B1(n_1238),
.B2(n_1243),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1233),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1238),
.A2(n_1290),
.B1(n_1262),
.B2(n_1252),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1243),
.A2(n_1249),
.B1(n_1174),
.B2(n_1165),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_1181),
.B2(n_1169),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1218),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1221),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1203),
.A2(n_1181),
.B1(n_1169),
.B2(n_1179),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1221),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1223),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1209),
.B(n_1213),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1223),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1206),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1202),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1202),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1157),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1157),
.A2(n_1195),
.B1(n_1239),
.B2(n_1225),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1225),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1157),
.A2(n_1151),
.B1(n_1281),
.B2(n_1227),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1255),
.B1(n_1271),
.B2(n_1266),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1251),
.A2(n_1278),
.B1(n_1234),
.B2(n_1239),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1225),
.A2(n_1274),
.B1(n_956),
.B2(n_1260),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1234),
.A2(n_1009),
.B1(n_1260),
.B2(n_1257),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1239),
.A2(n_1132),
.B1(n_1140),
.B2(n_1127),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1235),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1170),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1274),
.A2(n_956),
.B1(n_1260),
.B2(n_1257),
.Y(n_1395)
);

BUFx2_ASAP7_75t_SL g1396 ( 
.A(n_1173),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1173),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1235),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1143),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1257),
.A2(n_1027),
.B(n_671),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1146),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1257),
.B(n_1260),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1247),
.A2(n_1027),
.B1(n_1289),
.B2(n_1230),
.Y(n_1403)
);

CKINVDCx8_ASAP7_75t_R g1404 ( 
.A(n_1197),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1235),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1257),
.A2(n_1009),
.B1(n_1260),
.B2(n_1291),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1143),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_1173),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1257),
.A2(n_1009),
.B1(n_1027),
.B2(n_686),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1257),
.A2(n_1009),
.B1(n_1260),
.B2(n_1291),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1381),
.Y(n_1411)
);

INVxp33_ASAP7_75t_L g1412 ( 
.A(n_1317),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1395),
.A2(n_1296),
.B1(n_1390),
.B2(n_1410),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1395),
.A2(n_1296),
.B1(n_1295),
.B2(n_1410),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1402),
.B(n_1335),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1339),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1381),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1388),
.A2(n_1387),
.B(n_1379),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1375),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1390),
.A2(n_1406),
.B1(n_1295),
.B2(n_1403),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1343),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1386),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1384),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1406),
.B(n_1400),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1409),
.B(n_1303),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1382),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1378),
.Y(n_1428)
);

CKINVDCx6p67_ASAP7_75t_R g1429 ( 
.A(n_1405),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1387),
.A2(n_1379),
.B(n_1364),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1381),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1391),
.B(n_1326),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1377),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1292),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1403),
.B(n_1309),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_SL g1436 ( 
.A(n_1404),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1300),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1304),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_SL g1439 ( 
.A(n_1324),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1377),
.B(n_1380),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1380),
.B(n_1305),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1394),
.Y(n_1442)
);

NAND2x1_ASAP7_75t_L g1443 ( 
.A(n_1326),
.B(n_1368),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1347),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1393),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1341),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1322),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1354),
.A2(n_1392),
.B(n_1322),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1352),
.A2(n_1362),
.B1(n_1325),
.B2(n_1313),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1374),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1401),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1298),
.A2(n_1311),
.B1(n_1308),
.B2(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1376),
.Y(n_1453)
);

INVx3_ASAP7_75t_SL g1454 ( 
.A(n_1346),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1345),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1385),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1391),
.B(n_1329),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_1312),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1385),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1370),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1349),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1312),
.B(n_1327),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1373),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1373),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1359),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1359),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1355),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1355),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1364),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1310),
.B(n_1308),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1369),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1298),
.B(n_1321),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1372),
.A2(n_1371),
.A3(n_1369),
.B(n_1389),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1371),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1342),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1321),
.B(n_1316),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1335),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1372),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1319),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1389),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1350),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1365),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1316),
.B(n_1329),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1353),
.B(n_1337),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1353),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1367),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1348),
.A2(n_1325),
.B1(n_1307),
.B2(n_1313),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1357),
.A2(n_1360),
.B(n_1328),
.Y(n_1489)
);

AOI21xp33_ASAP7_75t_L g1490 ( 
.A1(n_1363),
.A2(n_1323),
.B(n_1358),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1319),
.A2(n_1331),
.B(n_1407),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1429),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1443),
.B(n_1306),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1415),
.B(n_1478),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1456),
.B(n_1407),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1444),
.B(n_1356),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1420),
.B(n_1344),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1412),
.B(n_1297),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1451),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1456),
.B(n_1331),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1441),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1417),
.B(n_1397),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1414),
.A2(n_1344),
.B1(n_1338),
.B2(n_1299),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1416),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1439),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1426),
.B(n_1333),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1451),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1459),
.B(n_1407),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1413),
.A2(n_1332),
.B1(n_1294),
.B2(n_1333),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1452),
.A2(n_1408),
.B1(n_1396),
.B2(n_1366),
.C(n_1399),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1434),
.Y(n_1512)
);

AND2x6_ASAP7_75t_L g1513 ( 
.A(n_1463),
.B(n_1477),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1453),
.B(n_1351),
.Y(n_1514)
);

NAND4xp25_ASAP7_75t_L g1515 ( 
.A(n_1421),
.B(n_1330),
.C(n_1340),
.D(n_1336),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1453),
.B(n_1331),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1436),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1461),
.B(n_1399),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1434),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1441),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1463),
.A2(n_1366),
.B1(n_1399),
.B2(n_1340),
.C(n_1318),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1458),
.A2(n_1302),
.B(n_1328),
.C(n_1307),
.Y(n_1522)
);

AND2x6_ASAP7_75t_L g1523 ( 
.A(n_1477),
.B(n_1314),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_SL g1524 ( 
.A1(n_1473),
.A2(n_1361),
.B(n_1302),
.C(n_1314),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1422),
.B(n_1334),
.C(n_1361),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1432),
.A2(n_1333),
.B(n_1301),
.C(n_1398),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1441),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1455),
.B(n_1320),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1442),
.B(n_1315),
.Y(n_1529)
);

NAND4xp25_ASAP7_75t_L g1530 ( 
.A(n_1485),
.B(n_1301),
.C(n_1425),
.D(n_1487),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1441),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1429),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1484),
.B(n_1447),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1430),
.A2(n_1419),
.B(n_1411),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1447),
.B(n_1432),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1491),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1430),
.A2(n_1419),
.B(n_1479),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1480),
.B(n_1428),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1462),
.B(n_1466),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1476),
.B(n_1486),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1428),
.B(n_1454),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1424),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1418),
.A2(n_1433),
.B(n_1431),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1443),
.B(n_1440),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1486),
.B(n_1482),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1483),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1479),
.A2(n_1475),
.B(n_1472),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1449),
.A2(n_1472),
.B(n_1470),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1535),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1508),
.B(n_1450),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1512),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1493),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1550),
.B(n_1464),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1519),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1537),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1543),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1543),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1474),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1501),
.B(n_1418),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1538),
.B(n_1474),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1545),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1493),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1474),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1542),
.B(n_1474),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1550),
.B(n_1464),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1499),
.B(n_1427),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1516),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1530),
.A2(n_1448),
.B1(n_1450),
.B2(n_1457),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1546),
.Y(n_1572)
);

AND2x2_ASAP7_75t_SL g1573 ( 
.A(n_1534),
.B(n_1423),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1507),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1550),
.B(n_1465),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1520),
.B(n_1527),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1551),
.A2(n_1448),
.B1(n_1450),
.B2(n_1457),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1510),
.A2(n_1428),
.B1(n_1475),
.B2(n_1469),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1540),
.B(n_1469),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1493),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1503),
.A2(n_1468),
.B1(n_1460),
.B2(n_1446),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1576),
.Y(n_1583)
);

AOI33xp33_ASAP7_75t_L g1584 ( 
.A1(n_1577),
.A2(n_1531),
.A3(n_1536),
.B1(n_1516),
.B2(n_1532),
.B3(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1564),
.Y(n_1585)
);

AOI33xp33_ASAP7_75t_L g1586 ( 
.A1(n_1577),
.A2(n_1531),
.A3(n_1518),
.B1(n_1495),
.B2(n_1500),
.B3(n_1509),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1578),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1558),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1427),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.Y(n_1593)
);

NAND2x1_ASAP7_75t_L g1594 ( 
.A(n_1572),
.B(n_1547),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1570),
.B(n_1547),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1576),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1504),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1571),
.A2(n_1511),
.B1(n_1506),
.B2(n_1525),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1571),
.B(n_1494),
.C(n_1539),
.D(n_1514),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1564),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1557),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1555),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1547),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1579),
.A2(n_1513),
.B1(n_1515),
.B2(n_1523),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1579),
.A2(n_1526),
.B1(n_1496),
.B2(n_1521),
.C(n_1522),
.Y(n_1607)
);

NOR3xp33_ASAP7_75t_L g1608 ( 
.A(n_1582),
.B(n_1490),
.C(n_1526),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1553),
.A2(n_1513),
.B1(n_1523),
.B2(n_1497),
.Y(n_1609)
);

AND2x4_ASAP7_75t_SL g1610 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1541),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_1548),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1552),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1560),
.B(n_1481),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1597),
.B(n_1583),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1611),
.B(n_1574),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1588),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1625)
);

CKINVDCx14_ASAP7_75t_R g1626 ( 
.A(n_1595),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1612),
.B(n_1593),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1611),
.B(n_1574),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1615),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1613),
.B(n_1555),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1585),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1590),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1592),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1591),
.B(n_1569),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1598),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1597),
.B(n_1578),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1605),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1616),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1635),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1632),
.B(n_1584),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1635),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1633),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1627),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1635),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1600),
.C(n_1599),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1626),
.A2(n_1600),
.B(n_1608),
.C(n_1606),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1627),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1640),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1645),
.B(n_1533),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1640),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1598),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1585),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1640),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1622),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1622),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1632),
.A2(n_1608),
.B1(n_1594),
.B2(n_1606),
.C(n_1599),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1646),
.B(n_1610),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1623),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1624),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1646),
.B(n_1583),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1634),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1633),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1646),
.B(n_1583),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1634),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1620),
.B(n_1596),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1623),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1636),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1637),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1637),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1620),
.B(n_1596),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1623),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1617),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1621),
.B(n_1583),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1648),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1675),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1654),
.B(n_1603),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1655),
.A2(n_1607),
.B(n_1582),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1660),
.B(n_1618),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1660),
.B(n_1618),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1669),
.A2(n_1609),
.B1(n_1607),
.B2(n_1565),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1660),
.B(n_1618),
.Y(n_1699)
);

OAI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1649),
.A2(n_1563),
.B(n_1619),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1674),
.B(n_1651),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1659),
.B(n_1492),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1663),
.B(n_1619),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1650),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.B(n_1665),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1625),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1677),
.B(n_1647),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1647),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1671),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1650),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1625),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1625),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1687),
.B(n_1628),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1663),
.B(n_1662),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1549),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1653),
.Y(n_1716)
);

NAND2x1_ASAP7_75t_L g1717 ( 
.A(n_1690),
.B(n_1617),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1662),
.B(n_1619),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1672),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1653),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1657),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1672),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1643),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1683),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1657),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1691),
.Y(n_1727)
);

OAI31xp33_ASAP7_75t_L g1728 ( 
.A1(n_1700),
.A2(n_1652),
.A3(n_1656),
.B(n_1658),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1694),
.B(n_1652),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1700),
.A2(n_1658),
.B1(n_1656),
.B2(n_1563),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1701),
.B(n_1670),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1693),
.A2(n_1681),
.B(n_1670),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1715),
.A2(n_1689),
.B(n_1681),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1717),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1698),
.A2(n_1505),
.B(n_1517),
.C(n_1492),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1721),
.A2(n_1594),
.B1(n_1581),
.B2(n_1555),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1628),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1721),
.A2(n_1513),
.B1(n_1621),
.B2(n_1631),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1702),
.A2(n_1717),
.B(n_1715),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1705),
.B(n_1643),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1714),
.A2(n_1513),
.B1(n_1705),
.B2(n_1692),
.Y(n_1741)
);

OAI32xp33_ASAP7_75t_L g1742 ( 
.A1(n_1714),
.A2(n_1689),
.A3(n_1631),
.B1(n_1630),
.B2(n_1638),
.Y(n_1742)
);

OAI322xp33_ASAP7_75t_L g1743 ( 
.A1(n_1703),
.A2(n_1638),
.A3(n_1680),
.B1(n_1686),
.B2(n_1685),
.C1(n_1684),
.C2(n_1667),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1691),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1695),
.A2(n_1563),
.B1(n_1513),
.B2(n_1581),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1692),
.B(n_1643),
.Y(n_1746)
);

OAI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1707),
.A2(n_1689),
.B1(n_1673),
.B2(n_1686),
.C(n_1685),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1697),
.Y(n_1748)
);

OAI32xp33_ASAP7_75t_L g1749 ( 
.A1(n_1703),
.A2(n_1630),
.A3(n_1638),
.B1(n_1684),
.B2(n_1680),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1695),
.B(n_1696),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1697),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

OAI321xp33_ASAP7_75t_L g1753 ( 
.A1(n_1729),
.A2(n_1715),
.A3(n_1718),
.B1(n_1699),
.B2(n_1696),
.C(n_1708),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1727),
.Y(n_1754)
);

AND2x4_ASAP7_75t_SL g1755 ( 
.A(n_1750),
.B(n_1715),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1735),
.A2(n_1715),
.B(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1731),
.Y(n_1757)
);

OAI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1732),
.A2(n_1699),
.B(n_1706),
.Y(n_1758)
);

OA21x2_ASAP7_75t_SL g1759 ( 
.A1(n_1737),
.A2(n_1617),
.B(n_1642),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1730),
.A2(n_1718),
.B1(n_1505),
.B2(n_1615),
.Y(n_1760)
);

OAI322xp33_ASAP7_75t_L g1761 ( 
.A1(n_1747),
.A2(n_1726),
.A3(n_1716),
.B1(n_1704),
.B2(n_1722),
.C1(n_1720),
.C2(n_1710),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1746),
.B(n_1724),
.Y(n_1762)
);

OAI32xp33_ASAP7_75t_L g1763 ( 
.A1(n_1733),
.A2(n_1712),
.A3(n_1706),
.B1(n_1711),
.B2(n_1724),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1740),
.B(n_1711),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1734),
.Y(n_1765)
);

AOI21xp33_ASAP7_75t_L g1766 ( 
.A1(n_1742),
.A2(n_1716),
.B(n_1710),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1744),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1748),
.Y(n_1768)
);

OAI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1738),
.A2(n_1712),
.B(n_1720),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1741),
.B(n_1644),
.Y(n_1770)
);

AOI211x1_ASAP7_75t_SL g1771 ( 
.A1(n_1735),
.A2(n_1725),
.B(n_1723),
.C(n_1719),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1751),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1739),
.A2(n_1726),
.B(n_1722),
.C(n_1723),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1757),
.B(n_1752),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1738),
.C(n_1741),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1765),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1767),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1758),
.B(n_1728),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1772),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1772),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1762),
.Y(n_1782)
);

AO22x1_ASAP7_75t_L g1783 ( 
.A1(n_1771),
.A2(n_1734),
.B1(n_1517),
.B2(n_1454),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1756),
.A2(n_1745),
.B1(n_1736),
.B2(n_1488),
.C(n_1454),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1775),
.B(n_1769),
.C(n_1753),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1776),
.B(n_1764),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_SL g1788 ( 
.A(n_1782),
.B(n_1445),
.Y(n_1788)
);

NAND5xp2_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1770),
.C(n_1768),
.D(n_1759),
.E(n_1755),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1785),
.A2(n_1760),
.B1(n_1768),
.B2(n_1630),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1782),
.B(n_1778),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1777),
.B(n_1763),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1780),
.A2(n_1749),
.B(n_1773),
.C(n_1743),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1777),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1774),
.B(n_1761),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1792),
.B(n_1781),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1783),
.B1(n_1760),
.B2(n_1785),
.C(n_1784),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1791),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1795),
.B(n_1666),
.Y(n_1799)
);

AO221x1_ASAP7_75t_L g1800 ( 
.A1(n_1790),
.A2(n_1630),
.B1(n_1723),
.B2(n_1719),
.C(n_1725),
.Y(n_1800)
);

AOI322xp5_ASAP7_75t_L g1801 ( 
.A1(n_1797),
.A2(n_1786),
.A3(n_1793),
.B1(n_1787),
.B2(n_1794),
.C1(n_1788),
.C2(n_1789),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1796),
.B(n_1666),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1799),
.Y(n_1803)
);

OAI322xp33_ASAP7_75t_L g1804 ( 
.A1(n_1798),
.A2(n_1800),
.A3(n_1725),
.B1(n_1719),
.B2(n_1661),
.C1(n_1664),
.C2(n_1679),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1796),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1797),
.A2(n_1529),
.B(n_1483),
.C(n_1502),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1805),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_SL g1808 ( 
.A(n_1802),
.B(n_1667),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1803),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1806),
.B(n_1668),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1804),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1809),
.B1(n_1807),
.B2(n_1810),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1808),
.A2(n_1801),
.B1(n_1498),
.B2(n_1630),
.C(n_1679),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1809),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1814),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1815),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1816),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1818),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1817),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1819),
.B(n_1812),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1820),
.A2(n_1813),
.B1(n_1549),
.B2(n_1664),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1668),
.B1(n_1676),
.B2(n_1673),
.C(n_1661),
.Y(n_1823)
);

AOI32xp33_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1821),
.A3(n_1676),
.B1(n_1683),
.B2(n_1688),
.Y(n_1824)
);

XNOR2xp5_ASAP7_75t_L g1825 ( 
.A(n_1824),
.B(n_1489),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_R g1826 ( 
.A1(n_1825),
.A2(n_1688),
.B1(n_1617),
.B2(n_1615),
.C(n_1642),
.Y(n_1826)
);

AOI211xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1524),
.B(n_1615),
.C(n_1522),
.Y(n_1827)
);


endmodule