module fake_jpeg_27225_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_28),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_55),
.B1(n_58),
.B2(n_47),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_42),
.B1(n_49),
.B2(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_60),
.B1(n_52),
.B2(n_51),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_96),
.B1(n_48),
.B2(n_45),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_93),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_0),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.C(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_57),
.B1(n_56),
.B2(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_1),
.Y(n_98)
);

INVx2_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_96),
.B1(n_83),
.B2(n_82),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_85),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_4),
.C(n_6),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_87),
.B1(n_91),
.B2(n_56),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_117),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_88),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_2),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_102),
.B(n_106),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_127),
.B(n_7),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_102),
.B1(n_92),
.B2(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_126),
.B1(n_131),
.B2(n_8),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_88),
.C(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_114),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_129),
.B1(n_123),
.B2(n_25),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_24),
.B(n_39),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_13),
.B(n_16),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_23),
.B(n_38),
.C(n_32),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_125),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_17),
.B1(n_27),
.B2(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_10),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_142),
.C(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_144),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_120),
.C(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_135),
.B(n_137),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);


endmodule