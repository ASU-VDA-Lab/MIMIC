module real_jpeg_27995_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_0),
.B(n_219),
.Y(n_224)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_37),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_37),
.B1(n_73),
.B2(n_74),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_4),
.A2(n_73),
.B1(n_74),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_4),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_106),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_106),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_106),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_43),
.Y(n_118)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_73),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_8),
.B(n_73),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_101),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_8),
.A2(n_10),
.B(n_23),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_29),
.B(n_32),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_45),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_131),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_130),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_108),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_80),
.B2(n_107),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_54),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_38),
.B(n_53),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_21),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_34),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_22),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_23),
.A2(n_26),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_23),
.A2(n_25),
.B(n_28),
.C(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_25),
.A2(n_41),
.B(n_184),
.C(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_25),
.B(n_90),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_25),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_27),
.B(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_27),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_31),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_33),
.A2(n_65),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_33),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_34),
.B(n_192),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B(n_48),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_41),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_40),
.B(n_77),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_45),
.B(n_50),
.C(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_41),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_44),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_44),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_45),
.B(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_47),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_48),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_49),
.B(n_146),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_57),
.A2(n_58),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_58),
.B(n_183),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_59),
.B(n_62),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_59),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_60),
.B(n_87),
.Y(n_119)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_63),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_64),
.A2(n_90),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_66),
.B(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_71),
.B(n_78),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_105),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_91),
.C(n_97),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_82),
.B(n_89),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_83),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_118),
.B(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_85),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_97),
.B1(n_98),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_95),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_115),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_113),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_115),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_126),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_116),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_119),
.B(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_121),
.B(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_126),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_265),
.B(n_270),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_177),
.B(n_253),
.C(n_264),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_165),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_134),
.B(n_165),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_147),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_136),
.B(n_137),
.C(n_147),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_143),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_158),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_149),
.B(n_154),
.C(n_158),
.Y(n_262)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_166),
.A2(n_167),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.C(n_175),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_252),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_245),
.B(n_251),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_203),
.B(n_244),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_181),
.B(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.C(n_189),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_200),
.C(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_239),
.B(n_243),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_220),
.B(n_238),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_206),
.B(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_216),
.C(n_217),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_237),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_225),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_241),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_259),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);


endmodule