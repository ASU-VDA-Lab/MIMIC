module fake_netlist_1_2554_n_690 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_690, n_647);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_690;
output n_647;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_24), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_39), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_18), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_19), .Y(n_85) );
BUFx10_ASAP7_75t_L g86 ( .A(n_51), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_57), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_16), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_63), .Y(n_90) );
BUFx8_ASAP7_75t_SL g91 ( .A(n_21), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_12), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_64), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_1), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_18), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_50), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_70), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_15), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_19), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_78), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_34), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_43), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_22), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_10), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_23), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_61), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_4), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_56), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_31), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_48), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_77), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_10), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_46), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_49), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_45), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_67), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_89), .B(n_0), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_83), .B(n_0), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_89), .B(n_1), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_96), .B(n_2), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_86), .B(n_4), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_112), .B(n_5), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_80), .B(n_5), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_107), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_125), .B(n_6), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_107), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_112), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_108), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_114), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_114), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_100), .B(n_7), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_86), .B(n_8), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_86), .B(n_8), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_85), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_117), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_123), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_123), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_84), .B(n_9), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
NOR2x1p5_ASAP7_75t_L g172 ( .A(n_142), .B(n_84), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_170), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_129), .B(n_127), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_131), .B(n_118), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_163), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_147), .B(n_98), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_131), .B(n_135), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_163), .B(n_95), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_164), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_135), .B(n_106), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_130), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_130), .Y(n_195) );
OR2x6_ASAP7_75t_L g196 ( .A(n_164), .B(n_111), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_153), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_130), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_154), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_154), .B(n_127), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_154), .B(n_128), .Y(n_208) );
OR2x6_ASAP7_75t_L g209 ( .A(n_145), .B(n_99), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_150), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_136), .B(n_103), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_136), .B(n_101), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_137), .B(n_92), .Y(n_214) );
INVx5_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_137), .A2(n_92), .B1(n_94), .B2(n_99), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
INVx5_ASAP7_75t_L g220 ( .A(n_165), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_150), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_138), .B(n_116), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_138), .B(n_97), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_140), .B(n_110), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_140), .B(n_115), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_153), .A2(n_116), .B1(n_110), .B2(n_94), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_144), .B(n_109), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_144), .B(n_111), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_148), .B(n_85), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_148), .B(n_122), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_153), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_149), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_134), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_178), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_210), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_218), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_183), .B(n_132), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_174), .A2(n_151), .B1(n_169), .B2(n_149), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_233), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_233), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_233), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_231), .B(n_152), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_232), .B(n_155), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_196), .B(n_156), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_233), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_174), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_231), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_229), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_183), .B(n_155), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_174), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_192), .B(n_156), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_190), .Y(n_256) );
BUFx8_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_173), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_202), .B(n_105), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_229), .Y(n_260) );
AND2x4_ASAP7_75t_SL g261 ( .A(n_178), .B(n_87), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_181), .B(n_151), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_229), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_202), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_176), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_196), .B(n_158), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_175), .B(n_157), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_174), .A2(n_157), .B1(n_169), .B2(n_160), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_207), .A2(n_162), .B1(n_160), .B2(n_167), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_172), .B(n_162), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_182), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_222), .B(n_158), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_209), .B(n_167), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_222), .B(n_166), .Y(n_279) );
NAND2xp33_ASAP7_75t_R g280 ( .A(n_209), .B(n_161), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_193), .B(n_166), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_186), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_212), .B(n_159), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_207), .A2(n_168), .B1(n_171), .B2(n_159), .Y(n_285) );
INVx5_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
BUFx12f_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_208), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_176), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_187), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_186), .B(n_171), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_223), .B(n_171), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_225), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_208), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_179), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_197), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_257), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_269), .A2(n_200), .B(n_205), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_248), .B(n_214), .Y(n_303) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_265), .B(n_120), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_198), .B1(n_179), .B2(n_191), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_234), .A2(n_198), .B(n_199), .C(n_203), .Y(n_306) );
CKINVDCx11_ASAP7_75t_R g307 ( .A(n_287), .Y(n_307) );
BUFx5_ASAP7_75t_L g308 ( .A(n_273), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_257), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_248), .B(n_228), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_255), .B(n_227), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_237), .Y(n_312) );
OAI22x1_ASAP7_75t_L g313 ( .A1(n_248), .A2(n_226), .B1(n_228), .B2(n_206), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_248), .B(n_228), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_255), .B(n_227), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_191), .B(n_189), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_243), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_267), .B(n_217), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
NOR2x1_ASAP7_75t_SL g322 ( .A(n_254), .B(n_213), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_257), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_267), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_237), .Y(n_327) );
OR2x6_ASAP7_75t_SL g328 ( .A(n_261), .B(n_102), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_295), .B(n_213), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_267), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_290), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_267), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_257), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_254), .B(n_230), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_295), .B(n_208), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_261), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_254), .A2(n_217), .B1(n_124), .B2(n_168), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_237), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_256), .B(n_208), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_SL g341 ( .A1(n_296), .A2(n_168), .B(n_134), .C(n_139), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_253), .B(n_208), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_253), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_261), .B(n_141), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_289), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_243), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_268), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_139), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_263), .B(n_143), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_268), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_278), .A2(n_85), .B1(n_143), .B2(n_141), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_247), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_328), .A2(n_287), .B1(n_280), .B2(n_273), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_239), .B(n_294), .C(n_262), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
BUFx12f_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_328), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_320), .B(n_247), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_336), .A2(n_273), .B1(n_288), .B2(n_297), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_319), .A2(n_314), .B1(n_310), .B2(n_342), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_343), .B(n_259), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_302), .A2(n_275), .B(n_281), .C(n_258), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_349), .Y(n_363) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_315), .A2(n_274), .B1(n_278), .B2(n_299), .C1(n_296), .C2(n_258), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_341), .A2(n_299), .B(n_275), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_310), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_307), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_310), .A2(n_241), .B1(n_272), .B2(n_270), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_312), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_349), .Y(n_370) );
INVx5_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_303), .B(n_319), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_314), .B(n_250), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_278), .B1(n_274), .B2(n_283), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_312), .Y(n_375) );
AO21x1_ASAP7_75t_L g376 ( .A1(n_334), .A2(n_281), .B(n_291), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_325), .A2(n_251), .B1(n_285), .B2(n_288), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_303), .A2(n_274), .B1(n_283), .B2(n_276), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_251), .B(n_266), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_338), .B(n_274), .Y(n_380) );
O2A1O1Ixp5_ASAP7_75t_SL g381 ( .A1(n_323), .A2(n_246), .B(n_240), .C(n_236), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_325), .B(n_291), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g384 ( .A1(n_316), .A2(n_282), .B(n_284), .C(n_236), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_357), .A2(n_313), .B1(n_333), .B2(n_324), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_304), .B(n_344), .C(n_306), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_380), .A2(n_305), .B1(n_244), .B2(n_240), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_313), .B1(n_332), .B2(n_330), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_373), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_333), .B1(n_324), .B2(n_309), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_371), .B(n_301), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_372), .B(n_244), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_361), .A2(n_345), .B1(n_351), .B2(n_348), .C(n_329), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_384), .B(n_341), .C(n_334), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_380), .A2(n_301), .B1(n_309), .B2(n_335), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_371), .B(n_323), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_352), .B(n_358), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_352), .A2(n_134), .B(n_264), .C(n_260), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_372), .B(n_329), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_378), .A2(n_292), .B(n_252), .C(n_260), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_360), .B(n_335), .Y(n_403) );
OAI22xp33_ASAP7_75t_SL g404 ( .A1(n_363), .A2(n_335), .B1(n_337), .B2(n_350), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_290), .B1(n_266), .B2(n_292), .Y(n_406) );
INVxp33_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_356), .A2(n_288), .B1(n_297), .B2(n_337), .Y(n_408) );
INVx5_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_252), .B(n_264), .C(n_85), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_356), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_367), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_409), .B(n_371), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_393), .B(n_384), .Y(n_415) );
OAI22xp5_ASAP7_75t_SL g416 ( .A1(n_412), .A2(n_367), .B1(n_371), .B2(n_374), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_399), .A2(n_368), .B1(n_362), .B2(n_347), .C(n_376), .Y(n_417) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_387), .B(n_375), .Y(n_418) );
INVx3_ASAP7_75t_SL g419 ( .A(n_413), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_386), .A2(n_362), .B1(n_382), .B2(n_359), .C(n_298), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_391), .A2(n_373), .B(n_377), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_393), .B(n_365), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_404), .A2(n_322), .B1(n_373), .B2(n_365), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_405), .B(n_365), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_388), .Y(n_426) );
INVx8_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_387), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_385), .B(n_381), .C(n_121), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_389), .A2(n_379), .B(n_297), .C(n_238), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_405), .B(n_298), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_389), .A2(n_271), .B1(n_238), .B2(n_331), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_388), .B(n_376), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_395), .B(n_195), .C(n_204), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_411), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_401), .B(n_323), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_276), .B1(n_298), .B2(n_235), .C(n_290), .Y(n_438) );
OAI222xp33_ASAP7_75t_L g439 ( .A1(n_396), .A2(n_331), .B1(n_271), .B2(n_91), .C1(n_13), .C2(n_14), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_395), .A2(n_346), .B(n_318), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_394), .A2(n_331), .B1(n_290), .B2(n_339), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_346), .B(n_326), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_409), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_435), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_422), .B(n_403), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_444), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_425), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_422), .B(n_397), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_417), .B(n_410), .C(n_409), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_424), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_443), .B(n_403), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_443), .B(n_390), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_415), .B(n_390), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_414), .B(n_404), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_424), .B(n_392), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_390), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_433), .A2(n_409), .B1(n_390), .B2(n_392), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_428), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_439), .A2(n_408), .A3(n_402), .B(n_392), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_447), .A2(n_400), .B1(n_398), .B2(n_406), .C(n_409), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_415), .A2(n_398), .B1(n_397), .B2(n_290), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_427), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_435), .B(n_397), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_437), .B(n_398), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_441), .A2(n_398), .B(n_339), .Y(n_473) );
AOI33xp33_ASAP7_75t_L g474 ( .A1(n_423), .A2(n_11), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_444), .B(n_339), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_433), .B(n_17), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_448), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_436), .B(n_17), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_20), .Y(n_479) );
AOI33xp33_ASAP7_75t_L g480 ( .A1(n_438), .A2(n_177), .A3(n_201), .B1(n_194), .B2(n_242), .B3(n_245), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_414), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_420), .B(n_177), .C(n_201), .D(n_194), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_431), .B(n_339), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_418), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_414), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_427), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_416), .A2(n_235), .B1(n_211), .B2(n_216), .C(n_242), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_427), .Y(n_489) );
AOI33xp33_ASAP7_75t_L g490 ( .A1(n_419), .A2(n_242), .A3(n_245), .B1(n_318), .B2(n_321), .B3(n_326), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_446), .B(n_25), .Y(n_491) );
AOI33xp33_ASAP7_75t_L g492 ( .A1(n_419), .A2(n_321), .A3(n_27), .B1(n_28), .B2(n_29), .B3(n_30), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_442), .B(n_327), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_421), .A2(n_327), .B1(n_312), .B2(n_235), .C1(n_237), .C2(n_243), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_427), .B(n_327), .Y(n_495) );
INVxp33_ASAP7_75t_SL g496 ( .A(n_432), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g498 ( .A(n_474), .B(n_429), .C(n_430), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_492), .B(n_418), .C(n_434), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_494), .B(n_312), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_456), .B(n_442), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_458), .B(n_440), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_452), .Y(n_503) );
AOI221x1_ASAP7_75t_L g504 ( .A1(n_482), .A2(n_185), .B1(n_195), .B2(n_204), .C(n_327), .Y(n_504) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_476), .B(n_440), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_449), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_464), .B(n_460), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_452), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_476), .B(n_440), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_450), .B(n_26), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_450), .B(n_33), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_478), .B(n_36), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_478), .B(n_37), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_453), .B(n_38), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_481), .B(n_42), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_457), .B(n_44), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_487), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_467), .B(n_235), .C(n_58), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_470), .B(n_286), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_453), .B(n_54), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_486), .B(n_59), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_472), .B(n_60), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_460), .B(n_62), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_496), .B(n_65), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_453), .B(n_66), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_457), .B(n_68), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_470), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_489), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_453), .B(n_69), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_455), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_455), .B(n_71), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_477), .B(n_73), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_472), .B(n_74), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_494), .B(n_308), .Y(n_536) );
NOR2xp33_ASAP7_75t_R g537 ( .A(n_495), .B(n_79), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_461), .B(n_249), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_466), .A2(n_286), .A3(n_250), .B(n_237), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_471), .B(n_185), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_462), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_463), .B(n_249), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_466), .A2(n_237), .B1(n_195), .B2(n_204), .C(n_185), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_490), .B(n_308), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_463), .B(n_249), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_471), .B(n_211), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_463), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_459), .B(n_249), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_451), .Y(n_550) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_464), .B(n_220), .C(n_215), .D(n_216), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_506), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
AOI21xp33_ASAP7_75t_L g554 ( .A1(n_539), .A2(n_454), .B(n_479), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_542), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_501), .B(n_465), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_541), .B(n_468), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_530), .B(n_485), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_524), .B(n_495), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_529), .B(n_485), .Y(n_560) );
OAI31xp33_ASAP7_75t_L g561 ( .A1(n_526), .A2(n_454), .A3(n_479), .B(n_484), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_526), .A2(n_482), .B(n_488), .C(n_483), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_548), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_550), .B(n_468), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_542), .B(n_485), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_550), .B(n_465), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_507), .B(n_485), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_507), .B(n_469), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_500), .A2(n_473), .B(n_493), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_503), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_503), .B(n_469), .Y(n_572) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_537), .B(n_491), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_505), .B(n_497), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_505), .B(n_512), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_513), .B(n_491), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_493), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_507), .B(n_493), .Y(n_579) );
AOI211x1_ASAP7_75t_L g580 ( .A1(n_500), .A2(n_480), .B(n_493), .C(n_497), .Y(n_580) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_504), .A2(n_497), .B(n_475), .Y(n_581) );
AND3x2_ASAP7_75t_L g582 ( .A(n_519), .B(n_475), .C(n_308), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_511), .B(n_475), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_537), .Y(n_584) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_509), .A2(n_475), .B(n_195), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_510), .B(n_185), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_525), .B(n_216), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_507), .B(n_243), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_536), .A2(n_286), .B1(n_250), .B2(n_249), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_511), .B(n_204), .Y(n_590) );
NAND2x1_ASAP7_75t_L g591 ( .A(n_524), .B(n_216), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_536), .B(n_215), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_551), .A2(n_250), .B(n_286), .C(n_215), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_525), .B(n_308), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_524), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_502), .B(n_308), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_533), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_512), .B(n_215), .Y(n_599) );
AOI211x1_ASAP7_75t_L g600 ( .A1(n_544), .A2(n_308), .B(n_220), .C(n_286), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_584), .A2(n_498), .B1(n_535), .B2(n_514), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_558), .B(n_531), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_567), .B(n_534), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_559), .A2(n_499), .B1(n_516), .B2(n_545), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_552), .B(n_528), .Y(n_606) );
NAND4xp25_ASAP7_75t_SL g607 ( .A(n_561), .B(n_531), .C(n_527), .D(n_521), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_553), .B(n_547), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_579), .B(n_527), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_563), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_556), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_561), .A2(n_535), .B(n_515), .C(n_521), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_580), .B(n_535), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_573), .A2(n_515), .B1(n_549), .B2(n_523), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_569), .A2(n_554), .B1(n_577), .B2(n_592), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_566), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_591), .A2(n_545), .B(n_549), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_555), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_555), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_557), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_575), .B(n_540), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_597), .B(n_540), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_571), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_598), .B(n_540), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
OR2x6_ASAP7_75t_L g627 ( .A(n_559), .B(n_522), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_576), .B(n_538), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_560), .B(n_517), .Y(n_629) );
AOI211x1_ASAP7_75t_L g630 ( .A1(n_554), .A2(n_543), .B(n_546), .C(n_520), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_568), .B(n_520), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_572), .B(n_220), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_569), .B(n_220), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_565), .B(n_250), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_565), .B(n_578), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_590), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_596), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_599), .Y(n_638) );
XOR2x2_ASAP7_75t_L g639 ( .A(n_582), .B(n_583), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_596), .B(n_595), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_588), .B(n_592), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_586), .Y(n_642) );
OA21x2_ASAP7_75t_SL g643 ( .A1(n_562), .A2(n_570), .B(n_600), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_585), .B(n_594), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_589), .A2(n_593), .B(n_587), .C(n_586), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_589), .B(n_585), .Y(n_646) );
UNKNOWN g647 ( );
INVx1_ASAP7_75t_L g648 ( .A(n_581), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_552), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_552), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_567), .A2(n_552), .B1(n_580), .B2(n_92), .C(n_99), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_567), .A2(n_552), .B1(n_580), .B2(n_92), .C(n_99), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_552), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_630), .B(n_651), .C(n_652), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_612), .A2(n_613), .B(n_605), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_644), .Y(n_657) );
AOI222xp33_ASAP7_75t_L g658 ( .A1(n_613), .A2(n_653), .B1(n_616), .B2(n_604), .C1(n_605), .C2(n_612), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_601), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_646), .A2(n_607), .B(n_618), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_615), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_633), .A2(n_604), .B(n_602), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_653), .A2(n_616), .B1(n_654), .B2(n_650), .C(n_649), .Y(n_663) );
OAI21xp33_ASAP7_75t_SL g664 ( .A1(n_620), .A2(n_619), .B(n_627), .Y(n_664) );
XNOR2x2_ASAP7_75t_L g665 ( .A(n_639), .B(n_643), .Y(n_665) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_614), .B(n_648), .C(n_606), .D(n_632), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_606), .A2(n_638), .B(n_641), .C(n_611), .Y(n_667) );
AOI31xp33_ASAP7_75t_L g668 ( .A1(n_638), .A2(n_645), .A3(n_636), .B(n_631), .Y(n_668) );
OAI211xp5_ASAP7_75t_L g669 ( .A1(n_656), .A2(n_622), .B(n_628), .C(n_637), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_656), .A2(n_617), .B1(n_626), .B2(n_621), .C(n_610), .Y(n_670) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_668), .B(n_627), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g672 ( .A1(n_664), .A2(n_603), .A3(n_609), .B1(n_635), .B2(n_640), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_660), .A2(n_667), .B1(n_666), .B2(n_663), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_658), .B(n_647), .C(n_634), .D(n_642), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_657), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_665), .B(n_623), .Y(n_676) );
OR4x1_ASAP7_75t_L g677 ( .A(n_673), .B(n_660), .C(n_655), .D(n_662), .Y(n_677) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_671), .B(n_669), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_670), .B(n_661), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_675), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_629), .B(n_625), .C(n_608), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_678), .B(n_674), .Y(n_682) );
AO22x2_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_672), .B1(n_659), .B2(n_624), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_680), .Y(n_684) );
INVx4_ASAP7_75t_L g685 ( .A(n_684), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_682), .B(n_679), .C(n_681), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_685), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_687), .B(n_686), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_688), .Y(n_689) );
AOI21xp33_ASAP7_75t_SL g690 ( .A1(n_689), .A2(n_683), .B(n_627), .Y(n_690) );
endmodule