module fake_jpeg_30035_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_21),
.B1(n_18),
.B2(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_55),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_63),
.B1(n_38),
.B2(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_67),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_32),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_31),
.CON(n_65),
.SN(n_65)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_44),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_39),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_77),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_30),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_79),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_80),
.B1(n_110),
.B2(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_29),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_109),
.B1(n_31),
.B2(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_95),
.Y(n_115)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g132 ( 
.A(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_16),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_27),
.B1(n_34),
.B2(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_34),
.B1(n_27),
.B2(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_33),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_37),
.B1(n_46),
.B2(n_25),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_40),
.B1(n_52),
.B2(n_45),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_106),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_19),
.B(n_23),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_46),
.B1(n_37),
.B2(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_40),
.B1(n_58),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_127),
.B1(n_136),
.B2(n_69),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_37),
.B1(n_25),
.B2(n_24),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_37),
.B1(n_24),
.B2(n_28),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_40),
.B(n_43),
.C(n_45),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_28),
.B1(n_35),
.B2(n_45),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_19),
.B(n_23),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_23),
.B(n_19),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_35),
.B1(n_34),
.B2(n_27),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_78),
.B1(n_103),
.B2(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_70),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_168),
.B1(n_113),
.B2(n_128),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_92),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_117),
.B1(n_123),
.B2(n_118),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_69),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_169),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_74),
.B(n_107),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_171),
.B(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_97),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_99),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_81),
.B1(n_71),
.B2(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_104),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_71),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_121),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_137),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_184),
.C(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_174),
.B(n_13),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_125),
.B1(n_116),
.B2(n_139),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_181),
.B1(n_188),
.B2(n_198),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_137),
.C(n_122),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_152),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_131),
.B(n_128),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_203),
.B(n_159),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_162),
.B1(n_167),
.B2(n_148),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_122),
.C(n_130),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_133),
.B1(n_86),
.B2(n_94),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_133),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_132),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_127),
.B1(n_126),
.B2(n_26),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_161),
.A2(n_111),
.B1(n_81),
.B2(n_87),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_204),
.B1(n_132),
.B2(n_2),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_76),
.B(n_101),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_26),
.B1(n_87),
.B2(n_109),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_43),
.C(n_45),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_155),
.B1(n_160),
.B2(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_210),
.B1(n_230),
.B2(n_231),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_170),
.B(n_171),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_209),
.A2(n_213),
.B(n_215),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_157),
.B1(n_168),
.B2(n_171),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_189),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_165),
.B(n_142),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_174),
.A2(n_168),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_221),
.C(n_186),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_155),
.C(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_233),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_133),
.B1(n_43),
.B2(n_132),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_R g228 ( 
.A1(n_191),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_43),
.B1(n_132),
.B2(n_40),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_175),
.B1(n_176),
.B2(n_181),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_189),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_12),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_210),
.B1(n_232),
.B2(n_219),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_248),
.B1(n_253),
.B2(n_258),
.Y(n_266)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_201),
.B1(n_196),
.B2(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_178),
.B1(n_199),
.B2(n_202),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_250),
.B1(n_227),
.B2(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_202),
.B1(n_199),
.B2(n_194),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_209),
.A2(n_196),
.B1(n_194),
.B2(n_184),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_192),
.C(n_13),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_10),
.C(n_8),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_215),
.A2(n_192),
.B1(n_12),
.B2(n_10),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_272),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_208),
.B1(n_225),
.B2(n_206),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_261),
.A2(n_273),
.B1(n_244),
.B2(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_265),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_216),
.B(n_221),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_279),
.B(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_220),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_257),
.B(n_241),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_244),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_278),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_222),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_248),
.A2(n_217),
.B1(n_229),
.B2(n_230),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_1),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_1),
.C(n_2),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_237),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_243),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_286),
.Y(n_298)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_261),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_254),
.C(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_5),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_256),
.B(n_2),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_296),
.B(n_276),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_4),
.C(n_5),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_272),
.C(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_262),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_259),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_286),
.B(n_288),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_273),
.C(n_5),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_291),
.B(n_287),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_295),
.B1(n_281),
.B2(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_289),
.B(n_292),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_316),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_306),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_293),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_298),
.B(n_301),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_312),
.B(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_300),
.C(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_318),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_331),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_317),
.B(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_324),
.B(n_321),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_330),
.B(n_324),
.C(n_310),
.D(n_293),
.Y(n_334)
);

FAx1_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_333),
.CI(n_6),
.CON(n_335),
.SN(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_6),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_7),
.B(n_260),
.C(n_290),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_7),
.Y(n_338)
);


endmodule