module fake_netlist_6_2032_n_2142 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2142);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2142;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_474;
wire n_527;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_38),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_10),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_45),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_55),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_80),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_124),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_50),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_190),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_137),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_40),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_87),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_26),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_165),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_77),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_111),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_107),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_55),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_112),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_145),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_37),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_88),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_134),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_159),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_15),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_119),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_51),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_152),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_179),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_103),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_129),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_96),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_34),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_15),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_35),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_29),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_93),
.Y(n_285)
);

INVx4_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_78),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_139),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_19),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_169),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_59),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_189),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_140),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_183),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_120),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_73),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_172),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_123),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_214),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_37),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_69),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_122),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_104),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_22),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_69),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_180),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_195),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_27),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_197),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_213),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_207),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_5),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_132),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_62),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_24),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_98),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_21),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_194),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_110),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_136),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_95),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_150),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_54),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_4),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_121),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_17),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_126),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_54),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_77),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_1),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_162),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_135),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_117),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_85),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_48),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_198),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_174),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_56),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_7),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_56),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_218),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_196),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_68),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_83),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_204),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_86),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_164),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_16),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_29),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_142),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_202),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_127),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_94),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_130),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_171),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_76),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_2),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_49),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_18),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_31),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_14),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_27),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_191),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_133),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_66),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_113),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_154),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_46),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_100),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_63),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_43),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_97),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_19),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_82),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_65),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_70),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_178),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_182),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_11),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_17),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_14),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_211),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_166),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_57),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_193),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_153),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_219),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_0),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_149),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_81),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_62),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_34),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_25),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_44),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_99),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_46),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_84),
.Y(n_411)
);

BUFx2_ASAP7_75t_SL g412 ( 
.A(n_49),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_65),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_61),
.Y(n_414)
);

BUFx8_ASAP7_75t_SL g415 ( 
.A(n_173),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_52),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_161),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_118),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_33),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_212),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_125),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_106),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_108),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_48),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_36),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_25),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_33),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_38),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_90),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_188),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_5),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_147),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_72),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_72),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_176),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_76),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_75),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_167),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_91),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_280),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_280),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_280),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_280),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_281),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_235),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_280),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_280),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_415),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_222),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_229),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_257),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_221),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_257),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_235),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_222),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_226),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_253),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_257),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_222),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_257),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_257),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_222),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_282),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_220),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_282),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_318),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_318),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_227),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_246),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_400),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_237),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_232),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_237),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_236),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_400),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_223),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_423),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_244),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_420),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_238),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_244),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_423),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_269),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_269),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_312),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_239),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_245),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_296),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_271),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_299),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_248),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_249),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_304),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_268),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_332),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_224),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_271),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_230),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_224),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_254),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_278),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_420),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_285),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_241),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_278),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_284),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_284),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_241),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_420),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_420),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_291),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_353),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_291),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_294),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_258),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_259),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_261),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_225),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_294),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_301),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_263),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_264),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_301),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_268),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_309),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_306),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_306),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_265),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_266),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_322),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_314),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_314),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_272),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_335),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_322),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_335),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_362),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_373),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_309),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_373),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_324),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_250),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_387),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_387),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_391),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_455),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_550),
.B(n_276),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_276),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_459),
.B(n_324),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_511),
.B(n_230),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_493),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_451),
.B(n_365),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_454),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_493),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_460),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_493),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_510),
.B(n_342),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_454),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_463),
.B(n_532),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_325),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_520),
.B(n_230),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_461),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_472),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_342),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_444),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_480),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_440),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_457),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_517),
.B(n_345),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_462),
.Y(n_589)
);

BUFx8_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_526),
.B(n_228),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_345),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_496),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_325),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_441),
.A2(n_283),
.B1(n_340),
.B2(n_337),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_485),
.B(n_309),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_273),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_498),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_482),
.B(n_270),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_466),
.B(n_433),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_445),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_483),
.B(n_465),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_488),
.B(n_315),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_465),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_445),
.B(n_289),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_501),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_446),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_449),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_450),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_450),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_485),
.B(n_230),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_503),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_452),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_448),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_494),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_466),
.B(n_290),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_471),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_452),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_504),
.B(n_433),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_495),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_550),
.B(n_312),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_499),
.B(n_376),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_550),
.B(n_292),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_504),
.B(n_297),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_507),
.B(n_247),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_479),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_500),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_481),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_481),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_448),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_512),
.B(n_302),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_512),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_303),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_508),
.B(n_247),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_516),
.B(n_486),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_467),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_489),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_458),
.B(n_437),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_545),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_490),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_566),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_588),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_584),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_566),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_610),
.Y(n_657)
);

BUFx4f_ASAP7_75t_L g658 ( 
.A(n_560),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_600),
.A2(n_490),
.B1(n_533),
.B2(n_426),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_603),
.B(n_607),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_584),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_610),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_598),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_613),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_456),
.C(n_447),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_615),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_583),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_561),
.B(n_523),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_561),
.B(n_524),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_629),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_573),
.B(n_412),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_596),
.A2(n_525),
.B1(n_530),
.B2(n_529),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_586),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_586),
.Y(n_678)
);

AO21x2_ASAP7_75t_L g679 ( 
.A1(n_622),
.A2(n_255),
.B(n_252),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_586),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_615),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_640),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_572),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_L g684 ( 
.A(n_645),
.B(n_537),
.C(n_536),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_591),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_562),
.B(n_541),
.C(n_443),
.Y(n_686)
);

AO22x2_ASAP7_75t_L g687 ( 
.A1(n_599),
.A2(n_437),
.B1(n_252),
.B2(n_256),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_630),
.B(n_533),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_640),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_591),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_473),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_629),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_582),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_561),
.B(n_506),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_567),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_591),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_588),
.B(n_506),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_600),
.B(n_547),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_606),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_559),
.B(n_275),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_458),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_629),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_651),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_587),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_588),
.B(n_601),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_633),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_620),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_612),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_588),
.B(n_305),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_633),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_612),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_573),
.B(n_310),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_629),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_SL g716 ( 
.A1(n_571),
.A2(n_255),
.B1(n_274),
.B2(n_256),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_612),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_587),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_589),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_614),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_567),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_589),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_592),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_592),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_614),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_573),
.B(n_320),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_569),
.B(n_275),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_577),
.B(n_275),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_580),
.B(n_231),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_614),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_609),
.B(n_326),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_583),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_560),
.B(n_312),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_617),
.A2(n_267),
.B1(n_379),
.B2(n_375),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_593),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_565),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_616),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_635),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_616),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_638),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_619),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_574),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_629),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_594),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_R g750 ( 
.A(n_621),
.B(n_502),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_626),
.B(n_399),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_619),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_629),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_624),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_636),
.B(n_399),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_568),
.Y(n_757)
);

INVxp33_ASAP7_75t_SL g758 ( 
.A(n_599),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_571),
.B(n_502),
.Y(n_759)
);

AOI21x1_ASAP7_75t_L g760 ( 
.A1(n_609),
.A2(n_277),
.B(n_274),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_608),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_624),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_608),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_568),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_629),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_638),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_624),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_568),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_568),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_598),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_639),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_639),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_637),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_590),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_598),
.A2(n_279),
.B1(n_321),
.B2(n_250),
.Y(n_775)
);

NOR2x1p5_ASAP7_75t_L g776 ( 
.A(n_627),
.B(n_233),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_590),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_543),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_564),
.Y(n_779)
);

INVx8_ASAP7_75t_L g780 ( 
.A(n_562),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_643),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_632),
.B(n_329),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_563),
.B(n_575),
.Y(n_783)
);

OA22x2_ASAP7_75t_L g784 ( 
.A1(n_649),
.A2(n_549),
.B1(n_543),
.B2(n_491),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_562),
.A2(n_279),
.B1(n_401),
.B2(n_321),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_604),
.B(n_549),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_637),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_564),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_574),
.B(n_399),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_604),
.B(n_467),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_604),
.B(n_469),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_648),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_642),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_564),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_570),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_648),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_625),
.B(n_277),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_642),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_560),
.B(n_312),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_634),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_622),
.A2(n_298),
.B1(n_300),
.B2(n_288),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_585),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_574),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_585),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_642),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_625),
.B(n_288),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_701),
.B(n_632),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_773),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_707),
.B(n_641),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_653),
.B(n_641),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_703),
.B(n_644),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_661),
.B(n_579),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_801),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_746),
.B(n_805),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_801),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_804),
.Y(n_819)
);

OR2x6_ASAP7_75t_SL g820 ( 
.A(n_739),
.B(n_234),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_746),
.B(n_644),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_805),
.B(n_631),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_692),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_773),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_780),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_716),
.A2(n_606),
.B(n_631),
.C(n_595),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_780),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_787),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_780),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_804),
.B(n_560),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_664),
.A2(n_579),
.B1(n_409),
.B2(n_421),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_682),
.B(n_689),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_664),
.B(n_649),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_770),
.B(n_425),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_770),
.B(n_806),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_780),
.A2(n_331),
.B1(n_333),
.B2(n_330),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_787),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_732),
.B(n_585),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_759),
.B(n_695),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_698),
.B(n_585),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_790),
.Y(n_841)
);

NAND3x1_ASAP7_75t_L g842 ( 
.A(n_783),
.B(n_300),
.C(n_298),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_679),
.A2(n_317),
.B1(n_319),
.B2(n_316),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_655),
.B(n_605),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_656),
.B(n_605),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_771),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_658),
.B(n_312),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_795),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_794),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_652),
.B(n_605),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_775),
.B(n_312),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_786),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_794),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_709),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_799),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_771),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_652),
.B(n_605),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_799),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_772),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_316),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_670),
.B(n_240),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_782),
.B(n_625),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_772),
.B(n_570),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_781),
.B(n_570),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_808),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_781),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_791),
.B(n_581),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_808),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_790),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_791),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_671),
.B(n_242),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_682),
.B(n_646),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_793),
.B(n_581),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_792),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_793),
.B(n_581),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_657),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_797),
.B(n_317),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_679),
.A2(n_319),
.B1(n_328),
.B2(n_323),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_689),
.B(n_646),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_797),
.B(n_708),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_727),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_712),
.B(n_323),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_663),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_663),
.Y(n_884)
);

OR2x2_ASAP7_75t_SL g885 ( 
.A(n_667),
.B(n_686),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_688),
.B(n_243),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_658),
.A2(n_409),
.B1(n_421),
.B2(n_401),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_665),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_709),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_674),
.A2(n_336),
.B1(n_347),
.B2(n_344),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_792),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_741),
.B(n_742),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_744),
.B(n_328),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_766),
.B(n_411),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_665),
.B(n_338),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_666),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_684),
.B(n_251),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_802),
.A2(n_338),
.B(n_356),
.C(n_343),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_666),
.B(n_343),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_683),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_705),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_668),
.B(n_356),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_750),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_683),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_690),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_668),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_711),
.A2(n_364),
.B1(n_389),
.B2(n_359),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_681),
.B(n_359),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_778),
.B(n_627),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_690),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_669),
.B(n_309),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_674),
.A2(n_352),
.B1(n_355),
.B2(n_348),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_681),
.B(n_364),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_SL g914 ( 
.A(n_676),
.B(n_411),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_766),
.B(n_411),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_694),
.Y(n_916)
);

NOR2x1p5_ASAP7_75t_L g917 ( 
.A(n_739),
.B(n_260),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_798),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_674),
.A2(n_358),
.B1(n_363),
.B2(n_357),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_694),
.B(n_389),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_798),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_736),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_700),
.B(n_396),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_674),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_789),
.B(n_262),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_798),
.B(n_396),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_745),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_700),
.B(n_706),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_766),
.B(n_411),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_706),
.B(n_439),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_718),
.B(n_439),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_745),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_675),
.B(n_590),
.C(n_293),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_672),
.B(n_411),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_718),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_719),
.B(n_628),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_752),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_785),
.B(n_411),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_L g939 ( 
.A(n_807),
.B(n_366),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_672),
.B(n_590),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_795),
.Y(n_941)
);

AOI22x1_ASAP7_75t_L g942 ( 
.A1(n_807),
.A2(n_809),
.B1(n_723),
.B2(n_724),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_SL g943 ( 
.A1(n_758),
.A2(n_380),
.B1(n_402),
.B2(n_611),
.Y(n_943)
);

BUFx6f_ASAP7_75t_SL g944 ( 
.A(n_778),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_809),
.A2(n_422),
.B1(n_378),
.B2(n_381),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_752),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_733),
.B(n_371),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_723),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_659),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_702),
.B(n_623),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_672),
.B(n_367),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_724),
.B(n_725),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_725),
.B(n_628),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_753),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_699),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_735),
.B(n_628),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_784),
.A2(n_384),
.B1(n_386),
.B2(n_390),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_753),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_784),
.B(n_809),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_735),
.B(n_738),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_755),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_738),
.B(n_647),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_748),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_728),
.B(n_394),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_729),
.B(n_287),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_693),
.B(n_398),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_751),
.B(n_295),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_679),
.A2(n_371),
.B1(n_431),
.B2(n_558),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_748),
.B(n_647),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_756),
.B(n_307),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_687),
.A2(n_431),
.B1(n_371),
.B2(n_558),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_749),
.B(n_311),
.C(n_308),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_755),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_749),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_762),
.Y(n_975)
);

AND2x6_ASAP7_75t_SL g976 ( 
.A(n_778),
.B(n_489),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_659),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_693),
.B(n_403),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_839),
.B(n_660),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_903),
.B(n_758),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_832),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_881),
.B(n_812),
.Y(n_982)
);

CKINVDCx8_ASAP7_75t_R g983 ( 
.A(n_976),
.Y(n_983)
);

OR2x2_ASAP7_75t_SL g984 ( 
.A(n_933),
.B(n_774),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_909),
.Y(n_985)
);

AND2x6_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_827),
.Y(n_986)
);

BUFx5_ASAP7_75t_L g987 ( 
.A(n_974),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_876),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_825),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_909),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_881),
.A2(n_763),
.B(n_761),
.C(n_779),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_847),
.A2(n_760),
.B(n_763),
.C(n_761),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_823),
.B(n_730),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_854),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_852),
.B(n_777),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_825),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_813),
.B(n_659),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_814),
.B(n_721),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_901),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_883),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_884),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_889),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_872),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_922),
.B(n_784),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_810),
.A2(n_800),
.B1(n_734),
.B2(n_721),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_884),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_909),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_821),
.A2(n_800),
.B1(n_734),
.B2(n_721),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_949),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_822),
.A2(n_861),
.B1(n_871),
.B2(n_918),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_825),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_862),
.B(n_722),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_957),
.B(n_327),
.C(n_313),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_888),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_924),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_817),
.B(n_722),
.Y(n_1017)
);

INVx3_ASAP7_75t_SL g1018 ( 
.A(n_885),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_817),
.B(n_816),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_879),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_826),
.A2(n_815),
.B(n_886),
.C(n_965),
.Y(n_1021)
);

AO22x1_ASAP7_75t_L g1022 ( 
.A1(n_965),
.A2(n_777),
.B1(n_334),
.B2(n_341),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_896),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_841),
.B(n_693),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_827),
.B(n_774),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_906),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_944),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_906),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_891),
.B(n_776),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_722),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_974),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_827),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_841),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_819),
.B(n_764),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_869),
.B(n_704),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_811),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_959),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_815),
.B(n_576),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_911),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_869),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_874),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_834),
.B(n_874),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_949),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_827),
.B(n_704),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_835),
.B(n_764),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_921),
.B(n_829),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_977),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_928),
.B(n_764),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_834),
.A2(n_687),
.B(n_346),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_830),
.A2(n_715),
.B(n_704),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_824),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_944),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_947),
.B(n_491),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_829),
.B(n_715),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_952),
.B(n_768),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_829),
.B(n_846),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_828),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_843),
.A2(n_687),
.B1(n_431),
.B2(n_371),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_840),
.A2(n_754),
.B(n_715),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_837),
.Y(n_1060)
);

AO22x1_ASAP7_75t_L g1061 ( 
.A1(n_967),
.A2(n_405),
.B1(n_370),
.B2(n_369),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_856),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_SL g1063 ( 
.A(n_831),
.B(n_349),
.C(n_339),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_837),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_926),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_843),
.A2(n_687),
.B1(n_431),
.B2(n_762),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_926),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_829),
.B(n_754),
.Y(n_1068)
);

NOR2x2_ASAP7_75t_L g1069 ( 
.A(n_943),
.B(n_705),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_833),
.B(n_597),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_848),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_960),
.B(n_768),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_859),
.Y(n_1073)
);

NOR2x2_ASAP7_75t_L g1074 ( 
.A(n_971),
.B(n_602),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_878),
.A2(n_938),
.B1(n_851),
.B2(n_887),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_917),
.B(n_618),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_977),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_880),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_866),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_955),
.B(n_650),
.Y(n_1080)
);

AND2x6_ASAP7_75t_L g1081 ( 
.A(n_870),
.B(n_768),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_900),
.B(n_492),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_904),
.B(n_492),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_905),
.B(n_910),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_916),
.B(n_769),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_935),
.B(n_497),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_967),
.B(n_399),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_948),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_963),
.B(n_497),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_863),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_882),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_925),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_864),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_867),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_848),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_873),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_925),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_875),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_878),
.B(n_769),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_851),
.A2(n_767),
.B1(n_429),
.B2(n_654),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_938),
.A2(n_767),
.B1(n_429),
.B2(n_654),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_968),
.A2(n_429),
.B1(n_662),
.B2(n_673),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_861),
.B(n_754),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_820),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_848),
.Y(n_1105)
);

CKINVDCx11_ASAP7_75t_R g1106 ( 
.A(n_907),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_849),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_940),
.B(n_676),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_893),
.Y(n_1109)
);

BUFx4f_ASAP7_75t_L g1110 ( 
.A(n_860),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_849),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_853),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_853),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_855),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_838),
.B(n_769),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_871),
.B(n_760),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_848),
.B(n_795),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_941),
.Y(n_1118)
);

BUFx4f_ASAP7_75t_L g1119 ( 
.A(n_860),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_897),
.A2(n_696),
.B1(n_757),
.B2(n_779),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_892),
.B(n_662),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_941),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_842),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_855),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_858),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_858),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_897),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_865),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_886),
.B(n_696),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_941),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_SL g1131 ( 
.A(n_964),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_970),
.B(n_676),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_L g1133 ( 
.A(n_941),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_877),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_865),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_972),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_868),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_970),
.B(n_696),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_868),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_962),
.B(n_969),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_898),
.A2(n_779),
.B(n_788),
.C(n_677),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_927),
.B(n_932),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_950),
.B(n_676),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_932),
.B(n_937),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_937),
.B(n_673),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_844),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_845),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_890),
.B(n_747),
.Y(n_1149)
);

OAI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_971),
.A2(n_351),
.B(n_350),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_946),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_954),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_912),
.B(n_505),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_968),
.A2(n_429),
.B1(n_677),
.B2(n_678),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_982),
.A2(n_847),
.B1(n_899),
.B2(n_895),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_989),
.B(n_940),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1092),
.B(n_919),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_982),
.B(n_894),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1092),
.B(n_894),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1075),
.A2(n_920),
.B1(n_931),
.B2(n_923),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1021),
.A2(n_915),
.B(n_929),
.C(n_945),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1078),
.B(n_915),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1050),
.A2(n_942),
.B(n_857),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1087),
.A2(n_836),
.B1(n_929),
.B2(n_939),
.Y(n_1164)
);

INVxp33_ASAP7_75t_SL g1165 ( 
.A(n_1025),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1078),
.B(n_902),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_997),
.A2(n_966),
.B(n_951),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1042),
.B(n_1020),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1097),
.B(n_908),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1011),
.A2(n_978),
.B1(n_966),
.B2(n_951),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1012),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1097),
.A2(n_913),
.B(n_930),
.C(n_978),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_997),
.A2(n_934),
.B(n_850),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1130),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_980),
.B(n_936),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1075),
.A2(n_1019),
.B1(n_1099),
.B2(n_1127),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_1116),
.A2(n_914),
.B(n_973),
.C(n_961),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_989),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1068),
.A2(n_765),
.B(n_747),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_SL g1180 ( 
.A1(n_979),
.A2(n_535),
.B(n_505),
.C(n_509),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1087),
.A2(n_956),
.B(n_953),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1019),
.B(n_954),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1134),
.B(n_958),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_994),
.B(n_958),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1012),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1091),
.B(n_961),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1001),
.Y(n_1187)
);

OAI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1018),
.A2(n_385),
.B1(n_388),
.B2(n_392),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1038),
.B(n_372),
.C(n_361),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1116),
.A2(n_975),
.B(n_973),
.C(n_788),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1109),
.B(n_975),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1020),
.B(n_374),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_998),
.B(n_795),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1038),
.B(n_377),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_R g1195 ( 
.A(n_1014),
.B(n_404),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1004),
.B(n_1018),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1133),
.A2(n_765),
.B(n_747),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1103),
.A2(n_765),
.B(n_747),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1070),
.A2(n_438),
.B1(n_417),
.B2(n_418),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1140),
.A2(n_803),
.B(n_796),
.Y(n_1200)
);

INVxp33_ASAP7_75t_SL g1201 ( 
.A(n_1025),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_L g1202 ( 
.A(n_985),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1005),
.A2(n_430),
.B(n_435),
.C(n_432),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1140),
.A2(n_803),
.B(n_796),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1023),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1039),
.A2(n_696),
.B1(n_757),
.B2(n_795),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1012),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1000),
.A2(n_382),
.B1(n_434),
.B2(n_427),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_1027),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_L g1210 ( 
.A(n_990),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1028),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1049),
.A2(n_535),
.B(n_534),
.C(n_531),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_SL g1213 ( 
.A1(n_983),
.A2(n_383),
.B1(n_424),
.B2(n_419),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1099),
.A2(n_513),
.B(n_509),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_987),
.B(n_757),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_988),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_1053),
.B(n_92),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_999),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1005),
.A2(n_796),
.B1(n_757),
.B2(n_691),
.Y(n_1219)
);

OAI21xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1084),
.A2(n_552),
.B(n_513),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1084),
.A2(n_531),
.B(n_528),
.C(n_527),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1006),
.A2(n_685),
.B1(n_743),
.B2(n_740),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1150),
.A2(n_406),
.B(n_393),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1052),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1138),
.A2(n_697),
.B(n_743),
.C(n_740),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1050),
.A2(n_713),
.B(n_737),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_993),
.A2(n_522),
.B(n_521),
.C(n_519),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1080),
.B(n_395),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1033),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_995),
.B(n_1029),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1058),
.A2(n_1066),
.B1(n_998),
.B2(n_1110),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1058),
.A2(n_408),
.B1(n_410),
.B2(n_413),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1041),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1090),
.B(n_678),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1138),
.A2(n_710),
.B(n_737),
.C(n_731),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_984),
.A2(n_414),
.B1(n_397),
.B2(n_416),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1093),
.B(n_680),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1094),
.B(n_680),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_991),
.A2(n_515),
.B(n_514),
.C(n_557),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1096),
.B(n_1098),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1040),
.A2(n_515),
.B(n_514),
.C(n_557),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1062),
.A2(n_546),
.B(n_556),
.C(n_555),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_981),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1137),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1129),
.A2(n_685),
.B(n_731),
.C(n_726),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1066),
.A2(n_544),
.B1(n_519),
.B2(n_521),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1032),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1032),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1071),
.A2(n_803),
.B(n_726),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1104),
.A2(n_540),
.B1(n_555),
.B2(n_554),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1065),
.B(n_527),
.Y(n_1251)
);

OAI22x1_ASAP7_75t_L g1252 ( 
.A1(n_1123),
.A2(n_540),
.B1(n_554),
.B2(n_553),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_SL g1253 ( 
.A(n_1110),
.B(n_528),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1073),
.B(n_691),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1122),
.A2(n_720),
.B(n_717),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1016),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1032),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1037),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1008),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1119),
.A2(n_544),
.B1(n_534),
.B2(n_539),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1079),
.A2(n_546),
.B(n_539),
.C(n_542),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1132),
.A2(n_713),
.B(n_710),
.C(n_697),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1031),
.B(n_1),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1088),
.B(n_1082),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1037),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1137),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1002),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1136),
.B(n_3),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1007),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1082),
.B(n_542),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1095),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_989),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1014),
.A2(n_551),
.B(n_548),
.C(n_477),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1122),
.A2(n_551),
.B(n_548),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1083),
.B(n_469),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1003),
.B(n_4),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1153),
.B(n_6),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1131),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1083),
.A2(n_477),
.B(n_476),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1086),
.B(n_470),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1089),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1095),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_987),
.B(n_1067),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1013),
.B(n_470),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1013),
.B(n_474),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1106),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_987),
.B(n_286),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1129),
.A2(n_286),
.B(n_9),
.C(n_11),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_996),
.A2(n_217),
.B(n_210),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_996),
.A2(n_201),
.B(n_200),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1121),
.B(n_8),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1119),
.A2(n_1063),
.B(n_992),
.C(n_1009),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1074),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_987),
.B(n_192),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1015),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1076),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1010),
.B(n_186),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1017),
.A2(n_185),
.B1(n_184),
.B2(n_181),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_996),
.A2(n_177),
.B(n_175),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1059),
.A2(n_170),
.B(n_168),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1063),
.A2(n_13),
.B(n_20),
.C(n_21),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1026),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_986),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1167),
.A2(n_1115),
.B(n_1048),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1194),
.B(n_1022),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1224),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1164),
.A2(n_992),
.B(n_1121),
.C(n_1056),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1240),
.B(n_987),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1228),
.A2(n_1056),
.B(n_1017),
.C(n_1055),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1226),
.A2(n_1146),
.B(n_1108),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1258),
.B(n_1046),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1231),
.A2(n_1102),
.B1(n_1154),
.B2(n_1101),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_SL g1314 ( 
.A1(n_1170),
.A2(n_1125),
.B(n_1152),
.C(n_1151),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1175),
.B(n_1176),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1158),
.B(n_987),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1161),
.A2(n_1048),
.B(n_1072),
.C(n_1055),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_1168),
.Y(n_1319)
);

OR2x6_ASAP7_75t_L g1320 ( 
.A(n_1265),
.B(n_1046),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1182),
.B(n_1072),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1159),
.A2(n_1045),
.B(n_1030),
.C(n_1034),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1160),
.A2(n_1115),
.B(n_1059),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1163),
.A2(n_1146),
.B(n_1108),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1160),
.A2(n_1054),
.B(n_1044),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1155),
.A2(n_1173),
.B(n_1172),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1155),
.A2(n_1045),
.B(n_1149),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1166),
.B(n_1147),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1222),
.A2(n_1145),
.B(n_1142),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_SL g1330 ( 
.A(n_1268),
.B(n_1154),
.C(n_1102),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1209),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1232),
.A2(n_1101),
.B1(n_1100),
.B2(n_1030),
.C(n_1034),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1282),
.B(n_1046),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1162),
.B(n_1147),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1200),
.A2(n_1142),
.B(n_1145),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1285),
.B(n_1147),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1190),
.A2(n_1293),
.B(n_1235),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1229),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1157),
.A2(n_1085),
.B(n_1035),
.C(n_1024),
.Y(n_1339)
);

NOR4xp25_ASAP7_75t_L g1340 ( 
.A(n_1302),
.B(n_1141),
.C(n_1100),
.D(n_1085),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1259),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1218),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1165),
.A2(n_1061),
.B1(n_1081),
.B2(n_1148),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_1196),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1286),
.B(n_1148),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1178),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1205),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1259),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1287),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1201),
.B(n_1148),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_SL g1351 ( 
.A(n_1189),
.B(n_1120),
.C(n_1069),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1288),
.A2(n_1139),
.B(n_1111),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1211),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1296),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1214),
.A2(n_1180),
.B(n_1225),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1192),
.B(n_1294),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1245),
.A2(n_1113),
.B(n_1114),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1233),
.Y(n_1358)
);

AOI31xp67_ASAP7_75t_L g1359 ( 
.A1(n_1193),
.A2(n_1295),
.A3(n_1215),
.B(n_1292),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1230),
.B(n_1010),
.Y(n_1360)
);

AO32x2_ASAP7_75t_L g1361 ( 
.A1(n_1231),
.A2(n_1135),
.A3(n_1118),
.B1(n_1126),
.B2(n_1124),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1169),
.B(n_1043),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1204),
.A2(n_1144),
.B(n_1036),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1301),
.A2(n_1051),
.B(n_1060),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1243),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1304),
.B(n_1095),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_SL g1368 ( 
.A(n_1178),
.B(n_1105),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1281),
.B(n_1043),
.Y(n_1369)
);

CKINVDCx6p67_ASAP7_75t_R g1370 ( 
.A(n_1174),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1181),
.A2(n_1118),
.B(n_1105),
.Y(n_1371)
);

AOI211x1_ASAP7_75t_L g1372 ( 
.A1(n_1264),
.A2(n_1143),
.B(n_22),
.C(n_23),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1289),
.A2(n_1047),
.B(n_1077),
.C(n_1064),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1220),
.A2(n_1239),
.B(n_1237),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1255),
.A2(n_1128),
.B(n_1057),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1272),
.A2(n_986),
.B(n_1112),
.Y(n_1376)
);

INVx3_ASAP7_75t_SL g1377 ( 
.A(n_1278),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1253),
.A2(n_986),
.B(n_1107),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1277),
.B(n_1232),
.C(n_1199),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1177),
.A2(n_986),
.B(n_1117),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1156),
.A2(n_986),
.B(n_1081),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_1117),
.B(n_1081),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1234),
.B(n_1081),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1284),
.A2(n_1117),
.B(n_1081),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1256),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1238),
.A2(n_1117),
.B(n_163),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1183),
.B(n_1117),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1217),
.A2(n_1270),
.B1(n_1191),
.B2(n_1186),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1198),
.A2(n_160),
.B(n_155),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1267),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1203),
.A2(n_1223),
.B(n_1212),
.C(n_1263),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1219),
.A2(n_24),
.B1(n_28),
.B2(n_30),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1275),
.A2(n_32),
.B(n_35),
.C(n_39),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1269),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1298),
.B(n_39),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1185),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1303),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1233),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1283),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1290),
.A2(n_131),
.B(n_128),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1280),
.A2(n_1221),
.B(n_1279),
.C(n_1273),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1174),
.B(n_105),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1251),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1251),
.B(n_40),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1202),
.B(n_41),
.Y(n_1405)
);

INVx3_ASAP7_75t_SL g1406 ( 
.A(n_1184),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1254),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1252),
.B(n_41),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1262),
.A2(n_102),
.B(n_101),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1299),
.A2(n_42),
.B(n_43),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1179),
.A2(n_42),
.B(n_45),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1244),
.B(n_47),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1171),
.B(n_47),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1185),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1208),
.B(n_52),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1184),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1266),
.Y(n_1417)
);

OR2x2_ASAP7_75t_SL g1418 ( 
.A(n_1202),
.B(n_53),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1291),
.A2(n_58),
.B(n_59),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1300),
.A2(n_60),
.B(n_61),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1206),
.A2(n_60),
.B(n_63),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1271),
.B(n_64),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1260),
.A2(n_67),
.B(n_68),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1246),
.A2(n_1260),
.B1(n_1184),
.B2(n_1276),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1227),
.A2(n_67),
.B(n_70),
.C(n_71),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1210),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1197),
.A2(n_71),
.B(n_73),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1248),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1248),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_L g1430 ( 
.A(n_1171),
.B(n_74),
.Y(n_1430)
);

INVx5_ASAP7_75t_L g1431 ( 
.A(n_1283),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1241),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1271),
.B(n_1207),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1207),
.B(n_78),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1247),
.B(n_79),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1210),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1274),
.A2(n_1261),
.B(n_1242),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1257),
.A2(n_1246),
.B(n_1283),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1257),
.A2(n_1195),
.B(n_1297),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1188),
.B(n_1236),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1250),
.A2(n_1226),
.B(n_1163),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1213),
.B(n_1194),
.C(n_1087),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1226),
.A2(n_1163),
.B(n_1173),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1240),
.B(n_982),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1167),
.A2(n_982),
.B(n_658),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1233),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1161),
.A2(n_1021),
.B(n_982),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1194),
.A2(n_1021),
.B(n_982),
.C(n_1092),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1170),
.A2(n_1116),
.A3(n_1190),
.B(n_1293),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1161),
.A2(n_1021),
.B(n_982),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1170),
.A2(n_1116),
.A3(n_1190),
.B(n_1293),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_SL g1452 ( 
.A(n_1194),
.B(n_1087),
.C(n_739),
.Y(n_1452)
);

OAI22x1_ASAP7_75t_L g1453 ( 
.A1(n_1194),
.A2(n_1018),
.B1(n_1097),
.B2(n_1092),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1226),
.A2(n_1163),
.B(n_1173),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1194),
.B(n_980),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1161),
.A2(n_1021),
.B(n_982),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1240),
.A2(n_1301),
.B(n_1302),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1229),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_L g1459 ( 
.A(n_1194),
.B(n_1087),
.C(n_661),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1167),
.A2(n_982),
.B(n_658),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1168),
.B(n_1070),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1240),
.B(n_982),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1185),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1209),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1226),
.A2(n_1163),
.B(n_1173),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1317),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_L g1467 ( 
.A(n_1448),
.B(n_1316),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1458),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1326),
.A2(n_1454),
.B(n_1443),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1455),
.B(n_1459),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1380),
.A2(n_1460),
.B(n_1445),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1447),
.A2(n_1456),
.B(n_1450),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1444),
.B(n_1462),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1447),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1450),
.A2(n_1456),
.B(n_1305),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1315),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1441),
.A2(n_1465),
.B(n_1324),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1330),
.A2(n_1442),
.B1(n_1379),
.B2(n_1306),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1461),
.B(n_1319),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1391),
.A2(n_1310),
.B(n_1316),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1311),
.A2(n_1335),
.B(n_1364),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1365),
.A2(n_1329),
.B(n_1305),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1431),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1347),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1367),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1401),
.A2(n_1452),
.B(n_1410),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1334),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1349),
.Y(n_1489)
);

INVx8_ASAP7_75t_L g1490 ( 
.A(n_1431),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1307),
.B(n_1366),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1444),
.A2(n_1462),
.B1(n_1343),
.B2(n_1328),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1352),
.A2(n_1327),
.B(n_1382),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1355),
.A2(n_1375),
.B(n_1325),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1431),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1368),
.B(n_1431),
.Y(n_1496)
);

O2A1O1Ixp5_ASAP7_75t_L g1497 ( 
.A1(n_1410),
.A2(n_1313),
.B(n_1355),
.C(n_1374),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1328),
.B(n_1356),
.Y(n_1498)
);

AO31x2_ASAP7_75t_L g1499 ( 
.A1(n_1313),
.A2(n_1308),
.A3(n_1318),
.B(n_1322),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1357),
.A2(n_1376),
.B(n_1411),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1428),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1398),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1342),
.B(n_1338),
.Y(n_1504)
);

OAI222xp33_ASAP7_75t_L g1505 ( 
.A1(n_1415),
.A2(n_1424),
.B1(n_1392),
.B2(n_1423),
.C1(n_1404),
.C2(n_1405),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1374),
.A2(n_1332),
.B(n_1357),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1423),
.A2(n_1424),
.B1(n_1392),
.B2(n_1395),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1363),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1371),
.A2(n_1384),
.B(n_1314),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1457),
.A2(n_1420),
.B(n_1421),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1381),
.B(n_1320),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_SL g1512 ( 
.A1(n_1419),
.A2(n_1373),
.B(n_1400),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1367),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1402),
.A2(n_1440),
.B1(n_1403),
.B2(n_1336),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1358),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1407),
.B(n_1369),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1446),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1393),
.A2(n_1425),
.B(n_1309),
.C(n_1427),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1339),
.A2(n_1388),
.B(n_1437),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1351),
.A2(n_1440),
.B1(n_1453),
.B2(n_1350),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1386),
.A2(n_1438),
.B(n_1389),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1333),
.A2(n_1436),
.B1(n_1426),
.B2(n_1360),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1344),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1390),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1394),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1437),
.A2(n_1321),
.B(n_1383),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1385),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1321),
.A2(n_1432),
.B(n_1345),
.C(n_1336),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_SL g1530 ( 
.A1(n_1383),
.A2(n_1387),
.B(n_1345),
.C(n_1388),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1397),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1333),
.B(n_1417),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1378),
.B(n_1439),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1435),
.A2(n_1416),
.B1(n_1406),
.B2(n_1408),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1435),
.B(n_1354),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1337),
.A2(n_1387),
.B(n_1362),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1337),
.Y(n_1537)
);

CKINVDCx6p67_ASAP7_75t_R g1538 ( 
.A(n_1331),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1464),
.Y(n_1539)
);

OAI222xp33_ASAP7_75t_L g1540 ( 
.A1(n_1422),
.A2(n_1434),
.B1(n_1412),
.B2(n_1433),
.C1(n_1418),
.C2(n_1429),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1361),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1361),
.A2(n_1451),
.B(n_1449),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1413),
.A2(n_1430),
.B1(n_1344),
.B2(n_1341),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1346),
.B(n_1463),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1370),
.A2(n_1377),
.B1(n_1348),
.B2(n_1399),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1340),
.A2(n_1359),
.B(n_1346),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1361),
.Y(n_1547)
);

BUFx2_ASAP7_75t_R g1548 ( 
.A(n_1409),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1396),
.A2(n_1414),
.B(n_1409),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1463),
.B(n_1449),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1372),
.B(n_1451),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1368),
.B(n_1431),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1331),
.Y(n_1555)
);

AO22x2_ASAP7_75t_L g1556 ( 
.A1(n_1313),
.A2(n_1330),
.B1(n_1424),
.B2(n_1459),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1455),
.A2(n_1021),
.B(n_1194),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1353),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1353),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1353),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1353),
.Y(n_1562)
);

AO31x2_ASAP7_75t_L g1563 ( 
.A1(n_1326),
.A2(n_1313),
.A3(n_1323),
.B(n_1327),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1353),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1455),
.A2(n_1021),
.B(n_1194),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1455),
.B(n_982),
.Y(n_1566)
);

INVx3_ASAP7_75t_SL g1567 ( 
.A(n_1307),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1455),
.A2(n_1330),
.B1(n_1442),
.B2(n_1379),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1326),
.A2(n_1450),
.B(n_1447),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1368),
.B(n_1431),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1455),
.A2(n_1330),
.B1(n_1442),
.B2(n_1379),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1455),
.A2(n_1087),
.B1(n_982),
.B2(n_1442),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1574)
);

AOI22x1_ASAP7_75t_L g1575 ( 
.A1(n_1453),
.A2(n_1326),
.B1(n_1410),
.B2(n_1457),
.Y(n_1575)
);

BUFx8_ASAP7_75t_SL g1576 ( 
.A(n_1341),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1368),
.B(n_1431),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1455),
.A2(n_1330),
.B1(n_1442),
.B2(n_1379),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1455),
.A2(n_982),
.B1(n_1462),
.B2(n_1444),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1326),
.A2(n_1454),
.B(n_1443),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1331),
.Y(n_1584)
);

AO31x2_ASAP7_75t_L g1585 ( 
.A1(n_1326),
.A2(n_1313),
.A3(n_1323),
.B(n_1327),
.Y(n_1585)
);

AO21x2_ASAP7_75t_L g1586 ( 
.A1(n_1326),
.A2(n_1450),
.B(n_1447),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_SL g1588 ( 
.A1(n_1410),
.A2(n_1457),
.B(n_1419),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1326),
.A2(n_1454),
.B(n_1443),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1455),
.A2(n_982),
.B1(n_1462),
.B2(n_1444),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_SL g1591 ( 
.A1(n_1410),
.A2(n_1457),
.B(n_1419),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1455),
.A2(n_1021),
.B(n_1194),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1461),
.B(n_1168),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1455),
.A2(n_1330),
.B1(n_1442),
.B2(n_1379),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1455),
.A2(n_1021),
.B(n_1194),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_SL g1596 ( 
.A1(n_1410),
.A2(n_1457),
.B(n_1419),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1446),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1455),
.A2(n_982),
.B(n_1450),
.C(n_1447),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1455),
.A2(n_1330),
.B1(n_1442),
.B2(n_1379),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1461),
.B(n_1168),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1331),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1331),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_SL g1603 ( 
.A1(n_1410),
.A2(n_1457),
.B(n_1419),
.Y(n_1603)
);

INVx8_ASAP7_75t_L g1604 ( 
.A(n_1431),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1455),
.A2(n_1087),
.B1(n_982),
.B2(n_1442),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1367),
.Y(n_1606)
);

AO31x2_ASAP7_75t_L g1607 ( 
.A1(n_1326),
.A2(n_1313),
.A3(n_1323),
.B(n_1327),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1459),
.B(n_1455),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1455),
.B(n_982),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1326),
.A2(n_1450),
.B(n_1447),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1461),
.B(n_1168),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1455),
.A2(n_982),
.B(n_1450),
.C(n_1447),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1319),
.B(n_1461),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1441),
.A2(n_1454),
.B(n_1443),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1455),
.A2(n_1087),
.B1(n_1442),
.B2(n_600),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1459),
.B(n_1455),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1461),
.B(n_1168),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1331),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1319),
.B(n_1461),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1468),
.Y(n_1622)
);

OA22x2_ASAP7_75t_L g1623 ( 
.A1(n_1521),
.A2(n_1487),
.B1(n_1565),
.B2(n_1557),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1488),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1488),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1617),
.A2(n_1566),
.B1(n_1609),
.B2(n_1572),
.Y(n_1627)
);

NOR2xp67_ASAP7_75t_L g1628 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1497),
.A2(n_1483),
.B(n_1520),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1613),
.B(n_1619),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1569),
.A2(n_1572),
.B1(n_1594),
.B2(n_1580),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1466),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1468),
.Y(n_1633)
);

O2A1O1Ixp5_ASAP7_75t_L g1634 ( 
.A1(n_1592),
.A2(n_1595),
.B(n_1481),
.C(n_1476),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1473),
.A2(n_1614),
.B(n_1598),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1498),
.B(n_1535),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1546),
.A2(n_1494),
.B(n_1509),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1569),
.A2(n_1594),
.B1(n_1599),
.B2(n_1580),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_SL g1641 ( 
.A1(n_1517),
.A2(n_1474),
.B(n_1502),
.Y(n_1641)
);

BUFx12f_ASAP7_75t_L g1642 ( 
.A(n_1489),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1502),
.B(n_1514),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1471),
.B(n_1599),
.Y(n_1644)
);

OA22x2_ASAP7_75t_L g1645 ( 
.A1(n_1534),
.A2(n_1523),
.B1(n_1618),
.B2(n_1608),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1471),
.B(n_1608),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1479),
.A2(n_1507),
.B1(n_1605),
.B2(n_1573),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1568),
.B(n_1578),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1568),
.B(n_1578),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1573),
.A2(n_1605),
.B1(n_1505),
.B2(n_1556),
.C(n_1479),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1477),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1507),
.A2(n_1543),
.B1(n_1614),
.B2(n_1598),
.Y(n_1652)
);

INVx3_ASAP7_75t_SL g1653 ( 
.A(n_1555),
.Y(n_1653)
);

NOR2xp67_ASAP7_75t_L g1654 ( 
.A(n_1545),
.B(n_1470),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1532),
.B(n_1618),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1489),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1467),
.A2(n_1540),
.B(n_1519),
.C(n_1529),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1556),
.A2(n_1467),
.B1(n_1475),
.B2(n_1515),
.C(n_1492),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1532),
.B(n_1561),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1562),
.B(n_1564),
.Y(n_1661)
);

AOI31xp33_ASAP7_75t_L g1662 ( 
.A1(n_1543),
.A2(n_1515),
.A3(n_1555),
.B(n_1602),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1528),
.A2(n_1556),
.B1(n_1597),
.B2(n_1518),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1503),
.A2(n_1475),
.B1(n_1575),
.B2(n_1548),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_SL g1665 ( 
.A(n_1511),
.B(n_1533),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1503),
.Y(n_1666)
);

OA21x2_ASAP7_75t_L g1667 ( 
.A1(n_1482),
.A2(n_1493),
.B(n_1478),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1496),
.A2(n_1553),
.B(n_1579),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1570),
.A2(n_1612),
.B(n_1586),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1504),
.A2(n_1529),
.B1(n_1519),
.B2(n_1491),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1496),
.A2(n_1571),
.B(n_1579),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1567),
.Y(n_1672)
);

O2A1O1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1588),
.A2(n_1596),
.B(n_1591),
.C(n_1603),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1511),
.A2(n_1513),
.B1(n_1606),
.B2(n_1486),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1530),
.A2(n_1506),
.B(n_1522),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1508),
.B(n_1525),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1501),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1512),
.A2(n_1485),
.B1(n_1531),
.B2(n_1526),
.C(n_1537),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1500),
.A2(n_1499),
.B(n_1604),
.C(n_1490),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1574),
.A2(n_1581),
.B(n_1610),
.Y(n_1680)
);

CKINVDCx14_ASAP7_75t_R g1681 ( 
.A(n_1539),
.Y(n_1681)
);

OA22x2_ASAP7_75t_L g1682 ( 
.A1(n_1551),
.A2(n_1533),
.B1(n_1602),
.B2(n_1549),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1527),
.B(n_1499),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1536),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1527),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1567),
.B(n_1533),
.Y(n_1687)
);

O2A1O1Ixp5_ASAP7_75t_L g1688 ( 
.A1(n_1472),
.A2(n_1541),
.B(n_1547),
.C(n_1585),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1499),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1499),
.A2(n_1547),
.B1(n_1541),
.B2(n_1539),
.C(n_1584),
.Y(n_1690)
);

NOR2xp67_ASAP7_75t_L g1691 ( 
.A(n_1484),
.B(n_1495),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1484),
.A2(n_1495),
.B(n_1490),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1510),
.A2(n_1620),
.B(n_1601),
.C(n_1584),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1510),
.A2(n_1620),
.B(n_1601),
.C(n_1542),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1510),
.B(n_1469),
.C(n_1589),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1538),
.A2(n_1604),
.B1(n_1490),
.B2(n_1542),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1604),
.A2(n_1542),
.B1(n_1583),
.B2(n_1469),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1552),
.A2(n_1616),
.B(n_1587),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1563),
.B(n_1585),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1585),
.B(n_1607),
.Y(n_1700)
);

AOI21x1_ASAP7_75t_SL g1701 ( 
.A1(n_1607),
.A2(n_1554),
.B(n_1559),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1577),
.A2(n_1611),
.B(n_1607),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1576),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1576),
.B(n_1480),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1617),
.A2(n_1455),
.B1(n_1442),
.B2(n_1566),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1569),
.A2(n_1580),
.B(n_1594),
.C(n_1572),
.Y(n_1706)
);

AND2x6_ASAP7_75t_L g1707 ( 
.A(n_1550),
.B(n_1537),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1557),
.B(n_1455),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1557),
.B(n_1455),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_SL g1710 ( 
.A(n_1511),
.B(n_1533),
.Y(n_1710)
);

OA21x2_ASAP7_75t_L g1711 ( 
.A1(n_1497),
.A2(n_1483),
.B(n_1520),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1524),
.B(n_1342),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1466),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1565),
.Y(n_1715)
);

O2A1O1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1557),
.A2(n_1565),
.B(n_1595),
.C(n_1592),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1595),
.C(n_1565),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1565),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1719)
);

AND2x2_ASAP7_75t_SL g1720 ( 
.A(n_1467),
.B(n_1087),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1617),
.A2(n_1455),
.B1(n_1442),
.B2(n_1566),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1497),
.A2(n_1483),
.B(n_1520),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1565),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1724)
);

OA22x2_ASAP7_75t_L g1725 ( 
.A1(n_1521),
.A2(n_1487),
.B1(n_1565),
.B2(n_1557),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1565),
.Y(n_1726)
);

CKINVDCx16_ASAP7_75t_R g1727 ( 
.A(n_1489),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1539),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1557),
.B(n_1455),
.Y(n_1731)
);

NOR2xp67_ASAP7_75t_R g1732 ( 
.A(n_1489),
.B(n_777),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1489),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1557),
.A2(n_1592),
.B(n_1565),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1518),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1686),
.B(n_1689),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1655),
.B(n_1632),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1707),
.Y(n_1739)
);

BUFx4f_ASAP7_75t_SL g1740 ( 
.A(n_1642),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1685),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1682),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1683),
.B(n_1699),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1624),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1688),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1685),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1651),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1635),
.B(n_1719),
.Y(n_1749)
);

AO21x2_ASAP7_75t_L g1750 ( 
.A1(n_1675),
.A2(n_1695),
.B(n_1702),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1665),
.B(n_1710),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1682),
.B(n_1626),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1680),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1720),
.Y(n_1754)
);

AO21x2_ASAP7_75t_L g1755 ( 
.A1(n_1715),
.A2(n_1726),
.B(n_1723),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1684),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1629),
.B(n_1711),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1700),
.B(n_1638),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1629),
.B(n_1711),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1707),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1707),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1707),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1687),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1713),
.B(n_1724),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1730),
.B(n_1734),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1707),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1718),
.B(n_1735),
.Y(n_1767)
);

INVx4_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

OA21x2_ASAP7_75t_L g1769 ( 
.A1(n_1634),
.A2(n_1669),
.B(n_1717),
.Y(n_1769)
);

OR2x6_ASAP7_75t_L g1770 ( 
.A(n_1716),
.B(n_1636),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1667),
.Y(n_1771)
);

AO21x2_ASAP7_75t_L g1772 ( 
.A1(n_1717),
.A2(n_1697),
.B(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1676),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1629),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1667),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1729),
.B(n_1711),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1722),
.B(n_1660),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1666),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1659),
.A2(n_1678),
.B(n_1650),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1639),
.B(n_1646),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1679),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1698),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1708),
.B(n_1709),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_SL g1784 ( 
.A(n_1664),
.B(n_1670),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1679),
.Y(n_1785)
);

CKINVDCx12_ASAP7_75t_R g1786 ( 
.A(n_1704),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1623),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1631),
.A2(n_1640),
.B1(n_1647),
.B2(n_1709),
.C(n_1708),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1623),
.Y(n_1789)
);

OA21x2_ASAP7_75t_L g1790 ( 
.A1(n_1690),
.A2(n_1731),
.B(n_1652),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1658),
.Y(n_1791)
);

OAI21x1_ASAP7_75t_L g1792 ( 
.A1(n_1701),
.A2(n_1673),
.B(n_1641),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1661),
.Y(n_1793)
);

AO21x2_ASAP7_75t_L g1794 ( 
.A1(n_1694),
.A2(n_1673),
.B(n_1731),
.Y(n_1794)
);

OR2x6_ASAP7_75t_L g1795 ( 
.A(n_1694),
.B(n_1657),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1725),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1788),
.A2(n_1725),
.B1(n_1644),
.B2(n_1721),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1756),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1788),
.B(n_1693),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1753),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1751),
.B(n_1777),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1625),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1776),
.B(n_1663),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1737),
.B(n_1630),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1739),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1757),
.B(n_1649),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1757),
.B(n_1648),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1759),
.B(n_1637),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1751),
.B(n_1643),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1742),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1776),
.B(n_1674),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1747),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1781),
.B(n_1654),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1780),
.B(n_1657),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1741),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1773),
.B(n_1627),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1778),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1767),
.A2(n_1706),
.B(n_1693),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1791),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1748),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1739),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1745),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1744),
.B(n_1696),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1783),
.B(n_1645),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1773),
.B(n_1705),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1785),
.B(n_1645),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1793),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1755),
.B(n_1736),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1744),
.B(n_1677),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1760),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1802),
.B(n_1761),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1802),
.B(n_1761),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1797),
.A2(n_1795),
.B1(n_1662),
.B2(n_1767),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1802),
.B(n_1762),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1801),
.B(n_1762),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1801),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_R g1838 ( 
.A(n_1827),
.B(n_1656),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1813),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1799),
.A2(n_1749),
.B1(n_1765),
.B2(n_1796),
.C(n_1789),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1800),
.Y(n_1841)
);

AOI21xp33_ASAP7_75t_L g1842 ( 
.A1(n_1799),
.A2(n_1755),
.B(n_1770),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1815),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1810),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1818),
.A2(n_1796),
.B(n_1787),
.C(n_1789),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1801),
.B(n_1743),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1818),
.A2(n_1668),
.B(n_1671),
.C(n_1692),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1797),
.A2(n_1795),
.B1(n_1767),
.B2(n_1790),
.Y(n_1848)
);

OAI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1824),
.A2(n_1767),
.B1(n_1795),
.B2(n_1770),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1817),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1801),
.B(n_1763),
.Y(n_1851)
);

OR2x6_ASAP7_75t_L g1852 ( 
.A(n_1813),
.B(n_1795),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1801),
.B(n_1766),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1766),
.Y(n_1854)
);

AO21x2_ASAP7_75t_L g1855 ( 
.A1(n_1829),
.A2(n_1774),
.B(n_1782),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_SL g1856 ( 
.A(n_1813),
.B(n_1765),
.C(n_1796),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1817),
.B(n_1764),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1813),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1822),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1810),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1803),
.B(n_1758),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1827),
.A2(n_1795),
.B(n_1770),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1828),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1827),
.A2(n_1795),
.B1(n_1767),
.B2(n_1790),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1826),
.A2(n_1770),
.B(n_1784),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1826),
.A2(n_1789),
.B1(n_1787),
.B2(n_1794),
.C(n_1772),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1812),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1815),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1812),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1820),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1814),
.B(n_1764),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1814),
.A2(n_1784),
.B1(n_1790),
.B2(n_1779),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1821),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1816),
.A2(n_1790),
.B1(n_1779),
.B2(n_1768),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1814),
.A2(n_1768),
.B1(n_1779),
.B2(n_1794),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1820),
.Y(n_1876)
);

BUFx10_ASAP7_75t_L g1877 ( 
.A(n_1828),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1816),
.A2(n_1779),
.B1(n_1794),
.B2(n_1768),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1806),
.B(n_1752),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_SL g1880 ( 
.A(n_1798),
.B(n_1727),
.C(n_1733),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1806),
.B(n_1752),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1809),
.A2(n_1779),
.B1(n_1768),
.B2(n_1794),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1807),
.B(n_1738),
.Y(n_1883)
);

OR2x6_ASAP7_75t_L g1884 ( 
.A(n_1828),
.B(n_1754),
.Y(n_1884)
);

NOR3xp33_ASAP7_75t_SL g1885 ( 
.A(n_1838),
.B(n_1703),
.C(n_1798),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1837),
.B(n_1807),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1843),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1841),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1872),
.B(n_1809),
.Y(n_1889)
);

INVx4_ASAP7_75t_L g1890 ( 
.A(n_1858),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1870),
.Y(n_1891)
);

AO21x2_ASAP7_75t_L g1892 ( 
.A1(n_1842),
.A2(n_1750),
.B(n_1746),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1837),
.B(n_1821),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1870),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1865),
.A2(n_1775),
.B(n_1771),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1878),
.A2(n_1772),
.B(n_1803),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1852),
.B(n_1754),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1836),
.B(n_1808),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1836),
.B(n_1808),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1876),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1878),
.B(n_1866),
.C(n_1875),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1861),
.B(n_1811),
.Y(n_1904)
);

INVx4_ASAP7_75t_SL g1905 ( 
.A(n_1852),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1876),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1848),
.A2(n_1874),
.B(n_1849),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1868),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1871),
.B(n_1653),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1840),
.B(n_1809),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1844),
.Y(n_1911)
);

INVx6_ASAP7_75t_L g1912 ( 
.A(n_1877),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1850),
.B(n_1653),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1862),
.B(n_1809),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1861),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1877),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1857),
.B(n_1808),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1859),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1844),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1834),
.A2(n_1792),
.B(n_1769),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_SL g1921 ( 
.A(n_1852),
.B(n_1819),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1884),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1860),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1882),
.B(n_1809),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1854),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1839),
.Y(n_1926)
);

BUFx3_ASAP7_75t_L g1927 ( 
.A(n_1877),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1863),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1904),
.B(n_1860),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1891),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1905),
.B(n_1853),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1903),
.B(n_1864),
.C(n_1856),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1918),
.B(n_1804),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1891),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1905),
.B(n_1853),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1903),
.B(n_1852),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1904),
.B(n_1867),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1915),
.B(n_1804),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1905),
.B(n_1897),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1905),
.B(n_1879),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1926),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1887),
.B(n_1867),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1905),
.B(n_1879),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1897),
.B(n_1881),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1897),
.B(n_1881),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1917),
.B(n_1830),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1897),
.B(n_1873),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1901),
.B(n_1873),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1925),
.B(n_1804),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1888),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1894),
.Y(n_1951)
);

AOI322xp5_ASAP7_75t_L g1952 ( 
.A1(n_1907),
.A2(n_1845),
.A3(n_1880),
.B1(n_1833),
.B2(n_1832),
.C1(n_1835),
.C2(n_1854),
.Y(n_1952)
);

NAND2x1_ASAP7_75t_SL g1953 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1908),
.B(n_1869),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1894),
.Y(n_1955)
);

OR2x6_ASAP7_75t_L g1956 ( 
.A(n_1920),
.B(n_1754),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1902),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1902),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1888),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1888),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1911),
.B(n_1869),
.Y(n_1961)
);

AND2x2_ASAP7_75t_SL g1962 ( 
.A(n_1890),
.B(n_1769),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1911),
.B(n_1855),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1926),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1885),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1926),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1912),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1906),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1901),
.B(n_1832),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1901),
.B(n_1833),
.Y(n_1970)
);

OAI222xp33_ASAP7_75t_L g1971 ( 
.A1(n_1889),
.A2(n_1884),
.B1(n_1823),
.B2(n_1831),
.C1(n_1805),
.C2(n_1811),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1923),
.B(n_1855),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1896),
.B(n_1847),
.C(n_1769),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1907),
.A2(n_1772),
.B1(n_1754),
.B2(n_1769),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1922),
.B(n_1835),
.Y(n_1975)
);

NAND4xp25_ASAP7_75t_L g1976 ( 
.A(n_1896),
.B(n_1778),
.C(n_1823),
.D(n_1628),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1923),
.B(n_1855),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1924),
.A2(n_1884),
.B1(n_1763),
.B2(n_1672),
.C(n_1811),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1922),
.B(n_1851),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1921),
.B(n_1846),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1906),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1921),
.B(n_1846),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1893),
.B(n_1883),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1940),
.B(n_1893),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1932),
.B(n_1910),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1980),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_SL g1987 ( 
.A(n_1965),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1952),
.B(n_1899),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1940),
.B(n_1890),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1965),
.A2(n_1914),
.B(n_1920),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1933),
.B(n_1899),
.Y(n_1991)
);

O2A1O1Ixp33_ASAP7_75t_L g1992 ( 
.A1(n_1936),
.A2(n_1913),
.B(n_1909),
.C(n_1928),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1936),
.A2(n_1681),
.B(n_1732),
.Y(n_1993)
);

AOI21xp33_ASAP7_75t_SL g1994 ( 
.A1(n_1936),
.A2(n_1973),
.B(n_1978),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1938),
.B(n_1900),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1943),
.B(n_1890),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1963),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1941),
.B(n_1900),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1930),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1964),
.B(n_1966),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1939),
.B(n_1916),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1929),
.B(n_1919),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1975),
.B(n_1886),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1934),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1951),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1955),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1967),
.B(n_1681),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1957),
.Y(n_2009)
);

NOR2x1_ASAP7_75t_L g2010 ( 
.A(n_1936),
.B(n_1927),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1949),
.B(n_1946),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1958),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1953),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1974),
.A2(n_1898),
.B1(n_1890),
.B2(n_1912),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1968),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1976),
.B(n_1830),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1939),
.B(n_1728),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1981),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1980),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1972),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1961),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1961),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1975),
.B(n_1886),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1972),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2003),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2019),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2000),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1986),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_2019),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1987),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_2010),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2013),
.B(n_1980),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2013),
.B(n_1986),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2003),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_2001),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2021),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2022),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1999),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1986),
.B(n_1982),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1989),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_2004),
.B(n_1929),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1984),
.B(n_1982),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1984),
.B(n_1982),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2005),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_2023),
.B(n_1937),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1989),
.B(n_1931),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1997),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2006),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2007),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1996),
.B(n_1931),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1985),
.B(n_1942),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1997),
.Y(n_2052)
);

INVxp33_ASAP7_75t_L g2053 ( 
.A(n_2017),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1996),
.B(n_1935),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2046),
.B(n_2017),
.Y(n_2055)
);

OAI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_2030),
.A2(n_1990),
.B1(n_1994),
.B2(n_1988),
.C(n_1993),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2031),
.A2(n_2035),
.B1(n_1956),
.B2(n_2014),
.Y(n_2057)
);

OAI31xp33_ASAP7_75t_L g2058 ( 
.A1(n_2031),
.A2(n_1992),
.A3(n_1971),
.B(n_2001),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_2040),
.B(n_2008),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2052),
.Y(n_2060)
);

OAI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2035),
.A2(n_1956),
.B1(n_2016),
.B2(n_1898),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2052),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_2030),
.B(n_2008),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2026),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2040),
.A2(n_1956),
.B1(n_1998),
.B2(n_1898),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2027),
.B(n_2009),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2026),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2027),
.A2(n_1956),
.B1(n_1962),
.B2(n_2012),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2042),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2025),
.B(n_2015),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_L g2071 ( 
.A(n_2025),
.B(n_2018),
.C(n_1962),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_2053),
.B(n_1740),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2033),
.B(n_2029),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_R g2074 ( 
.A(n_2033),
.B(n_1943),
.Y(n_2074)
);

AND2x2_ASAP7_75t_SL g2075 ( 
.A(n_2051),
.B(n_1935),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2029),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2034),
.B(n_1983),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2051),
.A2(n_1892),
.B1(n_1947),
.B2(n_1948),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2055),
.B(n_2059),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_2063),
.B(n_2034),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2073),
.B(n_2033),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2073),
.B(n_2046),
.Y(n_2082)
);

NAND2xp33_ASAP7_75t_L g2083 ( 
.A(n_2069),
.B(n_2046),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2060),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2075),
.B(n_2050),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2064),
.B(n_2050),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2062),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2067),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2076),
.B(n_2077),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2072),
.B(n_2050),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_2056),
.B(n_2036),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2070),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2057),
.B(n_2054),
.Y(n_2093)
);

AOI221xp5_ASAP7_75t_L g2094 ( 
.A1(n_2091),
.A2(n_2058),
.B1(n_2071),
.B2(n_2066),
.C(n_2061),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2079),
.B(n_2054),
.Y(n_2095)
);

AOI221xp5_ASAP7_75t_L g2096 ( 
.A1(n_2091),
.A2(n_2036),
.B1(n_2037),
.B2(n_2068),
.C(n_2065),
.Y(n_2096)
);

OAI211xp5_ASAP7_75t_SL g2097 ( 
.A1(n_2080),
.A2(n_2068),
.B(n_2078),
.C(n_2037),
.Y(n_2097)
);

AOI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2080),
.A2(n_2032),
.B(n_2054),
.C(n_2044),
.Y(n_2098)
);

NAND3xp33_ASAP7_75t_SL g2099 ( 
.A(n_2085),
.B(n_2032),
.C(n_2078),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2093),
.A2(n_2074),
.B1(n_2032),
.B2(n_2043),
.Y(n_2100)
);

NAND4xp25_ASAP7_75t_L g2101 ( 
.A(n_2090),
.B(n_2082),
.C(n_2086),
.D(n_2089),
.Y(n_2101)
);

OAI21xp33_ASAP7_75t_SL g2102 ( 
.A1(n_2081),
.A2(n_2043),
.B(n_2042),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2092),
.B(n_2041),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_2083),
.A2(n_2028),
.B(n_2039),
.Y(n_2104)
);

OAI211xp5_ASAP7_75t_SL g2105 ( 
.A1(n_2088),
.A2(n_2038),
.B(n_2048),
.C(n_2044),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2095),
.Y(n_2106)
);

NOR4xp25_ASAP7_75t_L g2107 ( 
.A(n_2097),
.B(n_2084),
.C(n_2087),
.D(n_2028),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2104),
.Y(n_2108)
);

AOI222xp33_ASAP7_75t_L g2109 ( 
.A1(n_2099),
.A2(n_2087),
.B1(n_2049),
.B2(n_2048),
.C1(n_2038),
.C2(n_2047),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2094),
.A2(n_2043),
.B1(n_2042),
.B2(n_2039),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_2096),
.A2(n_2028),
.B(n_2049),
.Y(n_2111)
);

AOI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_2102),
.A2(n_2047),
.B1(n_2039),
.B2(n_2041),
.C(n_2045),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2106),
.B(n_2101),
.Y(n_2113)
);

OAI21xp33_ASAP7_75t_L g2114 ( 
.A1(n_2110),
.A2(n_2100),
.B(n_2103),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2107),
.B(n_2098),
.Y(n_2115)
);

CKINVDCx16_ASAP7_75t_R g2116 ( 
.A(n_2108),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2112),
.B(n_2045),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2109),
.Y(n_2118)
);

OAI21xp33_ASAP7_75t_L g2119 ( 
.A1(n_2111),
.A2(n_2105),
.B(n_2047),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2113),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2118),
.A2(n_2020),
.B1(n_2002),
.B2(n_2024),
.Y(n_2121)
);

AOI21xp5_ASAP7_75t_L g2122 ( 
.A1(n_2115),
.A2(n_2020),
.B(n_2002),
.Y(n_2122)
);

INVx2_ASAP7_75t_SL g2123 ( 
.A(n_2116),
.Y(n_2123)
);

OAI211xp5_ASAP7_75t_L g2124 ( 
.A1(n_2119),
.A2(n_1712),
.B(n_2024),
.C(n_1947),
.Y(n_2124)
);

OAI21xp33_ASAP7_75t_L g2125 ( 
.A1(n_2114),
.A2(n_1948),
.B(n_2011),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_2123),
.B(n_2117),
.Y(n_2126)
);

NAND4xp25_ASAP7_75t_L g2127 ( 
.A(n_2125),
.B(n_1622),
.C(n_1633),
.D(n_1991),
.Y(n_2127)
);

NOR3x1_ASAP7_75t_L g2128 ( 
.A(n_2124),
.B(n_1895),
.C(n_1977),
.Y(n_2128)
);

NOR3xp33_ASAP7_75t_L g2129 ( 
.A(n_2126),
.B(n_2120),
.C(n_2122),
.Y(n_2129)
);

OAI31xp33_ASAP7_75t_L g2130 ( 
.A1(n_2129),
.A2(n_2121),
.A3(n_2127),
.B(n_2128),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2130),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_2130),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_SL g2133 ( 
.A1(n_2131),
.A2(n_1786),
.B1(n_1912),
.B2(n_1633),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_1979),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2134),
.A2(n_2132),
.B(n_1995),
.Y(n_2135)
);

OAI22x1_ASAP7_75t_L g2136 ( 
.A1(n_2133),
.A2(n_1959),
.B1(n_1960),
.B2(n_1950),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_SL g2137 ( 
.A1(n_2135),
.A2(n_1912),
.B1(n_1916),
.B2(n_1927),
.Y(n_2137)
);

OAI21xp33_ASAP7_75t_L g2138 ( 
.A1(n_2137),
.A2(n_2136),
.B(n_1979),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2138),
.A2(n_1954),
.B(n_1942),
.Y(n_2139)
);

AOI322xp5_ASAP7_75t_L g2140 ( 
.A1(n_2139),
.A2(n_1950),
.A3(n_1959),
.B1(n_1960),
.B2(n_1927),
.C1(n_1970),
.C2(n_1969),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_SL g2141 ( 
.A1(n_2140),
.A2(n_1944),
.B(n_1945),
.C(n_1970),
.Y(n_2141)
);

AOI211xp5_ASAP7_75t_L g2142 ( 
.A1(n_2141),
.A2(n_1977),
.B(n_1691),
.C(n_1954),
.Y(n_2142)
);


endmodule