module real_jpeg_5389_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_89),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_107),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_107),
.B1(n_183),
.B2(n_275),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_1),
.A2(n_107),
.B1(n_297),
.B2(n_300),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_30),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_30),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_93),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_3),
.A2(n_260),
.B(n_262),
.C(n_266),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_3),
.B(n_287),
.C(n_289),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_3),
.B(n_129),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_3),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_3),
.B(n_49),
.Y(n_326)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_5),
.Y(n_314)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_5),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_43),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_43),
.B1(n_123),
.B2(n_127),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_43),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_9),
.Y(n_210)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_10),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_11),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_11),
.A2(n_66),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_11),
.A2(n_66),
.B1(n_267),
.B2(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_363),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_227),
.B(n_361),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_195),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_15),
.B(n_195),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_169),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_159),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_17),
.B(n_159),
.C(n_169),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_84),
.B2(n_85),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_18),
.B(n_86),
.C(n_120),
.Y(n_389)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_47),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_20),
.B(n_47),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_21),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_24),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_26),
.A2(n_35),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_26),
.B(n_35),
.Y(n_238)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_30),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_30),
.B(n_91),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_30),
.A2(n_263),
.B(n_265),
.Y(n_262)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_33),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_34),
.A2(n_172),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_35),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_38),
.B(n_40),
.Y(n_177)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_42),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_59),
.B(n_69),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_48),
.A2(n_166),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_48),
.B(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_70),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_49),
.B(n_274),
.Y(n_291)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_54),
.Y(n_300)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_57),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_57),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_59),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_62),
.Y(n_265)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_65),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_69),
.B(n_291),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_69),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_72),
.Y(n_285)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_76),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_76),
.B(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_131),
.B1(n_134),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_120),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_105),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_88),
.B(n_109),
.Y(n_243)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_88),
.Y(n_378)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_93),
.B(n_106),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_93),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_93),
.Y(n_377)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_103),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_109),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_139),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_121),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_122),
.Y(n_248)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_128),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_140),
.B(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_129),
.B(n_221),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_129),
.A2(n_247),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_130),
.B(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_133),
.Y(n_264)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_138),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_139),
.B(n_249),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_154),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_140),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_141),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_148),
.Y(n_268)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_154),
.Y(n_219)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_164),
.B1(n_165),
.B2(n_168),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_160),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_160),
.A2(n_168),
.B1(n_259),
.B2(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_160),
.B(n_165),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_160),
.A2(n_168),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_167),
.B(n_273),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_185),
.C(n_187),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_171),
.B(n_178),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_177),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_177),
.B(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_179),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_194),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_226),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_196),
.B(n_226),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_199),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_216),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_200),
.B(n_216),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_202),
.B(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_205),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_208),
.A3(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_347),
.B(n_358),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_278),
.B(n_346),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_254),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_230),
.B(n_254),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_240),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.C(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_269),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_255),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_258),
.A2(n_269),
.B1(n_270),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_258),
.Y(n_343)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_272),
.B(n_387),
.Y(n_386)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_340),
.B(n_345),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_330),
.B(n_339),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_306),
.B(n_329),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_292),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_292),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_284),
.B1(n_290),
.B2(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_304),
.C(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_315),
.B(n_328),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_310),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_324),
.B(n_327),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_333),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_344),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_350),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_356),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.CI(n_353),
.CON(n_350),
.SN(n_350)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_359),
.B(n_360),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_390),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_366),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_389),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_379),
.B2(n_380),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_372),
.B2(n_373),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B(n_378),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_386),
.B(n_388),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_381),
.B(n_386),
.Y(n_388)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);


endmodule