module fake_ariane_830_n_1557 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1557);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1557;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_1548;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_256),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_7),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_41),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_129),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_309),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_150),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_92),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_242),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_217),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_12),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_269),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_236),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_241),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_86),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_190),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_141),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_215),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_33),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_221),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_212),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_64),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_86),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_31),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_88),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_169),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_124),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_307),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_204),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_189),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_156),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_99),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_178),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_160),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_17),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_229),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_254),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_30),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_272),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_134),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_88),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_101),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_110),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_159),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_38),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_286),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_90),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_228),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_119),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_54),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_276),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_264),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_122),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_2),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_206),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_145),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_223),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_131),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_188),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_191),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_10),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_61),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_201),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_275),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_29),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_115),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_168),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_142),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_182),
.Y(n_395)
);

BUFx8_ASAP7_75t_SL g396 ( 
.A(n_128),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_257),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_16),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_38),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_167),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_239),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_21),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_175),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_3),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_93),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_216),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_85),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_253),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_126),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_35),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_219),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_163),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_282),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_108),
.Y(n_415)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_125),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_14),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_46),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_66),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_42),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_117),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_36),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_30),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_24),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_84),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_75),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_106),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_82),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_187),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_138),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_196),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_179),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_40),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_313),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_273),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_195),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_183),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_57),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_137),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_87),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_143),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_5),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_277),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_9),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_185),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_296),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_301),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_148),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_291),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_246),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_139),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_127),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_180),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_32),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_112),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_184),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_44),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_83),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_114),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_176),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_200),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_79),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_230),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_102),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_155),
.Y(n_467)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_44),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_79),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_306),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_74),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_294),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_237),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_57),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_194),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_283),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_73),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_220),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_170),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_54),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_15),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_181),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_166),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_238),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_13),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_69),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_70),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_36),
.Y(n_488)
);

INVx4_ASAP7_75t_R g489 ( 
.A(n_48),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_24),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_3),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_8),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_66),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_116),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_77),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_295),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_49),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_22),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_4),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_203),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_8),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_284),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_235),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_162),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_49),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_136),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_69),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_21),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_245),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_48),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_278),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_55),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_251),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_18),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_247),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_97),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_32),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_165),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_287),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_281),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_255),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_18),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_58),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_1),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_80),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_31),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_53),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_250),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_302),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_35),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_71),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_186),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_20),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_298),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_56),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_14),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_96),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_53),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_10),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_192),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_104),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_316),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_177),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_113),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_174),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_149),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_198),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_12),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_118),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_0),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_334),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_334),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_0),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_468),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_366),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_468),
.B(n_1),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_449),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_449),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_387),
.B(n_4),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_323),
.B(n_5),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_468),
.B(n_6),
.Y(n_561)
);

BUFx8_ASAP7_75t_L g562 ( 
.A(n_466),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_387),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_343),
.B(n_6),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_468),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_343),
.B(n_7),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_344),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_468),
.B(n_9),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_442),
.B(n_11),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_399),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_429),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_344),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_344),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_321),
.B(n_11),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_344),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_460),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_342),
.Y(n_579)
);

BUFx12f_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_436),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_325),
.B(n_13),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_369),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_396),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_15),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_353),
.B(n_16),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_369),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_369),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_339),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_354),
.B(n_19),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_333),
.B(n_359),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_357),
.B(n_19),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_361),
.B(n_20),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_369),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_363),
.B(n_22),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_333),
.B(n_23),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_367),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_368),
.B(n_23),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

CKINVDCx6p67_ASAP7_75t_R g604 ( 
.A(n_364),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_372),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_367),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_542),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_385),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_396),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_379),
.B(n_25),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_389),
.B(n_390),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_392),
.B(n_25),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_382),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_359),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_530),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_380),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_382),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_393),
.B(n_26),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_385),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_450),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_400),
.B(n_26),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_391),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_403),
.B(n_27),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_406),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_458),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_340),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_459),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_413),
.B(n_27),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_319),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_326),
.B(n_28),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_405),
.Y(n_631)
);

XNOR2x1_ASAP7_75t_L g632 ( 
.A(n_434),
.B(n_28),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_430),
.B(n_29),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_459),
.B(n_33),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_530),
.B(n_34),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_493),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_34),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_431),
.B(n_37),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_493),
.B(n_37),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_408),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_342),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_507),
.B(n_39),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_420),
.B(n_39),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_450),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_432),
.B(n_40),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_435),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_424),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_494),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_494),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_438),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_549),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_326),
.B(n_41),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_428),
.B(n_42),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_448),
.B(n_43),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_457),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_441),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_444),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_508),
.B(n_43),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_320),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_517),
.B(n_45),
.Y(n_661)
);

BUFx12f_ASAP7_75t_L g662 ( 
.A(n_329),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_464),
.B(n_45),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_462),
.B(n_46),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_495),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_467),
.B(n_47),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_47),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_335),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_548),
.B(n_50),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_371),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_345),
.Y(n_672)
);

BUFx12f_ASAP7_75t_L g673 ( 
.A(n_356),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_499),
.Y(n_674)
);

CKINVDCx11_ASAP7_75t_R g675 ( 
.A(n_411),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_473),
.B(n_50),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_510),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_512),
.B(n_51),
.Y(n_678)
);

BUFx12f_ASAP7_75t_L g679 ( 
.A(n_375),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_475),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_478),
.B(n_51),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_522),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_317),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_524),
.B(n_52),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_533),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_479),
.B(n_52),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_482),
.B(n_506),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_513),
.B(n_55),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_388),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_515),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_518),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_529),
.B(n_56),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_398),
.Y(n_695)
);

BUFx8_ASAP7_75t_SL g696 ( 
.A(n_411),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_547),
.B(n_58),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_338),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_417),
.B(n_59),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_418),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_384),
.B(n_386),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_419),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_330),
.B(n_59),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_318),
.B(n_60),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_332),
.B(n_348),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_338),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_422),
.B(n_60),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_338),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_519),
.B(n_61),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_705),
.A2(n_386),
.B1(n_427),
.B2(n_384),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_705),
.A2(n_463),
.B1(n_470),
.B2(n_427),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_630),
.A2(n_653),
.B1(n_709),
.B2(n_703),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_624),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_578),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_624),
.B(n_540),
.Y(n_715)
);

AOI22x1_ASAP7_75t_SL g716 ( 
.A1(n_586),
.A2(n_523),
.B1(n_531),
.B2(n_480),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_572),
.B(n_322),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_568),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_615),
.B(n_416),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_630),
.A2(n_470),
.B1(n_476),
.B2(n_463),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_624),
.B(n_324),
.Y(n_721)
);

NAND3x1_ASAP7_75t_L g722 ( 
.A(n_623),
.B(n_523),
.C(n_480),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_568),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_653),
.A2(n_503),
.B1(n_546),
.B2(n_476),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_560),
.A2(n_570),
.B1(n_701),
.B2(n_567),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_574),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_625),
.B(n_423),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_625),
.B(n_582),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_574),
.Y(n_732)
);

NAND3x1_ASAP7_75t_L g733 ( 
.A(n_635),
.B(n_531),
.C(n_503),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_570),
.A2(n_426),
.B1(n_446),
.B2(n_425),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_632),
.A2(n_489),
.B1(n_546),
.B2(n_469),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_703),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_709),
.A2(n_474),
.B1(n_477),
.B2(n_456),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_592),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_SL g739 ( 
.A1(n_701),
.A2(n_485),
.B1(n_486),
.B2(n_481),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_604),
.A2(n_488),
.B1(n_490),
.B2(n_487),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_683),
.B(n_327),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_581),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_625),
.B(n_491),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_683),
.B(n_328),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_564),
.A2(n_498),
.B1(n_501),
.B2(n_492),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_571),
.A2(n_514),
.B1(n_525),
.B2(n_505),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_572),
.B(n_331),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_572),
.B(n_573),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_581),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_572),
.B(n_336),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_637),
.A2(n_527),
.B1(n_535),
.B2(n_526),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_588),
.B(n_538),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_SL g753 ( 
.A1(n_555),
.A2(n_539),
.B1(n_341),
.B2(n_346),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_573),
.B(n_337),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_575),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_581),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_564),
.A2(n_347),
.B1(n_350),
.B2(n_349),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_567),
.A2(n_352),
.B1(n_355),
.B2(n_351),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_358),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_599),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_605),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_602),
.B(n_360),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_659),
.A2(n_362),
.B1(n_370),
.B2(n_365),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_609),
.A2(n_573),
.B1(n_603),
.B2(n_602),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_573),
.B(n_373),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_566),
.A2(n_376),
.B1(n_377),
.B2(n_374),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_616),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_611),
.A2(n_381),
.B1(n_383),
.B2(n_378),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_579),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_603),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_599),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_575),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_603),
.B(n_394),
.Y(n_773)
);

AND2x2_ASAP7_75t_SL g774 ( 
.A(n_634),
.B(n_395),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_661),
.A2(n_397),
.B1(n_402),
.B2(n_401),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_667),
.A2(n_404),
.B1(n_409),
.B2(n_407),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_643),
.A2(n_68),
.B1(n_65),
.B2(n_67),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_668),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_580),
.B(n_67),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_609),
.A2(n_412),
.B1(n_414),
.B2(n_410),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_665),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_575),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_551),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_669),
.A2(n_415),
.B1(n_433),
.B2(n_421),
.Y(n_784)
);

AND2x2_ASAP7_75t_SL g785 ( 
.A(n_634),
.B(n_437),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_643),
.A2(n_587),
.B1(n_559),
.B2(n_594),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_629),
.A2(n_689),
.B1(n_672),
.B2(n_707),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_677),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_577),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_L g790 ( 
.A1(n_576),
.A2(n_544),
.B1(n_543),
.B2(n_541),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_642),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_682),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_686),
.A2(n_537),
.B1(n_532),
.B2(n_528),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_702),
.B(n_440),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_686),
.A2(n_521),
.B1(n_520),
.B2(n_516),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_577),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_577),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_695),
.B(n_443),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_600),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_613),
.B(n_445),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_600),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_SL g802 ( 
.A1(n_699),
.A2(n_511),
.B1(n_509),
.B2(n_504),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_660),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_576),
.A2(n_502),
.B1(n_500),
.B2(n_496),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_600),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_585),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_695),
.B(n_447),
.Y(n_807)
);

AO22x2_ASAP7_75t_L g808 ( 
.A1(n_559),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_SL g809 ( 
.A(n_688),
.B(n_451),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_606),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_688),
.A2(n_484),
.B1(n_483),
.B2(n_472),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_647),
.B(n_452),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_SL g813 ( 
.A1(n_699),
.A2(n_465),
.B1(n_455),
.B2(n_454),
.Y(n_813)
);

NAND3x1_ASAP7_75t_L g814 ( 
.A(n_584),
.B(n_72),
.C(n_73),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_585),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_738),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_R g817 ( 
.A(n_752),
.B(n_594),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_761),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_710),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_799),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_720),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_781),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_788),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_725),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_711),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_792),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_714),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_713),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_799),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_794),
.B(n_671),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_712),
.B(n_587),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_801),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_736),
.B(n_693),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_801),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_736),
.B(n_662),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_671),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_805),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_810),
.Y(n_839)
);

XOR2xp5_ASAP7_75t_L g840 ( 
.A(n_791),
.B(n_696),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_798),
.B(n_671),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_726),
.Y(n_842)
);

XOR2xp5_ASAP7_75t_L g843 ( 
.A(n_769),
.B(n_675),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_726),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_783),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_783),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_718),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_815),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_724),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_730),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_778),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_732),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_729),
.A2(n_553),
.B(n_550),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_755),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_772),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_782),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_789),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_796),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_797),
.Y(n_860)
);

XOR2xp5_ASAP7_75t_L g861 ( 
.A(n_735),
.B(n_704),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_728),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_786),
.B(n_673),
.Y(n_863)
);

AND2x6_ASAP7_75t_L g864 ( 
.A(n_731),
.B(n_640),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_757),
.B(n_639),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_812),
.Y(n_867)
);

XNOR2xp5_ASAP7_75t_L g868 ( 
.A(n_733),
.B(n_562),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_728),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_728),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_749),
.B(n_644),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_774),
.B(n_679),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_713),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_806),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_803),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_750),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_785),
.B(n_640),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_743),
.A2(n_553),
.B(n_550),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_787),
.B(n_700),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_806),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_741),
.A2(n_561),
.B(n_556),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_759),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_762),
.Y(n_884)
);

XOR2xp5_ASAP7_75t_L g885 ( 
.A(n_735),
.B(n_704),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_739),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_716),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_773),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_744),
.B(n_613),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_800),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_754),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_719),
.B(n_627),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_754),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_719),
.B(n_627),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_765),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_765),
.B(n_613),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_742),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_717),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_747),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_756),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_770),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_563),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_793),
.B(n_617),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_745),
.B(n_583),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_727),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_760),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_760),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_751),
.B(n_614),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_715),
.B(n_551),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_614),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_811),
.B(n_644),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_771),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_716),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_795),
.B(n_639),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_814),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_820),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_862),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_876),
.B(n_763),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_876),
.B(n_775),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_816),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_865),
.B(n_771),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_832),
.B(n_654),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_864),
.B(n_776),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_852),
.B(n_784),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_864),
.B(n_790),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_829),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_865),
.B(n_777),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_818),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_890),
.B(n_878),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_862),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_822),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_823),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_878),
.B(n_777),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_824),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_819),
.B(n_758),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_864),
.B(n_804),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_808),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_819),
.B(n_768),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_827),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_864),
.B(n_654),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_864),
.B(n_663),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_841),
.B(n_663),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_832),
.B(n_684),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_820),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_830),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_882),
.A2(n_879),
.B(n_854),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_834),
.B(n_808),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_841),
.B(n_684),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_903),
.B(n_690),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_906),
.B(n_694),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_829),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_833),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_912),
.B(n_584),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_817),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_873),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_835),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_862),
.Y(n_958)
);

AND2x2_ASAP7_75t_SL g959 ( 
.A(n_912),
.B(n_589),
.Y(n_959)
);

BUFx4_ASAP7_75t_SL g960 ( 
.A(n_875),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_873),
.B(n_611),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_817),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_862),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_907),
.B(n_678),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_871),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_860),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_908),
.B(n_641),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_828),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_899),
.B(n_809),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_913),
.B(n_641),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_892),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_860),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_909),
.B(n_657),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_838),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_839),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_847),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_842),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_831),
.B(n_721),
.Y(n_978)
);

CKINVDCx12_ASAP7_75t_R g979 ( 
.A(n_863),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_836),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_832),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_831),
.B(n_900),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_883),
.B(n_589),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_894),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_884),
.B(n_593),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_911),
.B(n_657),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_848),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_867),
.B(n_685),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_916),
.B(n_593),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_897),
.A2(n_561),
.B(n_556),
.Y(n_990)
);

AND2x2_ASAP7_75t_SL g991 ( 
.A(n_916),
.B(n_866),
.Y(n_991)
);

AND2x2_ASAP7_75t_SL g992 ( 
.A(n_866),
.B(n_596),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_872),
.B(n_685),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_832),
.B(n_779),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_888),
.B(n_622),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_844),
.Y(n_996)
);

AND2x6_ASAP7_75t_L g997 ( 
.A(n_897),
.B(n_891),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_849),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_893),
.B(n_802),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_871),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_895),
.B(n_722),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_845),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_846),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_846),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_880),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_850),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_869),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_832),
.B(n_631),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_870),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_851),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_853),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_855),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_837),
.B(n_596),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_915),
.B(n_648),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_915),
.B(n_658),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_856),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_910),
.B(n_670),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_898),
.B(n_779),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_837),
.B(n_601),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_910),
.B(n_896),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_904),
.B(n_889),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_857),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_601),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_927),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_971),
.B(n_861),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_947),
.B(n_858),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_994),
.B(n_902),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_992),
.B(n_859),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_955),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_984),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_994),
.B(n_886),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_981),
.B(n_874),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_919),
.B(n_885),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_945),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_920),
.B(n_821),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_981),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_1018),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_925),
.B(n_821),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_994),
.B(n_886),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_981),
.B(n_825),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_918),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_950),
.B(n_825),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_927),
.B(n_826),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_952),
.B(n_956),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_952),
.B(n_826),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_1000),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_950),
.B(n_868),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_993),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_992),
.B(n_554),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_938),
.B(n_636),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_956),
.B(n_923),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_945),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_918),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_917),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_917),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_966),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_924),
.B(n_764),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1005),
.B(n_840),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_918),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1013),
.B(n_565),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_965),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_923),
.B(n_766),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_918),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1019),
.B(n_687),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_966),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_918),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_674),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_962),
.B(n_734),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_993),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_921),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_929),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_931),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_931),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_991),
.B(n_687),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_991),
.B(n_698),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_944),
.B(n_753),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_980),
.B(n_746),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_931),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_944),
.B(n_813),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_931),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_931),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_932),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_1008),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_938),
.B(n_843),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_972),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_972),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_944),
.B(n_552),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_958),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1008),
.B(n_877),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_706),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_954),
.B(n_610),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_990),
.A2(n_1021),
.B(n_982),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_958),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_922),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_928),
.B(n_881),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1014),
.B(n_636),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_935),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_934),
.B(n_552),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1015),
.B(n_552),
.Y(n_1105)
);

NOR2xp67_ASAP7_75t_SL g1106 ( 
.A(n_941),
.B(n_610),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_958),
.Y(n_1107)
);

BUFx5_ASAP7_75t_L g1108 ( 
.A(n_997),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_946),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_928),
.B(n_887),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1098),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1075),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_1043),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_1025),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1032),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_1084),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1039),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_1102),
.B(n_934),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1098),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1059),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1068),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1037),
.B(n_922),
.Y(n_1122)
);

BUFx4_ASAP7_75t_SL g1123 ( 
.A(n_1079),
.Y(n_1123)
);

BUFx4f_ASAP7_75t_SL g1124 ( 
.A(n_1024),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_1045),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1035),
.A2(n_954),
.B1(n_959),
.B2(n_936),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1073),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1045),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1104),
.B(n_999),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1044),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_1046),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1047),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1040),
.B(n_959),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1074),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1084),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1047),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1089),
.Y(n_1137)
);

CKINVDCx14_ASAP7_75t_R g1138 ( 
.A(n_1061),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1037),
.B(n_939),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1024),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1048),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1046),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1040),
.B(n_948),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1085),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_1033),
.Y(n_1145)
);

BUFx5_ASAP7_75t_L g1146 ( 
.A(n_1075),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1087),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1067),
.B(n_930),
.Y(n_1148)
);

CKINVDCx8_ASAP7_75t_R g1149 ( 
.A(n_1033),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1101),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1103),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_1084),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_1076),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1053),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1081),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1084),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1043),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1102),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1053),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1091),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1076),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1102),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1091),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1064),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1090),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1031),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1031),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1091),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_1029),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1038),
.B(n_958),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1056),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1038),
.B(n_958),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1109),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1057),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1081),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1043),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1070),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1041),
.Y(n_1178)
);

BUFx8_ASAP7_75t_SL g1179 ( 
.A(n_1082),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1055),
.Y(n_1180)
);

INVx6_ASAP7_75t_SL g1181 ( 
.A(n_1079),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1088),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1067),
.B(n_989),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_1140),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1124),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1120),
.Y(n_1186)
);

INVx6_ASAP7_75t_L g1187 ( 
.A(n_1169),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1139),
.A2(n_1035),
.B1(n_1049),
.B2(n_1001),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1160),
.B(n_1083),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1139),
.A2(n_1095),
.B1(n_1082),
.B2(n_1050),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1149),
.A2(n_1001),
.B1(n_1082),
.B2(n_1079),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1126),
.A2(n_1001),
.B1(n_1027),
.B2(n_1041),
.Y(n_1192)
);

CKINVDCx11_ASAP7_75t_R g1193 ( 
.A(n_1114),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1127),
.Y(n_1194)
);

BUFx2_ASAP7_75t_SL g1195 ( 
.A(n_1114),
.Y(n_1195)
);

INVx6_ASAP7_75t_L g1196 ( 
.A(n_1169),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1134),
.Y(n_1197)
);

BUFx2_ASAP7_75t_SL g1198 ( 
.A(n_1142),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1126),
.A2(n_1001),
.B1(n_1042),
.B2(n_1095),
.Y(n_1199)
);

BUFx2_ASAP7_75t_SL g1200 ( 
.A(n_1142),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1133),
.A2(n_562),
.B1(n_914),
.B2(n_887),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1124),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1135),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1130),
.A2(n_1042),
.B1(n_1071),
.B2(n_1110),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1169),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1164),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1129),
.A2(n_1071),
.B1(n_1110),
.B2(n_1080),
.Y(n_1207)
);

CKINVDCx11_ASAP7_75t_R g1208 ( 
.A(n_1125),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1148),
.A2(n_1050),
.B1(n_1072),
.B2(n_1077),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1144),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1135),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1135),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1115),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1182),
.A2(n_1070),
.B1(n_1065),
.B2(n_948),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1141),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1147),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1182),
.A2(n_1065),
.B1(n_1086),
.B2(n_997),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1117),
.Y(n_1218)
);

CKINVDCx6p67_ASAP7_75t_R g1219 ( 
.A(n_1145),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1183),
.A2(n_598),
.B(n_595),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1150),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1151),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1138),
.A2(n_1065),
.B1(n_1086),
.B2(n_997),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1149),
.Y(n_1224)
);

CKINVDCx14_ASAP7_75t_R g1225 ( 
.A(n_1138),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1143),
.A2(n_598),
.B(n_595),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1145),
.A2(n_914),
.B1(n_1077),
.B2(n_937),
.Y(n_1227)
);

OAI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1122),
.A2(n_1072),
.B1(n_926),
.B2(n_942),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1181),
.A2(n_1057),
.B1(n_1030),
.B2(n_943),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1166),
.B(n_1167),
.Y(n_1230)
);

INVx6_ASAP7_75t_L g1231 ( 
.A(n_1131),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1111),
.Y(n_1232)
);

BUFx8_ASAP7_75t_L g1233 ( 
.A(n_1128),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1153),
.A2(n_1051),
.B(n_1028),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1178),
.A2(n_997),
.B1(n_1100),
.B2(n_1060),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1181),
.A2(n_997),
.B1(n_1105),
.B2(n_974),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1164),
.Y(n_1237)
);

INVx11_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1119),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1179),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1179),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_SL g1242 ( 
.A(n_1123),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1113),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1131),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1153),
.B(n_1096),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1132),
.A2(n_1018),
.B1(n_1030),
.B2(n_1052),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1135),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1116),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1136),
.B(n_1099),
.Y(n_1249)
);

INVx11_ASAP7_75t_L g1250 ( 
.A(n_1181),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1177),
.A2(n_961),
.B1(n_1029),
.B2(n_740),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1238),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1190),
.A2(n_1161),
.B1(n_1028),
.B2(n_1174),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1190),
.A2(n_1158),
.B1(n_1162),
.B2(n_1118),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1206),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1185),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1209),
.B(n_1161),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1249),
.B(n_1154),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1244),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1194),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1197),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_SL g1262 ( 
.A(n_1240),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1199),
.A2(n_1163),
.B1(n_1168),
.B2(n_1160),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1186),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1251),
.A2(n_1118),
.B1(n_1159),
.B2(n_1154),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1234),
.B(n_1096),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1188),
.A2(n_1173),
.B1(n_974),
.B2(n_1118),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1192),
.A2(n_987),
.B1(n_998),
.B2(n_976),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1207),
.A2(n_987),
.B1(n_998),
.B2(n_976),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1213),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1219),
.A2(n_1215),
.B1(n_1213),
.B2(n_1226),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1210),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1227),
.A2(n_1012),
.B1(n_1022),
.B2(n_1006),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1226),
.A2(n_949),
.B1(n_985),
.B2(n_983),
.Y(n_1274)
);

OR2x2_ASAP7_75t_SL g1275 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1220),
.A2(n_1051),
.B1(n_621),
.B2(n_628),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1229),
.A2(n_969),
.B1(n_997),
.B2(n_1159),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1234),
.B(n_1175),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1243),
.Y(n_1279)
);

INVx4_ASAP7_75t_SL g1280 ( 
.A(n_1187),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1237),
.B(n_1099),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1216),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1221),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1222),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1220),
.A2(n_621),
.B1(n_628),
.B2(n_618),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1227),
.A2(n_1006),
.B1(n_1022),
.B2(n_1012),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1191),
.A2(n_633),
.B1(n_638),
.B2(n_612),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1217),
.A2(n_646),
.B1(n_664),
.B2(n_618),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1237),
.B(n_995),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1245),
.B(n_1175),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1204),
.A2(n_1093),
.B1(n_953),
.B2(n_957),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1224),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1232),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1239),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1245),
.A2(n_1063),
.B(n_969),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1185),
.B(n_780),
.Y(n_1296)
);

AOI222xp33_ASAP7_75t_L g1297 ( 
.A1(n_1214),
.A2(n_638),
.B1(n_681),
.B2(n_633),
.C1(n_655),
.C2(n_612),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1223),
.A2(n_676),
.B(n_655),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1230),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1205),
.B(n_1225),
.Y(n_1300)
);

INVx5_ASAP7_75t_SL g1301 ( 
.A(n_1250),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1201),
.A2(n_1093),
.B1(n_953),
.B2(n_957),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1246),
.A2(n_1137),
.B1(n_1165),
.B2(n_1121),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1228),
.A2(n_1137),
.B1(n_1165),
.B2(n_1121),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1184),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1196),
.A2(n_681),
.B1(n_676),
.B2(n_1108),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1195),
.B(n_1017),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1235),
.A2(n_646),
.B1(n_666),
.B2(n_664),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1236),
.A2(n_692),
.B(n_666),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1202),
.A2(n_692),
.B1(n_697),
.B2(n_968),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1218),
.A2(n_697),
.B(n_569),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1211),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1203),
.B(n_1113),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1242),
.A2(n_1171),
.B1(n_975),
.B2(n_1011),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1265),
.A2(n_1233),
.B1(n_1208),
.B2(n_1200),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1287),
.A2(n_1297),
.B1(n_1302),
.B2(n_1267),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1290),
.B(n_1211),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1273),
.A2(n_1058),
.B1(n_1233),
.B2(n_1010),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1271),
.B(n_1285),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1286),
.A2(n_1016),
.B1(n_951),
.B2(n_557),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1253),
.A2(n_1198),
.B1(n_1231),
.B2(n_978),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1270),
.B(n_1212),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1285),
.A2(n_951),
.B1(n_557),
.B2(n_558),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1288),
.A2(n_557),
.B1(n_558),
.B2(n_1078),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1274),
.A2(n_1241),
.B1(n_979),
.B2(n_1193),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1275),
.A2(n_1202),
.B1(n_979),
.B2(n_960),
.Y(n_1326)
);

NAND4xp25_ASAP7_75t_L g1327 ( 
.A(n_1274),
.B(n_569),
.C(n_988),
.D(n_1023),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1291),
.A2(n_1007),
.B1(n_652),
.B2(n_656),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1253),
.A2(n_1020),
.B1(n_1231),
.B2(n_1203),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1007),
.B1(n_652),
.B2(n_656),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1268),
.A2(n_680),
.B1(n_691),
.B2(n_651),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1257),
.B(n_1203),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1290),
.B(n_1247),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1295),
.A2(n_1063),
.B(n_597),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1306),
.A2(n_1248),
.B1(n_1170),
.B2(n_1172),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_680),
.B1(n_691),
.B2(n_651),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1254),
.A2(n_651),
.B1(n_1094),
.B2(n_1017),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1276),
.A2(n_1108),
.B1(n_1189),
.B2(n_606),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1308),
.A2(n_1276),
.B1(n_1269),
.B2(n_1299),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1308),
.A2(n_1094),
.B1(n_1009),
.B2(n_1036),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1293),
.B(n_1112),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1281),
.A2(n_1009),
.B1(n_1054),
.B2(n_1026),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1310),
.A2(n_1009),
.B1(n_1020),
.B2(n_608),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1310),
.A2(n_1009),
.B1(n_1020),
.B2(n_608),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_1278),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1307),
.A2(n_1009),
.B1(n_1020),
.B2(n_608),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1304),
.A2(n_619),
.B1(n_620),
.B2(n_606),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1314),
.A2(n_620),
.B1(n_645),
.B2(n_619),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1277),
.A2(n_1298),
.B1(n_1309),
.B2(n_1263),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1264),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1296),
.A2(n_1170),
.B1(n_1172),
.B2(n_1155),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1255),
.B(n_1189),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1266),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1260),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1261),
.B(n_72),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1311),
.B(n_1106),
.C(n_591),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1266),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1278),
.A2(n_620),
.B1(n_645),
.B2(n_619),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1295),
.A2(n_996),
.B(n_977),
.Y(n_1359)
);

OAI222xp33_ASAP7_75t_L g1360 ( 
.A1(n_1272),
.A2(n_1283),
.B1(n_1284),
.B2(n_1282),
.C1(n_1294),
.C2(n_1258),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1312),
.Y(n_1361)
);

AND4x1_ASAP7_75t_L g1362 ( 
.A(n_1300),
.B(n_988),
.C(n_75),
.D(n_74),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1279),
.B(n_1113),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1256),
.A2(n_1066),
.B1(n_1097),
.B2(n_1176),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1292),
.A2(n_1180),
.B1(n_1176),
.B2(n_1116),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1280),
.A2(n_650),
.B1(n_645),
.B2(n_986),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1313),
.A2(n_1002),
.B(n_1003),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1280),
.A2(n_986),
.B1(n_973),
.B2(n_967),
.Y(n_1368)
);

AOI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1280),
.A2(n_973),
.B1(n_964),
.B2(n_970),
.C1(n_967),
.C2(n_649),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1279),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1305),
.B(n_1146),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1259),
.A2(n_650),
.B1(n_1108),
.B2(n_649),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1259),
.A2(n_1108),
.B1(n_649),
.B2(n_1004),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1301),
.A2(n_1034),
.B1(n_617),
.B2(n_1146),
.Y(n_1374)
);

OAI222xp33_ASAP7_75t_L g1375 ( 
.A1(n_1262),
.A2(n_626),
.B1(n_1180),
.B2(n_453),
.C1(n_1152),
.C2(n_1156),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1252),
.A2(n_585),
.B1(n_590),
.B2(n_626),
.C(n_708),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1252),
.A2(n_1146),
.B1(n_626),
.B2(n_1157),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1332),
.A2(n_338),
.B(n_590),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_1157),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1333),
.B(n_1354),
.Y(n_1381)
);

OAI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_1362),
.A2(n_1319),
.B1(n_1316),
.B2(n_1325),
.C(n_1327),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1319),
.A2(n_1097),
.B(n_1156),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1349),
.A2(n_1157),
.B1(n_1107),
.B2(n_1092),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1339),
.A2(n_338),
.B1(n_1157),
.B2(n_590),
.Y(n_1385)
);

OAI221xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1321),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.C(n_80),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1322),
.B(n_76),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1356),
.B(n_1062),
.C(n_1055),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1062),
.C(n_1055),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1355),
.B(n_78),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1355),
.B(n_81),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1357),
.B(n_82),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1357),
.B(n_83),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1332),
.B(n_84),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1361),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1341),
.B(n_1371),
.C(n_1370),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1352),
.B(n_87),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1360),
.B(n_89),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1329),
.B(n_1062),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1315),
.A2(n_89),
.B(n_90),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1368),
.A2(n_1323),
.B1(n_1338),
.B2(n_1343),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1359),
.B(n_91),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1359),
.B(n_91),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_338),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1359),
.B(n_338),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1344),
.A2(n_1107),
.B1(n_1092),
.B2(n_1069),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1358),
.A2(n_963),
.B(n_1069),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1351),
.B(n_1107),
.C(n_963),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_963),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1375),
.A2(n_94),
.B(n_95),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_315),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1350),
.B(n_98),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1334),
.B(n_100),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1350),
.B(n_103),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1334),
.B(n_105),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1336),
.B(n_107),
.C(n_109),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1334),
.B(n_111),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1340),
.B(n_314),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_312),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1395),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1380),
.B(n_1335),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1381),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1400),
.B(n_1382),
.C(n_1386),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_L g1424 ( 
.A1(n_1394),
.A2(n_1373),
.B(n_1318),
.C(n_1377),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1396),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1394),
.B(n_1324),
.C(n_1376),
.Y(n_1426)
);

NOR3xp33_ASAP7_75t_SL g1427 ( 
.A(n_1410),
.B(n_1326),
.C(n_1365),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1402),
.Y(n_1428)
);

OAI211xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1397),
.A2(n_1369),
.B(n_1342),
.C(n_1372),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1404),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1387),
.A2(n_1346),
.B(n_1364),
.C(n_1366),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1384),
.B(n_1374),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1379),
.B(n_1337),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1403),
.B(n_1330),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1392),
.B(n_1320),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1398),
.A2(n_1348),
.B1(n_1347),
.B2(n_1331),
.C(n_1328),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1398),
.B(n_120),
.C(n_121),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1405),
.Y(n_1438)
);

NAND4xp75_ASAP7_75t_L g1439 ( 
.A(n_1399),
.B(n_130),
.C(n_132),
.D(n_133),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1393),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1401),
.A2(n_135),
.B1(n_140),
.B2(n_144),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1383),
.B(n_1409),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1390),
.B(n_146),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1405),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_1444)
);

AOI211x1_ASAP7_75t_L g1445 ( 
.A1(n_1391),
.A2(n_153),
.B(n_154),
.C(n_157),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1389),
.B(n_158),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1425),
.Y(n_1447)
);

NOR2x1_ASAP7_75t_L g1448 ( 
.A(n_1440),
.B(n_1408),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1438),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1428),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1438),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1422),
.B(n_1378),
.Y(n_1452)
);

AND2x4_ASAP7_75t_SL g1453 ( 
.A(n_1442),
.B(n_1411),
.Y(n_1453)
);

NAND4xp75_ASAP7_75t_SL g1454 ( 
.A(n_1443),
.B(n_1378),
.C(n_1407),
.D(n_1417),
.Y(n_1454)
);

XOR2x2_ASAP7_75t_L g1455 ( 
.A(n_1423),
.B(n_1385),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1421),
.B(n_1378),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1443),
.B(n_1388),
.Y(n_1459)
);

NOR4xp25_ASAP7_75t_L g1460 ( 
.A(n_1441),
.B(n_1385),
.C(n_1399),
.D(n_1418),
.Y(n_1460)
);

XOR2xp5_ASAP7_75t_L g1461 ( 
.A(n_1433),
.B(n_1412),
.Y(n_1461)
);

NAND4xp75_ASAP7_75t_SL g1462 ( 
.A(n_1423),
.B(n_1407),
.C(n_1415),
.D(n_1413),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1434),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1435),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1458),
.Y(n_1465)
);

XOR2x2_ASAP7_75t_L g1466 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1466)
);

AO22x2_ASAP7_75t_L g1467 ( 
.A1(n_1447),
.A2(n_1445),
.B1(n_1424),
.B2(n_1426),
.Y(n_1467)
);

XNOR2x1_ASAP7_75t_L g1468 ( 
.A(n_1455),
.B(n_1439),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1448),
.Y(n_1469)
);

XOR2x2_ASAP7_75t_L g1470 ( 
.A(n_1461),
.B(n_1441),
.Y(n_1470)
);

CKINVDCx8_ASAP7_75t_R g1471 ( 
.A(n_1459),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1452),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1453),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1463),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1451),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1464),
.B(n_1429),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1451),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1471),
.A2(n_1469),
.B1(n_1467),
.B2(n_1468),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1475),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1474),
.Y(n_1480)
);

XNOR2x1_ASAP7_75t_L g1481 ( 
.A(n_1466),
.B(n_1462),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_SL g1482 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1482)
);

OA22x2_ASAP7_75t_L g1483 ( 
.A1(n_1469),
.A2(n_1450),
.B1(n_1432),
.B2(n_1456),
.Y(n_1483)
);

AO22x1_ASAP7_75t_L g1484 ( 
.A1(n_1476),
.A2(n_1460),
.B1(n_1454),
.B2(n_1427),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1475),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1467),
.A2(n_1457),
.B1(n_1427),
.B2(n_1431),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1470),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1467),
.A2(n_1444),
.B1(n_1446),
.B2(n_1419),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1472),
.A2(n_1444),
.B1(n_1436),
.B2(n_1414),
.Y(n_1489)
);

OA22x2_ASAP7_75t_L g1490 ( 
.A1(n_1477),
.A2(n_1406),
.B1(n_1416),
.B2(n_164),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1465),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1478),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1488),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1491),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1479),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1485),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1489),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1486),
.Y(n_1499)
);

OA22x2_ASAP7_75t_L g1500 ( 
.A1(n_1493),
.A2(n_1487),
.B1(n_1481),
.B2(n_1484),
.Y(n_1500)
);

AND4x1_ASAP7_75t_L g1501 ( 
.A(n_1499),
.B(n_1482),
.C(n_1490),
.D(n_1483),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1494),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1495),
.Y(n_1503)
);

OA22x2_ASAP7_75t_L g1504 ( 
.A1(n_1498),
.A2(n_193),
.B1(n_197),
.B2(n_199),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1497),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1492),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1503),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1502),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1500),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1506),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1504),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1505),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1501),
.B(n_1496),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1513),
.A2(n_1509),
.B1(n_1511),
.B2(n_1512),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1508),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1510),
.B(n_202),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1507),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1517),
.B(n_310),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1514),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1515),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1516),
.B(n_209),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1520),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1518),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1519),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_1524)
);

BUFx2_ASAP7_75t_SL g1525 ( 
.A(n_1521),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1521),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1526),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1525),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1523),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1522),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1524),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1522),
.A2(n_218),
.B1(n_222),
.B2(n_224),
.Y(n_1532)
);

BUFx4f_ASAP7_75t_SL g1533 ( 
.A(n_1522),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1526),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1527),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_1535)
);

AND4x2_ASAP7_75t_L g1536 ( 
.A(n_1533),
.B(n_231),
.C(n_232),
.D(n_233),
.Y(n_1536)
);

AO22x2_ASAP7_75t_L g1537 ( 
.A1(n_1528),
.A2(n_234),
.B1(n_240),
.B2(n_243),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1534),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1531),
.A2(n_252),
.B1(n_258),
.B2(n_260),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1530),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1529),
.A2(n_261),
.B1(n_262),
.B2(n_266),
.Y(n_1541)
);

OAI22x1_ASAP7_75t_L g1542 ( 
.A1(n_1532),
.A2(n_267),
.B1(n_268),
.B2(n_271),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1540),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1537),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1537),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1542),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1536),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1547),
.A2(n_1539),
.B1(n_1538),
.B2(n_1535),
.Y(n_1548)
);

OAI22x1_ASAP7_75t_L g1549 ( 
.A1(n_1543),
.A2(n_1541),
.B1(n_274),
.B2(n_279),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1549),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1548),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1550),
.A2(n_1544),
.B1(n_1545),
.B2(n_1546),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1551),
.A2(n_280),
.B1(n_285),
.B2(n_288),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1552),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1553),
.B(n_289),
.Y(n_1555)
);

AOI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1554),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.C(n_297),
.Y(n_1556)
);

AOI211xp5_ASAP7_75t_L g1557 ( 
.A1(n_1556),
.A2(n_1555),
.B(n_303),
.C(n_304),
.Y(n_1557)
);


endmodule