module fake_jpeg_3635_n_226 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_18),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_63),
.B1(n_80),
.B2(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_0),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_0),
.Y(n_89)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_58),
.B(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_66),
.B1(n_79),
.B2(n_78),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_76),
.B1(n_75),
.B2(n_69),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_78),
.B1(n_87),
.B2(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_57),
.B1(n_80),
.B2(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_76),
.B1(n_75),
.B2(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_56),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_84),
.B1(n_82),
.B2(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_120),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_89),
.B1(n_82),
.B2(n_62),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_112),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_118),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_64),
.C(n_65),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_91),
.B(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_88),
.B1(n_60),
.B2(n_77),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_123),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_72),
.B1(n_71),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_94),
.B1(n_96),
.B2(n_69),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_139),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_134),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_1),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_115),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_2),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_2),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_7),
.Y(n_167)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_81),
.B1(n_70),
.B2(n_6),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_159),
.B1(n_162),
.B2(n_171),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_125),
.B(n_131),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_36),
.C(n_26),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_163),
.C(n_162),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_81),
.B1(n_70),
.B2(n_50),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_81),
.B1(n_70),
.B2(n_49),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_167),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_44),
.C(n_43),
.Y(n_163)
);

XOR2x2_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_7),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_40),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_177),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_170),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_151),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_128),
.B(n_131),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_189),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_125),
.B(n_37),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_125),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_198),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_184),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_158),
.B1(n_150),
.B2(n_171),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_209)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_192),
.A3(n_200),
.B1(n_193),
.B2(n_197),
.C1(n_191),
.C2(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_172),
.A3(n_189),
.B1(n_182),
.B2(n_177),
.C1(n_176),
.C2(n_185),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_154),
.B(n_159),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_27),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_186),
.A3(n_164),
.B1(n_175),
.B2(n_179),
.C1(n_147),
.C2(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_15),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_206),
.B(n_209),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_213),
.B(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_214),
.C(n_28),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_219),
.B1(n_31),
.B2(n_33),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_24),
.Y(n_223)
);

OAI321xp33_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_34),
.A3(n_35),
.B1(n_21),
.B2(n_22),
.C(n_19),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_19),
.B(n_20),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_21),
.Y(n_226)
);


endmodule