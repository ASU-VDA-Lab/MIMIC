module fake_jpeg_12509_n_164 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_14),
.A2(n_2),
.B(n_4),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_50),
.B(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_52),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_13),
.Y(n_59)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_22),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_64),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_12),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_26),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_20),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_10),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_60),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_92),
.B(n_102),
.C(n_104),
.D(n_81),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_72),
.C(n_57),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_63),
.B1(n_70),
.B2(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_101),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_72),
.B1(n_75),
.B2(n_69),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_62),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_82),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_78),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_79),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_79),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_79),
.B1(n_81),
.B2(n_88),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_97),
.B1(n_102),
.B2(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_129),
.B(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_131),
.Y(n_142)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_115),
.B1(n_105),
.B2(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_135),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_121),
.B(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_107),
.B(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_111),
.B1(n_117),
.B2(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_127),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_149),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_140),
.B(n_130),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_149),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_145),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_154),
.A2(n_157),
.B(n_153),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_133),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_129),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.C(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_142),
.Y(n_163)
);

NAND2x1_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_143),
.Y(n_164)
);


endmodule