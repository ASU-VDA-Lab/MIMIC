module fake_jpeg_14765_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_21),
.B1(n_27),
.B2(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_30),
.B2(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_28),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_44),
.B1(n_51),
.B2(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_15),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_59),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_37),
.B1(n_31),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_50),
.B1(n_45),
.B2(n_34),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_42),
.B(n_43),
.C(n_47),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_20),
.B(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_69),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_27),
.B(n_33),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_72),
.C(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_50),
.B1(n_45),
.B2(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_15),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_97),
.B1(n_73),
.B2(n_17),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_98),
.B(n_101),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_73),
.B1(n_60),
.B2(n_80),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_36),
.A3(n_35),
.B1(n_34),
.B2(n_26),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_95),
.B(n_65),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_35),
.B1(n_22),
.B2(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_22),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_106),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_124),
.B1(n_58),
.B2(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_114),
.Y(n_141)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_69),
.C(n_72),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_113),
.C(n_67),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_102),
.C(n_86),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_121),
.B(n_123),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_118),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_119),
.B(n_15),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_57),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_70),
.B1(n_76),
.B2(n_74),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_94),
.B1(n_79),
.B2(n_88),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_76),
.C(n_0),
.D(n_2),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_93),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_76),
.B(n_67),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_16),
.B1(n_15),
.B2(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_132),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_97),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_138),
.C(n_120),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_90),
.B1(n_81),
.B2(n_80),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_133),
.B1(n_122),
.B2(n_108),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_146),
.B1(n_123),
.B2(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_87),
.B1(n_96),
.B2(n_16),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_140),
.B1(n_145),
.B2(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_87),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_147),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_15),
.B(n_1),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_143),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_58),
.B1(n_93),
.B2(n_0),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_9),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_114),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_108),
.B1(n_123),
.B2(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_112),
.C(n_111),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_113),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_162),
.C(n_139),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_113),
.C(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_10),
.C(n_2),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_128),
.B1(n_141),
.B2(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_0),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_14),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_143),
.B(n_131),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_109),
.B(n_3),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_130),
.B1(n_145),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_152),
.B1(n_145),
.B2(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_150),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_168),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_172),
.C(n_166),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_182),
.C(n_184),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_156),
.C(n_157),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_164),
.B1(n_149),
.B2(n_153),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_186),
.B(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_148),
.C(n_165),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_13),
.Y(n_198)
);

OA21x2_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_9),
.B(n_4),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_168),
.C(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_13),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_176),
.C(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_196),
.C(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_198),
.B1(n_6),
.B2(n_11),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_184),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_185),
.B1(n_183),
.B2(n_170),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_200),
.B(n_204),
.C(n_191),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_203),
.B(n_190),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_179),
.A3(n_169),
.B1(n_170),
.B2(n_175),
.C1(n_6),
.C2(n_11),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_209),
.B(n_12),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_196),
.B(n_192),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_208),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_192),
.B(n_190),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_6),
.C(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_0),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_213),
.Y(n_216)
);


endmodule