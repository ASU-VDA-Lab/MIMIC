module fake_jpeg_3434_n_392 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_45),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_51),
.B(n_54),
.Y(n_128)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_6),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_15),
.B(n_6),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_0),
.CON(n_65),
.SN(n_65)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_84),
.B(n_1),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_72),
.Y(n_119)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_9),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_74),
.B(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_10),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_93),
.Y(n_136)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_10),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_19),
.Y(n_144)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_19),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_26),
.B1(n_31),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_141),
.B1(n_149),
.B2(n_65),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_31),
.B1(n_41),
.B2(n_22),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_100),
.A2(n_104),
.B1(n_117),
.B2(n_118),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_39),
.B1(n_27),
.B2(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_27),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_130),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_108),
.A2(n_107),
.B(n_129),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_39),
.B1(n_42),
.B2(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_42),
.B1(n_28),
.B2(n_23),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_92),
.B1(n_94),
.B2(n_60),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_143),
.B1(n_25),
.B2(n_2),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_28),
.C(n_42),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_12),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_53),
.A2(n_19),
.B1(n_42),
.B2(n_28),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_48),
.A2(n_19),
.B1(n_42),
.B2(n_25),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_53),
.A2(n_25),
.B1(n_11),
.B2(n_3),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_81),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_57),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_152),
.B(n_166),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_163),
.Y(n_203)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_161),
.A2(n_112),
.B1(n_131),
.B2(n_142),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_87),
.B1(n_76),
.B2(n_75),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_179),
.B1(n_131),
.B2(n_137),
.Y(n_216)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_52),
.B(n_73),
.C(n_91),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_99),
.A3(n_119),
.B1(n_101),
.B2(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_101),
.A2(n_61),
.B1(n_58),
.B2(n_56),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_175),
.B1(n_124),
.B2(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_183),
.Y(n_204)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_181),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_189),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_182),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_25),
.B1(n_12),
.B2(n_4),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_103),
.A2(n_5),
.B(n_12),
.C(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_186),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_5),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_139),
.A2(n_5),
.B(n_14),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_134),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_192),
.Y(n_213)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_112),
.B1(n_121),
.B2(n_131),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_2),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_111),
.B(n_2),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_216),
.B1(n_225),
.B2(n_205),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_126),
.B1(n_122),
.B2(n_139),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_205),
.B1(n_223),
.B2(n_155),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_113),
.B1(n_140),
.B2(n_102),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_215),
.C(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_177),
.C(n_152),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_148),
.C(n_111),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_160),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_190),
.B1(n_181),
.B2(n_140),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_113),
.B1(n_137),
.B2(n_106),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_192),
.B(n_132),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_168),
.B1(n_166),
.B2(n_189),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_228),
.A2(n_245),
.B1(n_217),
.B2(n_209),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_231),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_184),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_218),
.C(n_208),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_194),
.B(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_170),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_194),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_251),
.B1(n_252),
.B2(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_183),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_153),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_247),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_198),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_188),
.B1(n_178),
.B2(n_169),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_180),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_191),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_202),
.B1(n_206),
.B2(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_207),
.A2(n_135),
.B1(n_102),
.B2(n_106),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_262),
.C(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_219),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_260),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_204),
.C(n_208),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_237),
.B1(n_228),
.B2(n_245),
.Y(n_287)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_219),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_227),
.B(n_197),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_229),
.B(n_253),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_209),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_251),
.B1(n_250),
.B2(n_228),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_212),
.C(n_182),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_159),
.C(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_221),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_277),
.Y(n_293)
);

AOI21x1_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_231),
.B(n_235),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_278),
.A2(n_283),
.B(n_295),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_299),
.B1(n_298),
.B2(n_266),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_289),
.C(n_265),
.Y(n_302)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_259),
.B(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_241),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_285),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_234),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_290),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_288),
.B1(n_297),
.B2(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_245),
.B1(n_247),
.B2(n_239),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_232),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_244),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_298),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_274),
.B1(n_258),
.B2(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_242),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_252),
.B1(n_253),
.B2(n_233),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_307),
.B1(n_271),
.B2(n_291),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_311),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_284),
.B1(n_292),
.B2(n_282),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_281),
.A2(n_274),
.B1(n_255),
.B2(n_259),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_262),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.C(n_316),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_259),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_222),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_286),
.B(n_285),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_315),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_294),
.C(n_280),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_268),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_264),
.C(n_268),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_319),
.C(n_283),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_279),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_269),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_299),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_328),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_337),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_318),
.B1(n_320),
.B2(n_309),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_SL g327 ( 
.A1(n_302),
.A2(n_295),
.B(n_278),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_310),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_269),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_222),
.C(n_246),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_334),
.C(n_335),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_221),
.B(n_199),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_330),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_304),
.B1(n_300),
.B2(n_319),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_199),
.C(n_197),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_211),
.C(n_214),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_226),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_335),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_351),
.Y(n_356)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_317),
.B1(n_310),
.B2(n_303),
.Y(n_346)
);

AO221x1_ASAP7_75t_L g359 ( 
.A1(n_346),
.A2(n_253),
.B1(n_214),
.B2(n_211),
.C(n_132),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_328),
.C(n_334),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_348),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_323),
.B(n_301),
.CI(n_306),
.CON(n_348),
.SN(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_195),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_349),
.B(n_337),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_211),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_321),
.C(n_322),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_354),
.Y(n_364)
);

OAI321xp33_ASAP7_75t_L g355 ( 
.A1(n_340),
.A2(n_332),
.A3(n_350),
.B1(n_338),
.B2(n_351),
.C(n_344),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_346),
.B1(n_348),
.B2(n_342),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_322),
.C(n_332),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_361),
.Y(n_367)
);

NAND2x1_ASAP7_75t_SL g363 ( 
.A(n_359),
.B(n_348),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_SL g360 ( 
.A1(n_351),
.A2(n_195),
.B(n_132),
.C(n_185),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_356),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_158),
.C(n_156),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_368),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_366),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_341),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_362),
.A2(n_356),
.B(n_339),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_369),
.A2(n_360),
.B(n_157),
.Y(n_375)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_360),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_374),
.B(n_376),
.Y(n_381)
);

AOI21xp33_ASAP7_75t_L g379 ( 
.A1(n_375),
.A2(n_377),
.B(n_368),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_364),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_360),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_165),
.B(n_187),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_378),
.A2(n_173),
.B(n_142),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_373),
.B(n_363),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_382),
.B(n_383),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_369),
.B(n_162),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_377),
.B(n_171),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_386),
.A2(n_387),
.B(n_173),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_SL g387 ( 
.A1(n_380),
.A2(n_173),
.B(n_14),
.C(n_147),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_176),
.Y(n_388)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_389),
.A3(n_147),
.B1(n_109),
.B2(n_116),
.C1(n_135),
.C2(n_385),
.Y(n_390)
);

NOR3xp33_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_109),
.C(n_116),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_114),
.B1(n_147),
.B2(n_14),
.Y(n_392)
);


endmodule