module fake_jpeg_2474_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx2_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_51),
.Y(n_58)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_33),
.B1(n_15),
.B2(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_0),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_36),
.B1(n_46),
.B2(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_53),
.B(n_41),
.C(n_43),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_74),
.B(n_38),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_36),
.B(n_44),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_61),
.B1(n_60),
.B2(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_80),
.B1(n_0),
.B2(n_1),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_81),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_46),
.B1(n_44),
.B2(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_42),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_39),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_32),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_73),
.B(n_38),
.C(n_71),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_9),
.B(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_99),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_21),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_2),
.B(n_3),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_97),
.B(n_102),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_88),
.B1(n_10),
.B2(n_11),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_5),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_12),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_88),
.C(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_9),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_104),
.C(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_109),
.B1(n_104),
.B2(n_27),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_113),
.B1(n_116),
.B2(n_109),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_127),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_120),
.B1(n_125),
.B2(n_123),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_129),
.B1(n_118),
.B2(n_117),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_126),
.B(n_25),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_22),
.C(n_28),
.Y(n_133)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_30),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_31),
.Y(n_136)
);


endmodule