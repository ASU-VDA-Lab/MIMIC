module real_jpeg_26377_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_5),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_152),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_152),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_152),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_7),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_7),
.A2(n_31),
.B1(n_122),
.B2(n_150),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_150),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_150),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_8),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_105),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_52),
.C(n_55),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_83),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_8),
.A2(n_88),
.B1(n_229),
.B2(n_232),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_10),
.A2(n_32),
.B1(n_42),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_10),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_159),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_159),
.Y(n_229)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_12),
.A2(n_68),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_14),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_14),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_139)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_106),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_84),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_20),
.A2(n_71),
.B1(n_72),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_20),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_43),
.B2(n_44),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_21),
.A2(n_22),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_45),
.C(n_61),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_34),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_23),
.A2(n_101),
.B1(n_158),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_29),
.B1(n_39),
.B2(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_24),
.A2(n_27),
.B(n_156),
.C(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_26),
.A2(n_27),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_26),
.B(n_29),
.C(n_32),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_26),
.B(n_50),
.C(n_64),
.Y(n_245)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g244 ( 
.A(n_27),
.B(n_155),
.CON(n_244),
.SN(n_244)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_30),
.Y(n_118)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_32),
.B(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_35),
.B(n_105),
.Y(n_104)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_39),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_40),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_40),
.A2(n_105),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_40),
.A2(n_105),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_40),
.A2(n_105),
.B1(n_165),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_45),
.A2(n_46),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_47),
.A2(n_54),
.B1(n_205),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_47),
.A2(n_74),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_49),
.A2(n_65),
.B(n_243),
.C(n_245),
.Y(n_242)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_50),
.B(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_79),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_54),
.A2(n_76),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_54),
.B(n_155),
.Y(n_227)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_56),
.B(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_58),
.A2(n_77),
.B(n_98),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_69),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_67),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_62),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_62),
.A2(n_83),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_62),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_62),
.A2(n_83),
.B1(n_191),
.B2(n_244),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_62),
.A2(n_69),
.B(n_114),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_66),
.A2(n_168),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_66),
.A2(n_82),
.B(n_115),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_72),
.A2(n_73),
.B(n_80),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_75),
.A2(n_77),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_75),
.A2(n_77),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_75),
.A2(n_77),
.B1(n_96),
.B2(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_84),
.B(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_99),
.B(n_100),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_85),
.A2(n_86),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_87),
.A2(n_94),
.B1(n_99),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_87),
.A2(n_99),
.B1(n_100),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_93),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_88),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_88),
.A2(n_141),
.B1(n_222),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_88),
.A2(n_93),
.B(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_89),
.A2(n_137),
.B1(n_140),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_89),
.B(n_139),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_89),
.A2(n_210),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_91),
.B(n_155),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_100),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_104),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_101),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_103),
.B(n_105),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_328),
.B(n_333),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_313),
.B(n_327),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_294),
.B(n_312),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_193),
.B(n_276),
.C(n_293),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_177),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_132),
.B(n_177),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_160),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_146),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_134),
.B(n_146),
.C(n_160),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_135),
.B(n_144),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_143),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_145),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_153),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_179),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_169),
.B2(n_176),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_163),
.B(n_166),
.C(n_176),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_184),
.B(n_186),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_178),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_180),
.B(n_182),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_186),
.B(n_209),
.Y(n_282)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_275),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_270),
.B(n_274),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_255),
.B(n_269),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_238),
.B(n_254),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_218),
.B(n_237),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_202),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_213),
.C(n_216),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_217),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_225),
.B(n_236),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_230),
.B(n_235),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_253),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_253),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_248),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_249),
.C(n_250),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_247),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_265),
.C(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_292),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_286),
.C(n_292),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_285),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_296),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_311),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_309),
.B2(n_310),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_310),
.C(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_306),
.C(n_308),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_322),
.B2(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_322),
.C(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);


endmodule