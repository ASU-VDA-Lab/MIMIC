module real_jpeg_30593_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx3_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_0),
.A2(n_47),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g162 ( 
.A1(n_0),
.A2(n_47),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_0),
.B(n_25),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_0),
.A2(n_47),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_0),
.A2(n_260),
.A3(n_265),
.B1(n_268),
.B2(n_276),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_0),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_0),
.B(n_155),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_1),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g412 ( 
.A(n_1),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_2),
.B(n_219),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_2),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_102),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_6),
.A2(n_102),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22x1_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_39),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_39),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_9),
.A2(n_39),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_11),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_11),
.A2(n_86),
.B1(n_173),
.B2(n_177),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_86),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_13),
.Y(n_219)
);

OAI211xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_220),
.B(n_467),
.C(n_469),
.Y(n_14)
);

NAND2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_217),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_16),
.B(n_218),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_215),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_193),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_18),
.B(n_193),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.C(n_156),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_19),
.A2(n_20),
.B1(n_132),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_59),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_21),
.B(n_317),
.C(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_22),
.A2(n_23),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_23),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_43),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g191 ( 
.A(n_24),
.B(n_192),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_24),
.A2(n_35),
.B1(n_192),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_52),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_32),
.Y(n_141)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_33),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_38),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_44),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_44),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_47),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_47),
.B(n_329),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_47),
.A2(n_64),
.B(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_47),
.B(n_90),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_48),
.B(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_51),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_58),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_88),
.B2(n_131),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_60),
.B(n_131),
.C(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_60),
.B(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_83),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_62),
.B(n_318),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_70),
.C(n_78),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_64),
.A2(n_70),
.B(n_79),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_66),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_70)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_70),
.A2(n_146),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_71),
.Y(n_244)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_72),
.Y(n_339)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_74),
.Y(n_358)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_145),
.B1(n_154),
.B2(n_155),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_85),
.Y(n_330)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_100),
.B(n_113),
.Y(n_88)
);

HB1xp67_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_120),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_135),
.B1(n_142),
.B2(n_143),
.Y(n_134)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_90),
.A2(n_142),
.B(n_143),
.Y(n_417)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_93),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_101),
.A2(n_119),
.B1(n_206),
.B2(n_213),
.Y(n_205)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

AOI22x1_ASAP7_75t_L g320 ( 
.A1(n_114),
.A2(n_119),
.B1(n_136),
.B2(n_213),
.Y(n_320)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_117),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_117),
.Y(n_299)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_130),
.Y(n_275)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_132),
.Y(n_463)
);

HB1xp67_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_133),
.B(n_452),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_134),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_144),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_153),
.Y(n_255)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g247 ( 
.A1(n_154),
.A2(n_155),
.B1(n_248),
.B2(n_256),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g341 ( 
.A1(n_154),
.A2(n_155),
.B1(n_256),
.B2(n_342),
.Y(n_341)
);

XOR2x2_ASAP7_75t_L g461 ( 
.A(n_156),
.B(n_462),
.Y(n_461)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_188),
.B(n_189),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_158),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_171),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_159),
.A2(n_171),
.B1(n_188),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_159),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_161),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_162),
.Y(n_256)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_166),
.Y(n_267)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_171),
.B(n_190),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_172),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_175),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_179),
.B(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_180),
.A2(n_387),
.B1(n_409),
.B2(n_413),
.Y(n_408)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_181),
.A2(n_236),
.B1(n_241),
.B2(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_187),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_187),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_195),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_195),
.B(n_418),
.C(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_214),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_201),
.A2(n_202),
.B1(n_319),
.B2(n_320),
.Y(n_440)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_202),
.B(n_227),
.Y(n_397)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_217),
.B(n_470),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_220),
.B(n_468),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_459),
.B(n_466),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_423),
.B(n_456),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_377),
.Y(n_222)
);

OAI21x1_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_322),
.B(n_376),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_283),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_225),
.B(n_283),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_246),
.C(n_257),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_226),
.B(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_227),
.B(n_230),
.C(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_227),
.B(n_420),
.C(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_227),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B(n_245),
.Y(n_229)
);

OAI211xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_232),
.B(n_235),
.C(n_240),
.Y(n_245)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_231),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_231),
.B(n_354),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_235),
.B(n_240),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_240),
.A2(n_387),
.B(n_393),
.Y(n_386)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_246),
.A2(n_247),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_246),
.B(n_308),
.C(n_346),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_246),
.A2(n_257),
.B1(n_258),
.B2(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_246),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_246),
.B(n_408),
.Y(n_439)
);

INVx3_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_247),
.Y(n_374)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_282),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_259),
.B(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_315),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_312),
.B2(n_313),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_285),
.B(n_315),
.C(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_308),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_287),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_291),
.B(n_300),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_308),
.B(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_360),
.Y(n_361)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_349),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_320),
.B1(n_340),
.B2(n_351),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_319),
.B(n_340),
.C(n_367),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_320),
.B(n_422),
.C(n_447),
.Y(n_446)
);

AOI21x1_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_370),
.B(n_375),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_364),
.B(n_369),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_347),
.B(n_363),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_343),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g363 ( 
.A(n_326),
.B(n_343),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_340),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_340),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_331),
.B(n_335),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_351),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_386),
.Y(n_418)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI21x1_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_352),
.B(n_362),
.Y(n_347)
);

AOI21x1_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_359),
.B(n_361),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_366),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_372),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_398),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_381),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_394),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_402),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_402),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_394),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B(n_403),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_404),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_419),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_414),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_431),
.C(n_432),
.Y(n_430)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_410),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND4xp25_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.C(n_429),
.D(n_444),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_433),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_438),
.C(n_441),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_441),
.B2(n_442),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_444),
.A2(n_457),
.B(n_458),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_454),
.B(n_455),
.Y(n_444)
);

NOR3xp33_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_454),
.C(n_455),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_448),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_451),
.C(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_449),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_460),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_464),
.Y(n_466)
);


endmodule