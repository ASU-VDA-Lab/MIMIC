module real_aes_8614_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_241;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g434 ( .A(n_0), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_1), .A2(n_120), .B(n_123), .C(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g186 ( .A(n_2), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_3), .A2(n_115), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_4), .B(n_196), .Y(n_513) );
AOI21xp33_ASAP7_75t_L g197 ( .A1(n_5), .A2(n_115), .B(n_198), .Y(n_197) );
AND2x6_ASAP7_75t_L g120 ( .A(n_6), .B(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_7), .A2(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_8), .B(n_41), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_9), .A2(n_31), .B1(n_104), .B2(n_105), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g448 ( .A(n_10), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_11), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g203 ( .A(n_12), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_13), .B(n_156), .Y(n_469) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
INVx1_ASAP7_75t_L g174 ( .A(n_15), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_16), .A2(n_129), .B(n_175), .C(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_17), .B(n_196), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_18), .B(n_131), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_19), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_20), .B(n_549), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_21), .A2(n_155), .B(n_189), .C(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_22), .B(n_196), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_23), .B(n_156), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_24), .A2(n_171), .B(n_173), .C(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_25), .B(n_156), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_26), .Y(n_498) );
INVx1_ASAP7_75t_L g487 ( .A(n_27), .Y(n_487) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_29), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_30), .B(n_156), .Y(n_187) );
INVx1_ASAP7_75t_L g104 ( .A(n_31), .Y(n_104) );
INVx1_ASAP7_75t_L g545 ( .A(n_32), .Y(n_545) );
INVx1_ASAP7_75t_L g213 ( .A(n_33), .Y(n_213) );
INVx2_ASAP7_75t_L g118 ( .A(n_34), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_35), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_36), .A2(n_155), .B(n_204), .C(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_L g546 ( .A(n_37), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_38), .A2(n_120), .B(n_123), .C(n_126), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_39), .A2(n_123), .B(n_486), .C(n_491), .Y(n_485) );
CKINVDCx14_ASAP7_75t_R g509 ( .A(n_40), .Y(n_509) );
INVx1_ASAP7_75t_L g211 ( .A(n_42), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_43), .A2(n_133), .B(n_201), .C(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_44), .B(n_156), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_45), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_46), .Y(n_542) );
INVx1_ASAP7_75t_L g476 ( .A(n_47), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_48), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_49), .B(n_115), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_50), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_51), .A2(n_123), .B1(n_189), .B2(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_52), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_53), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_54), .A2(n_201), .B(n_202), .C(n_204), .Y(n_200) );
CKINVDCx14_ASAP7_75t_R g445 ( .A(n_55), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_56), .Y(n_251) );
INVx1_ASAP7_75t_L g199 ( .A(n_57), .Y(n_199) );
INVx1_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_59), .Y(n_140) );
INVx1_ASAP7_75t_SL g512 ( .A(n_60), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_61), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_62), .B(n_196), .Y(n_480) );
INVx1_ASAP7_75t_L g501 ( .A(n_63), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_SL g221 ( .A1(n_64), .A2(n_131), .B(n_204), .C(n_222), .Y(n_221) );
INVxp67_ASAP7_75t_L g223 ( .A(n_65), .Y(n_223) );
INVx1_ASAP7_75t_L g719 ( .A(n_66), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_67), .A2(n_115), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_68), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_69), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_70), .A2(n_115), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g244 ( .A(n_71), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_72), .A2(n_166), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g455 ( .A(n_73), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_74), .Y(n_484) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_75), .A2(n_76), .B1(n_728), .B2(n_729), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_75), .Y(n_729) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_76), .A2(n_101), .B1(n_715), .B2(n_724), .C1(n_734), .C2(n_740), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_76), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_77), .A2(n_120), .B(n_123), .C(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_78), .A2(n_115), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g458 ( .A(n_79), .Y(n_458) );
AOI222xp33_ASAP7_75t_SL g102 ( .A1(n_80), .A2(n_103), .B1(n_106), .B2(n_706), .C1(n_707), .C2(n_711), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_81), .B(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx1_ASAP7_75t_L g467 ( .A(n_83), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_84), .B(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_85), .A2(n_120), .B(n_123), .C(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g432 ( .A(n_86), .Y(n_432) );
OR2x2_ASAP7_75t_L g705 ( .A(n_86), .B(n_433), .Y(n_705) );
OR2x2_ASAP7_75t_L g723 ( .A(n_86), .B(n_714), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_87), .A2(n_123), .B(n_500), .C(n_503), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_88), .B(n_149), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_89), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_90), .A2(n_120), .B(n_123), .C(n_152), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_91), .Y(n_161) );
INVx1_ASAP7_75t_L g220 ( .A(n_92), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g168 ( .A(n_93), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_94), .B(n_128), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_95), .B(n_145), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_96), .B(n_145), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_97), .A2(n_115), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g479 ( .A(n_98), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_99), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g706 ( .A(n_103), .Y(n_706) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_431), .B1(n_436), .B2(n_705), .Y(n_106) );
INVx2_ASAP7_75t_L g708 ( .A(n_107), .Y(n_708) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_400), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_293), .C(n_366), .Y(n_108) );
OAI211xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_178), .B(n_225), .C(n_277), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_146), .Y(n_111) );
AND2x2_ASAP7_75t_L g241 ( .A(n_112), .B(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g260 ( .A(n_112), .Y(n_260) );
INVx2_ASAP7_75t_L g275 ( .A(n_112), .Y(n_275) );
INVx1_ASAP7_75t_L g305 ( .A(n_112), .Y(n_305) );
AND2x2_ASAP7_75t_L g355 ( .A(n_112), .B(n_276), .Y(n_355) );
AOI32xp33_ASAP7_75t_L g382 ( .A1(n_112), .A2(n_310), .A3(n_383), .B1(n_385), .B2(n_386), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_112), .B(n_231), .Y(n_388) );
AND2x2_ASAP7_75t_L g415 ( .A(n_112), .B(n_258), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_112), .B(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_142), .Y(n_112) );
AOI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_122), .B(n_135), .Y(n_113) );
BUFx2_ASAP7_75t_L g166 ( .A(n_115), .Y(n_166) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_116), .B(n_120), .Y(n_183) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g490 ( .A(n_117), .Y(n_490) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g124 ( .A(n_118), .Y(n_124) );
INVx1_ASAP7_75t_L g190 ( .A(n_118), .Y(n_190) );
INVx1_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx3_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_119), .Y(n_131) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_119), .Y(n_172) );
INVx4_ASAP7_75t_SL g176 ( .A(n_120), .Y(n_176) );
BUFx3_ASAP7_75t_L g491 ( .A(n_120), .Y(n_491) );
INVx5_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
AND2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
BUFx3_ASAP7_75t_L g134 ( .A(n_124), .Y(n_134) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B(n_132), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_128), .A2(n_186), .B(n_187), .C(n_188), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_128), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_128), .A2(n_171), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_129), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_129), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_129), .B(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_132), .A2(n_247), .B(n_248), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_L g466 ( .A1(n_132), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_132), .A2(n_468), .B(n_501), .C(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g249 ( .A(n_135), .Y(n_249) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_136), .A2(n_181), .B(n_191), .Y(n_180) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_136), .A2(n_208), .B(n_215), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_136), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_138), .B(n_139), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
NOR2xp33_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx3_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_144), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_144), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_144), .A2(n_497), .B(n_504), .Y(n_496) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_145), .A2(n_218), .B(n_224), .Y(n_217) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_145), .Y(n_452) );
AND2x2_ASAP7_75t_L g304 ( .A(n_146), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g326 ( .A(n_146), .Y(n_326) );
AND2x2_ASAP7_75t_L g411 ( .A(n_146), .B(n_241), .Y(n_411) );
AND2x2_ASAP7_75t_L g414 ( .A(n_146), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_163), .Y(n_146) );
INVx2_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_147), .B(n_258), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_147), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g310 ( .A(n_147), .Y(n_310) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_160), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_148), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g549 ( .A(n_148), .Y(n_549) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_149), .A2(n_165), .B(n_177), .Y(n_164) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_149), .A2(n_443), .B(n_449), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_149), .A2(n_183), .B(n_484), .C(n_485), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_159), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_155), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_162), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_162), .B(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_162), .A2(n_463), .B(n_470), .Y(n_462) );
AND2x2_ASAP7_75t_L g252 ( .A(n_163), .B(n_233), .Y(n_252) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
AND2x2_ASAP7_75t_L g276 ( .A(n_164), .B(n_258), .Y(n_276) );
AND2x2_ASAP7_75t_L g345 ( .A(n_164), .B(n_242), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_176), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_169), .A2(n_176), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_169), .A2(n_176), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_SL g444 ( .A1(n_169), .A2(n_176), .B(n_445), .C(n_446), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_169), .A2(n_176), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_169), .A2(n_176), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_169), .A2(n_176), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g541 ( .A1(n_169), .A2(n_176), .B(n_542), .C(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_171), .B(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_171), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_171), .B(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g210 ( .A1(n_172), .A2(n_211), .B1(n_212), .B2(n_213), .Y(n_210) );
INVx2_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_176), .A2(n_183), .B1(n_209), .B2(n_214), .Y(n_208) );
INVx1_ASAP7_75t_L g503 ( .A(n_176), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_193), .Y(n_178) );
OR2x2_ASAP7_75t_L g239 ( .A(n_179), .B(n_207), .Y(n_239) );
INVx1_ASAP7_75t_L g318 ( .A(n_179), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_179), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_179), .B(n_206), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_179), .B(n_330), .Y(n_384) );
AND2x2_ASAP7_75t_L g392 ( .A(n_179), .B(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
AND2x2_ASAP7_75t_L g299 ( .A(n_180), .B(n_207), .Y(n_299) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_183), .A2(n_244), .B(n_245), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_183), .A2(n_464), .B(n_465), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_183), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_193), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g426 ( .A(n_193), .Y(n_426) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_206), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_194), .B(n_270), .Y(n_292) );
OR2x2_ASAP7_75t_L g321 ( .A(n_194), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g353 ( .A(n_194), .B(n_333), .Y(n_353) );
INVx1_ASAP7_75t_SL g373 ( .A(n_194), .Y(n_373) );
AND2x2_ASAP7_75t_L g377 ( .A(n_194), .B(n_238), .Y(n_377) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_195), .B(n_206), .Y(n_230) );
AND2x2_ASAP7_75t_L g237 ( .A(n_195), .B(n_217), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g280 ( .A(n_195), .B(n_262), .Y(n_280) );
INVx1_ASAP7_75t_SL g287 ( .A(n_195), .Y(n_287) );
BUFx2_ASAP7_75t_L g298 ( .A(n_195), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_195), .B(n_229), .Y(n_314) );
AND2x2_ASAP7_75t_L g329 ( .A(n_195), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g393 ( .A(n_195), .B(n_207), .Y(n_393) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_205), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_206), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g317 ( .A(n_206), .B(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_206), .A2(n_335), .B1(n_338), .B2(n_341), .C(n_346), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_206), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
INVx3_ASAP7_75t_L g262 ( .A(n_207), .Y(n_262) );
INVx2_ASAP7_75t_L g468 ( .A(n_212), .Y(n_468) );
BUFx2_ASAP7_75t_L g272 ( .A(n_217), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_217), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g303 ( .A(n_217), .Y(n_303) );
OR2x2_ASAP7_75t_L g322 ( .A(n_217), .B(n_262), .Y(n_322) );
INVx3_ASAP7_75t_L g330 ( .A(n_217), .Y(n_330) );
AND2x2_ASAP7_75t_L g333 ( .A(n_217), .B(n_262), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_231), .B1(n_235), .B2(n_240), .C(n_253), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_228), .B(n_302), .Y(n_427) );
OR2x2_ASAP7_75t_L g430 ( .A(n_228), .B(n_261), .Y(n_430) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OAI221xp5_ASAP7_75t_SL g253 ( .A1(n_229), .A2(n_254), .B1(n_261), .B2(n_263), .C(n_266), .Y(n_253) );
AND2x2_ASAP7_75t_L g270 ( .A(n_229), .B(n_262), .Y(n_270) );
AND2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_229), .B(n_286), .Y(n_285) );
NAND2x1_ASAP7_75t_L g328 ( .A(n_229), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g380 ( .A(n_229), .B(n_322), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_231), .A2(n_340), .B1(n_369), .B2(n_371), .Y(n_368) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AOI322xp5_ASAP7_75t_L g277 ( .A1(n_232), .A2(n_241), .A3(n_278), .B1(n_281), .B2(n_284), .C1(n_288), .C2(n_291), .Y(n_277) );
OR2x2_ASAP7_75t_L g289 ( .A(n_232), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_233), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g268 ( .A(n_233), .B(n_242), .Y(n_268) );
INVx1_ASAP7_75t_L g283 ( .A(n_233), .Y(n_283) );
AND2x2_ASAP7_75t_L g349 ( .A(n_233), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g259 ( .A(n_234), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g350 ( .A(n_234), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_234), .B(n_258), .Y(n_424) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_238), .B(n_373), .Y(n_372) );
INVx3_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g324 ( .A(n_239), .B(n_271), .Y(n_324) );
OR2x2_ASAP7_75t_L g421 ( .A(n_239), .B(n_272), .Y(n_421) );
INVx1_ASAP7_75t_L g402 ( .A(n_240), .Y(n_402) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_252), .Y(n_240) );
INVx4_ASAP7_75t_L g290 ( .A(n_241), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_241), .B(n_309), .Y(n_315) );
INVx2_ASAP7_75t_L g258 ( .A(n_242), .Y(n_258) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B(n_250), .Y(n_242) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_249), .A2(n_539), .B(n_547), .Y(n_538) );
INVx1_ASAP7_75t_L g556 ( .A(n_249), .Y(n_556) );
INVx1_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_252), .B(n_312), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g327 ( .A1(n_254), .A2(n_328), .B(n_331), .Y(n_327) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
INVx1_ASAP7_75t_L g339 ( .A(n_258), .Y(n_339) );
INVx1_ASAP7_75t_L g265 ( .A(n_259), .Y(n_265) );
AND2x2_ASAP7_75t_L g267 ( .A(n_259), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g363 ( .A(n_260), .B(n_349), .Y(n_363) );
AND2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_345), .Y(n_385) );
BUFx2_ASAP7_75t_L g337 ( .A(n_262), .Y(n_337) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AOI32xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .A3(n_270), .B1(n_271), .B2(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g347 ( .A(n_267), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_267), .A2(n_395), .B1(n_396), .B2(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_270), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_270), .B(n_329), .Y(n_370) );
AND2x2_ASAP7_75t_L g417 ( .A(n_270), .B(n_302), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_271), .B(n_318), .Y(n_365) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g418 ( .A(n_273), .Y(n_418) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g343 ( .A(n_274), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_276), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g390 ( .A(n_276), .B(n_310), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_276), .B(n_305), .Y(n_397) );
INVx1_ASAP7_75t_SL g379 ( .A(n_278), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_279), .B(n_330), .Y(n_357) );
NOR4xp25_ASAP7_75t_L g403 ( .A(n_279), .B(n_302), .C(n_404), .D(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_280), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g360 ( .A(n_283), .Y(n_360) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_286), .A2(n_377), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g302 ( .A(n_287), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND4xp25_ASAP7_75t_SL g293 ( .A(n_294), .B(n_319), .C(n_334), .D(n_354), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_300), .B(n_304), .C(n_306), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g386 ( .A(n_299), .B(n_329), .Y(n_386) );
AND2x2_ASAP7_75t_L g395 ( .A(n_299), .B(n_373), .Y(n_395) );
INVx3_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_302), .B(n_337), .Y(n_399) );
AND2x2_ASAP7_75t_L g311 ( .A(n_305), .B(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_315), .B2(n_316), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x2_ASAP7_75t_L g409 ( .A(n_309), .B(n_355), .Y(n_409) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_311), .B(n_360), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_312), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_325), .C(n_327), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_320), .A2(n_355), .B1(n_356), .B2(n_358), .C(n_361), .Y(n_354) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_328), .A2(n_413), .B1(n_416), .B2(n_418), .C(n_419), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_329), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_337), .B(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_342), .A2(n_362), .B1(n_364), .B2(n_365), .Y(n_361) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_351), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_362), .A2(n_388), .B1(n_426), .B2(n_427), .C(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_374), .C(n_394), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_378), .C(n_387), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_381), .C(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g406 ( .A(n_384), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g428 ( .A1(n_385), .A2(n_411), .B(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_391), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI21xp5_ASAP7_75t_SL g420 ( .A1(n_397), .A2(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .C(n_425), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_408), .C(n_410), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
CKINVDCx14_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g710 ( .A(n_431), .Y(n_710) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NOR2x2_ASAP7_75t_L g713 ( .A(n_432), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_433), .Y(n_714) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_SL g707 ( .A1(n_437), .A2(n_705), .B1(n_708), .B2(n_709), .Y(n_707) );
XOR2xp5_ASAP7_75t_L g726 ( .A(n_437), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_635), .Y(n_437) );
NAND5xp2_ASAP7_75t_L g438 ( .A(n_439), .B(n_550), .C(n_582), .D(n_599), .E(n_622), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_481), .B1(n_514), .B2(n_518), .C(n_522), .Y(n_439) );
INVx1_ASAP7_75t_L g662 ( .A(n_440), .Y(n_662) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_460), .Y(n_440) );
AND3x2_ASAP7_75t_L g637 ( .A(n_441), .B(n_462), .C(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_450), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_442), .B(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g529 ( .A(n_442), .Y(n_529) );
AND2x2_ASAP7_75t_L g533 ( .A(n_442), .B(n_472), .Y(n_533) );
INVx2_ASAP7_75t_L g559 ( .A(n_442), .Y(n_559) );
OR2x2_ASAP7_75t_L g570 ( .A(n_442), .B(n_473), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_442), .B(n_461), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_442), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g649 ( .A(n_442), .B(n_473), .Y(n_649) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
AND2x2_ASAP7_75t_L g590 ( .A(n_450), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_450), .B(n_461), .Y(n_609) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g521 ( .A(n_451), .B(n_461), .Y(n_521) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_451), .Y(n_528) );
AND2x2_ASAP7_75t_L g576 ( .A(n_451), .B(n_473), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_451), .B(n_460), .C(n_559), .Y(n_601) );
AND2x2_ASAP7_75t_L g666 ( .A(n_451), .B(n_462), .Y(n_666) );
AND2x2_ASAP7_75t_L g700 ( .A(n_451), .B(n_461), .Y(n_700) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_459), .Y(n_451) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_452), .A2(n_474), .B(n_480), .Y(n_473) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_452), .A2(n_507), .B(n_513), .Y(n_506) );
INVxp67_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_461), .B(n_559), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_461), .B(n_590), .Y(n_598) );
AND2x2_ASAP7_75t_L g648 ( .A(n_461), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g676 ( .A(n_461), .Y(n_676) );
INVx4_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g583 ( .A(n_462), .B(n_576), .Y(n_583) );
BUFx3_ASAP7_75t_L g615 ( .A(n_462), .Y(n_615) );
INVx2_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_473), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_481), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_494), .Y(n_481) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_515), .Y(n_514) );
INVx3_ASAP7_75t_SL g525 ( .A(n_482), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_482), .B(n_554), .Y(n_586) );
OR2x2_ASAP7_75t_L g605 ( .A(n_482), .B(n_495), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_482), .B(n_562), .Y(n_610) );
AND2x2_ASAP7_75t_L g613 ( .A(n_482), .B(n_555), .Y(n_613) );
AND2x2_ASAP7_75t_L g625 ( .A(n_482), .B(n_506), .Y(n_625) );
AND2x2_ASAP7_75t_L g641 ( .A(n_482), .B(n_496), .Y(n_641) );
AND2x4_ASAP7_75t_L g644 ( .A(n_482), .B(n_516), .Y(n_644) );
OR2x2_ASAP7_75t_L g661 ( .A(n_482), .B(n_597), .Y(n_661) );
OR2x2_ASAP7_75t_L g692 ( .A(n_482), .B(n_538), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_482), .B(n_620), .Y(n_694) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_490), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_536), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_494), .B(n_555), .Y(n_687) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
AND2x2_ASAP7_75t_L g524 ( .A(n_495), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g554 ( .A(n_495), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_538), .Y(n_562) );
AND2x2_ASAP7_75t_L g580 ( .A(n_495), .B(n_516), .Y(n_580) );
OR2x2_ASAP7_75t_L g597 ( .A(n_495), .B(n_555), .Y(n_597) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g517 ( .A(n_496), .Y(n_517) );
AND2x2_ASAP7_75t_L g620 ( .A(n_496), .B(n_506), .Y(n_620) );
INVx2_ASAP7_75t_L g516 ( .A(n_506), .Y(n_516) );
INVx1_ASAP7_75t_L g632 ( .A(n_506), .Y(n_632) );
AND2x2_ASAP7_75t_L g682 ( .A(n_506), .B(n_525), .Y(n_682) );
AND2x2_ASAP7_75t_L g535 ( .A(n_515), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_525), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_515), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_L g553 ( .A(n_516), .B(n_525), .Y(n_553) );
OR2x2_ASAP7_75t_L g669 ( .A(n_517), .B(n_643), .Y(n_669) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_520), .B(n_649), .Y(n_655) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
OAI32xp33_ASAP7_75t_L g611 ( .A1(n_521), .A2(n_612), .A3(n_614), .B1(n_616), .B2(n_617), .Y(n_611) );
OR2x2_ASAP7_75t_L g628 ( .A(n_521), .B(n_570), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g653 ( .A1(n_521), .A2(n_531), .B(n_558), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_526), .B1(n_531), .B2(n_534), .Y(n_522) );
INVxp33_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_524), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_525), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g579 ( .A(n_525), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g679 ( .A(n_525), .B(n_620), .Y(n_679) );
OR2x2_ASAP7_75t_L g703 ( .A(n_525), .B(n_597), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_526), .A2(n_585), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_530), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g563 ( .A(n_528), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_528), .B(n_533), .Y(n_581) );
AND2x2_ASAP7_75t_L g603 ( .A(n_529), .B(n_576), .Y(n_603) );
INVx1_ASAP7_75t_L g616 ( .A(n_529), .Y(n_616) );
OR2x2_ASAP7_75t_L g621 ( .A(n_529), .B(n_555), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_532), .B(n_570), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_533), .A2(n_552), .B1(n_557), .B2(n_561), .Y(n_551) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_536), .A2(n_594), .B1(n_601), .B2(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g678 ( .A(n_536), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_538), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g697 ( .A(n_538), .B(n_580), .Y(n_697) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_540), .A2(n_548), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_563), .B1(n_564), .B2(n_569), .C(n_571), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_553), .B(n_555), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_554), .A2(n_660), .B(n_661), .C(n_662), .Y(n_659) );
AND2x2_ASAP7_75t_L g664 ( .A(n_554), .B(n_644), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_SL g702 ( .A1(n_554), .A2(n_643), .B(n_703), .C(n_704), .Y(n_702) );
BUFx3_ASAP7_75t_L g594 ( .A(n_555), .Y(n_594) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_558), .B(n_615), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_558), .A2(n_678), .B(n_680), .C(n_686), .Y(n_677) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVxp67_ASAP7_75t_L g638 ( .A(n_560), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_562), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_566), .A2(n_583), .B(n_584), .C(n_592), .Y(n_582) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g667 ( .A(n_570), .Y(n_667) );
OR2x2_ASAP7_75t_L g684 ( .A(n_570), .B(n_614), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_578), .B2(n_581), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_573), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
OR2x2_ASAP7_75t_L g671 ( .A(n_575), .B(n_615), .Y(n_671) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g626 ( .A(n_576), .B(n_616), .Y(n_626) );
INVx1_ASAP7_75t_L g634 ( .A(n_577), .Y(n_634) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_580), .B(n_594), .Y(n_642) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_590), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g699 ( .A(n_591), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_598), .Y(n_592) );
INVx1_ASAP7_75t_L g629 ( .A(n_593), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_594), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_594), .B(n_625), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_594), .B(n_620), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_594), .B(n_641), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_594), .A2(n_604), .B(n_644), .C(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_604), .B1(n_606), .B2(n_610), .C(n_611), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_608), .B(n_616), .Y(n_690) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_610), .A2(n_625), .B(n_627), .C(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_613), .B(n_620), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_614), .B(n_667), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g614 ( .A(n_615), .Y(n_614) );
INVxp33_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AOI21xp33_ASAP7_75t_SL g630 ( .A1(n_619), .A2(n_631), .B(n_633), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_619), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_620), .B(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_627), .B2(n_629), .C(n_630), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_626), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g660 ( .A(n_632), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g635 ( .A(n_636), .B(n_663), .C(n_677), .D(n_688), .E(n_701), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_646), .C(n_659), .Y(n_636) );
INVx2_ASAP7_75t_SL g683 ( .A(n_637), .Y(n_683) );
NAND4xp25_ASAP7_75t_SL g639 ( .A(n_640), .B(n_642), .C(n_643), .D(n_645), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_645), .A2(n_647), .B(n_650), .C(n_656), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_648), .A2(n_689), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_672), .Y(n_663) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_671), .A2(n_694), .B1(n_696), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .Y(n_716) );
NOR2xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_SL g739 ( .A(n_718), .Y(n_739) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
OA21x2_ASAP7_75t_L g741 ( .A1(n_720), .A2(n_732), .B(n_739), .Y(n_741) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_723), .Y(n_730) );
BUFx2_ASAP7_75t_L g732 ( .A(n_723), .Y(n_732) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_730), .B(n_731), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
CKINVDCx6p67_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
endmodule