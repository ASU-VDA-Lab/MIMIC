module fake_jpeg_14609_n_368 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_368);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_368;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_38),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_48),
.B(n_62),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_94),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_19),
.B1(n_27),
.B2(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_68),
.A2(n_73),
.B1(n_75),
.B2(n_84),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_19),
.B1(n_22),
.B2(n_34),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_19),
.B1(n_22),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_29),
.B1(n_26),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_27),
.B1(n_16),
.B2(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_44),
.B1(n_64),
.B2(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_28),
.B1(n_35),
.B2(n_18),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_28),
.B1(n_35),
.B2(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_32),
.B1(n_24),
.B2(n_20),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_86),
.A2(n_88),
.B1(n_92),
.B2(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_87),
.B(n_111),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_24),
.B1(n_20),
.B2(n_16),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_29),
.B1(n_26),
.B2(n_4),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_91),
.A2(n_14),
.B1(n_28),
.B2(n_34),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_29),
.B(n_26),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_110),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_108),
.B1(n_99),
.B2(n_71),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_40),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_5),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_115),
.A2(n_129),
.B1(n_157),
.B2(n_121),
.Y(n_183)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_6),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_120),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_122),
.B1(n_132),
.B2(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_124),
.B(n_125),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_9),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_101),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_111),
.Y(n_128)
);

CKINVDCx11_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_9),
.B1(n_11),
.B2(n_73),
.Y(n_129)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_11),
.B1(n_103),
.B2(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_139),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_135),
.Y(n_181)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_66),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_137),
.B(n_149),
.Y(n_206)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_136),
.B1(n_128),
.B2(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_105),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_67),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_84),
.C(n_107),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_134),
.C(n_122),
.Y(n_187)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_96),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_71),
.B(n_85),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_159),
.CI(n_160),
.CON(n_184),
.SN(n_184)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_112),
.B(n_109),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_65),
.B(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_150),
.B1(n_130),
.B2(n_138),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_54),
.B1(n_46),
.B2(n_50),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_163),
.B1(n_159),
.B2(n_155),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_172),
.B(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_186),
.B1(n_195),
.B2(n_190),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_168),
.B(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_171),
.A2(n_182),
.B1(n_201),
.B2(n_168),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_143),
.B(n_132),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_149),
.B1(n_148),
.B2(n_123),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_175),
.A2(n_174),
.B1(n_181),
.B2(n_198),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_196),
.B(n_199),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_156),
.B1(n_147),
.B2(n_152),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_208),
.Y(n_223)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_194),
.Y(n_215)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_135),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_203),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_119),
.B(n_118),
.CI(n_134),
.CON(n_199),
.SN(n_199)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_199),
.B(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_137),
.A2(n_155),
.B1(n_152),
.B2(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_205),
.B1(n_208),
.B2(n_161),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_117),
.Y(n_202)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_127),
.A2(n_145),
.B1(n_146),
.B2(n_116),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_146),
.A2(n_141),
.B1(n_143),
.B2(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_218),
.B1(n_220),
.B2(n_230),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_186),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_212),
.A2(n_219),
.B(n_221),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_214),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_239),
.B(n_241),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_165),
.B1(n_186),
.B2(n_184),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_192),
.C(n_194),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_R g224 ( 
.A(n_199),
.B(n_190),
.C(n_206),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_232),
.B(n_243),
.Y(n_265)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_238),
.Y(n_260)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_184),
.B1(n_171),
.B2(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_173),
.B(n_170),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_174),
.B(n_176),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_235),
.B1(n_247),
.B2(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_237),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_196),
.B1(n_180),
.B2(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_179),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_177),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_176),
.A2(n_177),
.B(n_185),
.C(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_185),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_189),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_250),
.C(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_216),
.C(n_218),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_252),
.A2(n_264),
.B(n_274),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_224),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_262),
.C(n_268),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_217),
.C(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_237),
.C(n_212),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_242),
.B(n_243),
.CI(n_239),
.CON(n_271),
.SN(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_210),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_243),
.B(n_214),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_238),
.C(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_271),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_239),
.B(n_228),
.C(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_287),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_227),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_292),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_239),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_260),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_294),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_278),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_305),
.C(n_268),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_266),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_271),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_263),
.B(n_265),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_304),
.B(n_274),
.Y(n_311)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_267),
.B1(n_276),
.B2(n_272),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_248),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_254),
.B(n_272),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_251),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_253),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_262),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_311),
.A2(n_288),
.B(n_306),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_265),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_315),
.C(n_317),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_249),
.C(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_249),
.C(n_273),
.Y(n_317)
);

XNOR2x2_ASAP7_75t_SL g319 ( 
.A(n_293),
.B(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_280),
.A2(n_255),
.B1(n_276),
.B2(n_292),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_303),
.B1(n_284),
.B2(n_298),
.Y(n_338)
);

XOR2x2_ASAP7_75t_SL g326 ( 
.A(n_282),
.B(n_255),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_330),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_297),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_310),
.C(n_312),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_321),
.B(n_294),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_332),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_296),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_334),
.A2(n_337),
.B(n_288),
.Y(n_345)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_285),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_309),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_338),
.A2(n_340),
.B1(n_283),
.B2(n_287),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_286),
.B1(n_281),
.B2(n_303),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_329),
.A2(n_324),
.B1(n_319),
.B2(n_280),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_343),
.B1(n_351),
.B2(n_337),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_281),
.B1(n_284),
.B2(n_308),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_333),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_345),
.A2(n_334),
.B(n_330),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_307),
.C(n_317),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_333),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_338),
.B(n_299),
.CI(n_320),
.CON(n_347),
.SN(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_340),
.B(n_320),
.CI(n_323),
.CON(n_348),
.SN(n_348)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_350),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_356),
.C(n_357),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_356),
.B(n_346),
.C(n_335),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_344),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_353),
.A2(n_339),
.B1(n_336),
.B2(n_345),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_352),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.C(n_358),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_361),
.B1(n_341),
.B2(n_315),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_365),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_SL g367 ( 
.A1(n_366),
.A2(n_341),
.B1(n_327),
.B2(n_349),
.C(n_343),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_349),
.C(n_351),
.Y(n_368)
);


endmodule