module fake_jpeg_123_n_304 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_23),
.B1(n_41),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_81),
.B1(n_86),
.B2(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_88),
.B1(n_96),
.B2(n_105),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_40),
.B1(n_29),
.B2(n_35),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_97),
.B1(n_101),
.B2(n_1),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_29),
.C(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_40),
.B1(n_42),
.B2(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_90),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_36),
.B1(n_32),
.B2(n_24),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_26),
.B1(n_42),
.B2(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_36),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_32),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_40),
.B1(n_23),
.B2(n_31),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_109),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_107),
.B1(n_1),
.B2(n_5),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_15),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_112),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_99),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_137),
.Y(n_165)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_132),
.Y(n_154)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_97),
.B1(n_77),
.B2(n_111),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_94),
.B1(n_87),
.B2(n_84),
.Y(n_172)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_138),
.B1(n_146),
.B2(n_84),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_14),
.Y(n_132)
);

CKINVDCx10_ASAP7_75t_R g133 ( 
.A(n_83),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_133),
.Y(n_151)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_70),
.B(n_6),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_143),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

O2A1O1Ixp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_80),
.B(n_106),
.C(n_67),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_168),
.C(n_179),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_156),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_108),
.A3(n_107),
.B1(n_67),
.B2(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_98),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_79),
.Y(n_164)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_10),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_94),
.B(n_87),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_142),
.B(n_10),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_173),
.B1(n_13),
.B2(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_93),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_94),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_167),
.Y(n_193)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_140),
.C(n_127),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_146),
.B(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_200),
.B(n_202),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_123),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_185),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_141),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_93),
.B1(n_121),
.B2(n_128),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_202),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_131),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_165),
.B1(n_162),
.B2(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_171),
.B1(n_174),
.B2(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_126),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_151),
.A2(n_13),
.B(n_153),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_168),
.B(n_149),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_169),
.B1(n_160),
.B2(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_161),
.B1(n_174),
.B2(n_151),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_227),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_226),
.B(n_182),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_190),
.B(n_149),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_179),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_231),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_189),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_183),
.C(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_243),
.C(n_212),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_220),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_200),
.B(n_191),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_245),
.B(n_222),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_192),
.B1(n_195),
.B2(n_180),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_243),
.B1(n_230),
.B2(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_184),
.C(n_188),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_184),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_237),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_225),
.B1(n_230),
.B2(n_219),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_232),
.B1(n_240),
.B2(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_212),
.C(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_263),
.C(n_234),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_245),
.B(n_236),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_218),
.C(n_211),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_271),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_274),
.B1(n_252),
.B2(n_248),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_260),
.B(n_258),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_238),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_229),
.B(n_232),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_237),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_235),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_255),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_251),
.B1(n_256),
.B2(n_254),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_280),
.B(n_283),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_289),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_276),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_269),
.B(n_270),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_278),
.B1(n_281),
.B2(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_281),
.C(n_275),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_241),
.B1(n_275),
.B2(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_292),
.B1(n_257),
.B2(n_214),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_294),
.B(n_293),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_300),
.A3(n_297),
.B1(n_227),
.B2(n_228),
.C1(n_231),
.C2(n_214),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_218),
.B(n_244),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_302),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_213),
.Y(n_304)
);


endmodule