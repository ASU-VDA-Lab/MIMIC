module real_jpeg_25110_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_1),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_1),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_59),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_80),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_80),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_66),
.B1(n_69),
.B2(n_80),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_47),
.B1(n_54),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_5),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_88),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_88),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_66),
.B1(n_69),
.B2(n_88),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_148),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_7),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_177),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_177),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_7),
.A2(n_66),
.B1(n_69),
.B2(n_177),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_9),
.A2(n_49),
.B1(n_66),
.B2(n_69),
.Y(n_186)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_11),
.A2(n_45),
.B1(n_54),
.B2(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_11),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_120),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_120),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_11),
.A2(n_66),
.B1(n_69),
.B2(n_120),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_12),
.A2(n_48),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_12),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_146),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_146),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_12),
.A2(n_66),
.B1(n_69),
.B2(n_146),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_79),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_13),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_13),
.B(n_56),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_13),
.B(n_29),
.C(n_31),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_229),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_13),
.B(n_38),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_229),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_13),
.B(n_66),
.C(n_68),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_13),
.A2(n_101),
.B(n_289),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_15),
.A2(n_41),
.B1(n_66),
.B2(n_69),
.Y(n_108)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_16),
.B(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_95),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_22),
.B(n_81),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B1(n_60),
.B2(n_61),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_38),
.B(n_39),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_25),
.A2(n_38),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_25),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_25),
.A2(n_38),
.B1(n_196),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_26),
.A2(n_27),
.B1(n_92),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_26),
.A2(n_27),
.B1(n_124),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_26),
.A2(n_195),
.B(n_197),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_26),
.A2(n_197),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_27),
.A2(n_142),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_27),
.A2(n_181),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_28),
.A2(n_29),
.B1(n_67),
.B2(n_68),
.Y(n_71)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_29),
.B(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_35),
.B1(n_52),
.B2(n_53),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_34),
.A2(n_48),
.A3(n_53),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_35),
.B(n_52),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_35),
.B(n_255),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_38),
.B(n_182),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_55),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_48),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_50),
.A2(n_56),
.B1(n_145),
.B2(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_50),
.A2(n_150),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_77),
.B1(n_78),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_87),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_119),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_55),
.A2(n_117),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.C(n_76),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_86),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_63),
.A2(n_85),
.B1(n_90),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B(n_72),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_70),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_64),
.A2(n_70),
.B1(n_111),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_64),
.A2(n_70),
.B1(n_261),
.B2(n_263),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_64),
.B(n_226),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_65),
.A2(n_73),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_65),
.A2(n_126),
.B1(n_140),
.B2(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_65),
.A2(n_188),
.B(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_65),
.A2(n_225),
.B(n_262),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_65),
.B(n_229),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_69),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_70),
.B(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_144),
.B(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_82),
.A2(n_86),
.B1(n_160),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_86),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_86),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI31xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_161),
.A3(n_167),
.B(n_346),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_151),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_97),
.B(n_151),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_121),
.C(n_129),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_98),
.A2(n_121),
.B1(n_122),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_98),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_100),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_100),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_108),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_108),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_101),
.A2(n_134),
.B1(n_135),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_101),
.A2(n_205),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_101),
.B(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_101),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_107),
.B(n_229),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B(n_128),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_126),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_126),
.A2(n_277),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_129),
.A2(n_130),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.C(n_143),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_131),
.A2(n_132),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_141),
.B(n_143),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_162),
.A2(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_163),
.B(n_166),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_339),
.B(n_345),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_214),
.B(n_338),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_207),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_170),
.B(n_207),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_189),
.C(n_191),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_171),
.A2(n_172),
.B1(n_189),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_183),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_179),
.C(n_183),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_184),
.B(n_187),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_189),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_191),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_198),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_194),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_198),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_202),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_203),
.A2(n_300),
.B1(n_302),
.B2(n_304),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_209),
.B(n_210),
.C(n_213),
.Y(n_344)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_247),
.B(n_332),
.C(n_337),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_241),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_231),
.C(n_232),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_217),
.A2(n_218),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_223),
.C(n_227),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_231),
.B(n_232),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_326),
.B(n_331),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_278),
.B(n_325),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_267),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_267),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.C(n_264),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_256),
.Y(n_274)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_264),
.B1(n_265),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_274),
.C(n_275),
.Y(n_330)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_319),
.B(n_324),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_297),
.B(n_318),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_291),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_291),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_295),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_307),
.B(n_317),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_305),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_303),
.B(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_312),
.B(n_316),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_344),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_344),
.Y(n_345)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);


endmodule