module fake_jpeg_5526_n_80 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_15),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx11_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_0),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_20),
.B1(n_19),
.B2(n_21),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_17),
.B1(n_13),
.B2(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_34),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_27),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_36),
.C(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_52),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_31),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_13),
.B(n_1),
.C(n_2),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_66),
.B(n_67),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_42),
.C(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_38),
.C(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_43),
.B1(n_62),
.B2(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_62),
.B1(n_54),
.B2(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_1),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_74),
.B1(n_70),
.B2(n_4),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_4),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_72),
.B(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_7),
.Y(n_80)
);


endmodule