module fake_netlist_5_41_n_2201 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2201);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2201;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx5_ASAP7_75t_L g220 ( 
.A(n_76),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_91),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_167),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_125),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_25),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_112),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_130),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_6),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_78),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_48),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_71),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_47),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_98),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_154),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_7),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_101),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_135),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_121),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_145),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_70),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_139),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_102),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_194),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_126),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_26),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_73),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_88),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_86),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_161),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_214),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_146),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_59),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_179),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_142),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_23),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_51),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_94),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_17),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_97),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_32),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_21),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_123),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_69),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_176),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_150),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_15),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_47),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_188),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_92),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_96),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_192),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_175),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_42),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_113),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_32),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_166),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_84),
.Y(n_306)
);

BUFx2_ASAP7_75t_SL g307 ( 
.A(n_50),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_117),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_54),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_111),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_24),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_37),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_83),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_106),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_9),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_210),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_138),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_43),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_10),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_172),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_83),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_201),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_5),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_85),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_87),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_67),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_207),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_70),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_198),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_17),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_39),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_66),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_80),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_140),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_3),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_129),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_52),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_170),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_151),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_79),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_12),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_168),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_13),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_16),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_60),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_66),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_25),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_165),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_40),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_14),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_132),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_181),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_107),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_67),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_184),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_57),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_72),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_105),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_19),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_73),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_21),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_35),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_206),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_215),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_58),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_40),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_56),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_159),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_191),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_23),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_74),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_110),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_155),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_19),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_2),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_77),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_133),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_11),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_35),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_74),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_65),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_29),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_114),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_62),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_103),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_199),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_44),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_29),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_11),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_163),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_28),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_58),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_16),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_41),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_81),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_120),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_197),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_216),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_209),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_119),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_63),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_26),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_108),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_53),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_75),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_183),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_219),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_38),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_82),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_63),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_45),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_1),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_39),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_57),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_128),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_80),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_137),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_72),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_78),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_95),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_3),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_180),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_136),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_9),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_148),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_13),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_30),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_272),
.B(n_316),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_231),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_220),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_220),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_258),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_296),
.B(n_0),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_301),
.B(n_1),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_220),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_262),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_343),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_220),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_240),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_220),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_220),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_272),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_240),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_220),
.Y(n_449)
);

BUFx5_ASAP7_75t_L g450 ( 
.A(n_221),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_228),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_316),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_230),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_232),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_254),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_220),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_220),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_233),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_234),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_292),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_236),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_312),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_324),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_324),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_238),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_337),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_241),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_254),
.B(n_2),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_221),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_321),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_225),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_247),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_331),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_256),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_335),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_225),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_341),
.B(n_4),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_263),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_235),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_244),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_355),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_239),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_244),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_245),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_341),
.B(n_4),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_245),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_264),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_239),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_249),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_249),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_251),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_251),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_274),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_259),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_277),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_353),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_255),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_259),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_278),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_373),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_278),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_279),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_353),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_287),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_268),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_280),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_273),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_287),
.Y(n_514)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_417),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_289),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_403),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_411),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_289),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_295),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_281),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_285),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_295),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_307),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_293),
.B(n_5),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_288),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_268),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_290),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_304),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_298),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_298),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_300),
.Y(n_532)
);

INVxp33_ASAP7_75t_SL g533 ( 
.A(n_322),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_327),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_333),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_334),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_339),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_356),
.B(n_6),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_300),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_346),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_356),
.B(n_7),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_302),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_293),
.B(n_8),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_401),
.B(n_8),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_302),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_338),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_338),
.Y(n_547)
);

CKINVDCx14_ASAP7_75t_R g548 ( 
.A(n_271),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_337),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_360),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_404),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_348),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_434),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_511),
.B(n_404),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_461),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_441),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_466),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_435),
.A2(n_362),
.B(n_359),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_455),
.B(n_401),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_467),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_482),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_460),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_440),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_475),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_494),
.B(n_255),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_488),
.B(n_328),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_435),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_448),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_488),
.B(n_328),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_448),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_478),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_443),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_445),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_446),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_474),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_487),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_506),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_517),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_533),
.B(n_222),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_436),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_518),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_436),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_456),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_529),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_527),
.Y(n_599)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_551),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_451),
.B(n_453),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_456),
.A2(n_420),
.B(n_357),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_503),
.B(n_405),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_483),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_405),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_485),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_486),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_489),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_442),
.B(n_357),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_490),
.B(n_420),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_548),
.B(n_223),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_450),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_454),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_454),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_224),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_458),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_450),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_458),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_459),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_492),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_459),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_495),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_464),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_468),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_464),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_469),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_450),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_470),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_471),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_472),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_471),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_472),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_450),
.B(n_227),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_477),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_497),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_549),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_477),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_479),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_605),
.A2(n_433),
.B1(n_541),
.B2(n_538),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_586),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_589),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_573),
.B(n_608),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_605),
.A2(n_433),
.B1(n_544),
.B2(n_491),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_593),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_592),
.B(n_479),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_614),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_484),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_605),
.B(n_502),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_609),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_574),
.B(n_450),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_595),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_565),
.B(n_484),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_627),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_574),
.B(n_450),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_610),
.Y(n_669)
);

BUFx8_ASAP7_75t_SL g670 ( 
.A(n_553),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_611),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_624),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_574),
.B(n_450),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_612),
.B(n_473),
.C(n_493),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_575),
.B(n_498),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_616),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_SL g677 ( 
.A1(n_637),
.A2(n_253),
.B1(n_365),
.B2(n_294),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_596),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_598),
.A2(n_439),
.B1(n_452),
.B2(n_447),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_564),
.A2(n_502),
.B1(n_480),
.B2(n_465),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_575),
.B(n_578),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_500),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_578),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_578),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_607),
.B(n_493),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_577),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_583),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_576),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_623),
.B(n_499),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_602),
.B(n_499),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_555),
.A2(n_515),
.B1(n_501),
.B2(n_512),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_569),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_564),
.A2(n_509),
.B1(n_505),
.B2(n_507),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_576),
.B(n_359),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_616),
.B(n_501),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_641),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_569),
.B(n_508),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_626),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_569),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_640),
.B(n_504),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_613),
.B(n_510),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_613),
.B(n_514),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_617),
.B(n_508),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_577),
.B(n_512),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_516),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_571),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_642),
.B(n_519),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_582),
.B(n_522),
.C(n_521),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_571),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_617),
.B(n_521),
.Y(n_712)
);

INVx4_ASAP7_75t_SL g713 ( 
.A(n_600),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_593),
.B(n_520),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_628),
.B(n_523),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_584),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_593),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_584),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_603),
.B(n_530),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_593),
.B(n_273),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_604),
.B(n_522),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_585),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_606),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_619),
.B(n_526),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_635),
.B(n_374),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_558),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_619),
.B(n_526),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_593),
.B(n_273),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_564),
.A2(n_531),
.B1(n_539),
.B2(n_532),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_606),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_571),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_621),
.B(n_528),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_606),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_559),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_557),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_606),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_542),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_621),
.B(n_534),
.C(n_528),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_571),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_581),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_581),
.B(n_273),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_581),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_581),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_554),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_622),
.B(n_534),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_588),
.B(n_273),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_588),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_564),
.A2(n_546),
.B1(n_547),
.B2(n_545),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_556),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_622),
.B(n_271),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_556),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_588),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_568),
.A2(n_537),
.B1(n_552),
.B2(n_540),
.Y(n_757)
);

BUFx4f_ASAP7_75t_L g758 ( 
.A(n_588),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_604),
.B(n_537),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_588),
.B(n_540),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_560),
.Y(n_761)
);

INVx4_ASAP7_75t_SL g762 ( 
.A(n_559),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_603),
.A2(n_543),
.B1(n_525),
.B2(n_385),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_579),
.B(n_552),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_625),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_561),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_550),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_629),
.B(n_307),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_559),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_563),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_567),
.B(n_242),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_599),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_SL g773 ( 
.A(n_625),
.B(n_271),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_630),
.B(n_370),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_559),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_630),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_634),
.B(n_308),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_634),
.B(n_313),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_559),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_566),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_566),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_639),
.B(n_313),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_566),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_549),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_615),
.B(n_317),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_615),
.B(n_620),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_639),
.B(n_271),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_340),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_566),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_566),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_645),
.A2(n_438),
.B1(n_349),
.B2(n_358),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_646),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_631),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_644),
.A2(n_360),
.B1(n_385),
.B2(n_384),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_631),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_633),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_633),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_620),
.B(n_229),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_572),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_599),
.B(n_276),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_636),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_638),
.B(n_332),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_638),
.B(n_350),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_237),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_650),
.B(n_361),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_650),
.B(n_362),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_777),
.B(n_788),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_655),
.B(n_378),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_684),
.B(n_367),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_658),
.B(n_601),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_654),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_657),
.B(n_243),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_682),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_720),
.A2(n_366),
.B1(n_380),
.B2(n_330),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_767),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_684),
.B(n_367),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_695),
.B(n_273),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_652),
.A2(n_368),
.B1(n_377),
.B2(n_389),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_685),
.B(n_368),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_720),
.B(n_352),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_685),
.B(n_377),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_691),
.A2(n_299),
.B1(n_246),
.B2(n_428),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_702),
.B(n_785),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_681),
.B(n_647),
.C(n_674),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_654),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_656),
.B(n_572),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_804),
.B(n_389),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_694),
.A2(n_390),
.B1(n_391),
.B2(n_402),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_754),
.B(n_248),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_665),
.B(n_773),
.C(n_658),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_695),
.B(n_273),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_664),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_767),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_804),
.B(n_390),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_651),
.A2(n_513),
.B(n_402),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_784),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_782),
.B(n_379),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_L g841 ( 
.A1(n_689),
.A2(n_391),
.B(n_425),
.C(n_430),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_804),
.B(n_425),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_648),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_782),
.B(n_382),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_760),
.A2(n_323),
.B1(n_252),
.B2(n_257),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_774),
.B(n_601),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_656),
.B(n_250),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_649),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_720),
.A2(n_286),
.B1(n_310),
.B2(n_314),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_701),
.B(n_430),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_701),
.B(n_260),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_768),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_727),
.B(n_261),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_774),
.B(n_580),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_668),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_668),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_761),
.B(n_265),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_659),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_768),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_660),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_669),
.A2(n_297),
.B1(n_427),
.B2(n_266),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_671),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_692),
.B(n_267),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_799),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_679),
.B(n_383),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_675),
.A2(n_310),
.B(n_380),
.C(n_375),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_709),
.B(n_332),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_672),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_680),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_778),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_757),
.B(n_270),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_699),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_791),
.B(n_693),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_695),
.A2(n_730),
.B1(n_752),
.B2(n_763),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_741),
.B(n_386),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_716),
.B(n_388),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_683),
.A2(n_345),
.B1(n_275),
.B2(n_282),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_651),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_710),
.B(n_394),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_715),
.Y(n_881)
);

BUFx6f_ASAP7_75t_SL g882 ( 
.A(n_676),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_761),
.B(n_766),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_766),
.B(n_291),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_787),
.B(n_397),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_806),
.B(n_686),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_688),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_715),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_688),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_797),
.B(n_303),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_793),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_580),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_695),
.Y(n_894)
);

OAI221xp5_ASAP7_75t_L g895 ( 
.A1(n_794),
.A2(n_283),
.B1(n_226),
.B2(n_269),
.C(n_286),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_689),
.B(n_305),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_793),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_768),
.A2(n_387),
.B1(n_325),
.B2(n_326),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_770),
.B(n_306),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_768),
.A2(n_408),
.B1(n_309),
.B2(n_311),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_687),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_796),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_670),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_700),
.B(n_591),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_651),
.B(n_352),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_690),
.B(n_398),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_796),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_786),
.B(n_315),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_765),
.B(n_363),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_677),
.B(n_726),
.C(n_705),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_719),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_703),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_798),
.B(n_318),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_801),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_719),
.Y(n_915)
);

AND2x2_ASAP7_75t_SL g916 ( 
.A(n_687),
.B(n_352),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_698),
.B(n_399),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_407),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_764),
.B(n_410),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_801),
.B(n_347),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_709),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_722),
.Y(n_922)
);

CKINVDCx14_ASAP7_75t_R g923 ( 
.A(n_799),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_803),
.Y(n_924)
);

AO221x1_ASAP7_75t_L g925 ( 
.A1(n_718),
.A2(n_352),
.B1(n_354),
.B2(n_364),
.C(n_351),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_765),
.B(n_363),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_802),
.B(n_372),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_764),
.B(n_413),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_722),
.B(n_376),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_696),
.B(n_415),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_706),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_803),
.B(n_384),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_661),
.B(n_381),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_703),
.A2(n_226),
.B1(n_269),
.B2(n_330),
.Y(n_934)
);

INVxp33_ASAP7_75t_L g935 ( 
.A(n_772),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_661),
.B(n_395),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_740),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_661),
.B(n_412),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_800),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_803),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_759),
.B(n_422),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_709),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_759),
.B(n_276),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_663),
.B(n_352),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_734),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_L g946 ( 
.A(n_734),
.B(n_416),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_706),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_803),
.A2(n_418),
.B1(n_421),
.B2(n_423),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_704),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_663),
.A2(n_550),
.B(n_283),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_704),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_717),
.B(n_424),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_653),
.B(n_431),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_805),
.B(n_276),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_718),
.B(n_432),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_740),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_748),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_718),
.B(n_276),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_737),
.B(n_429),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_748),
.B(n_284),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_707),
.B(n_284),
.Y(n_961)
);

INVx8_ASAP7_75t_L g962 ( 
.A(n_670),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_712),
.B(n_429),
.Y(n_963)
);

AND2x4_ASAP7_75t_SL g964 ( 
.A(n_676),
.B(n_562),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_707),
.B(n_284),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_753),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_725),
.B(n_314),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_676),
.B(n_284),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_733),
.B(n_319),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_758),
.A2(n_375),
.B(n_320),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_879),
.A2(n_758),
.B(n_743),
.Y(n_971)
);

AO22x1_ASAP7_75t_L g972 ( 
.A1(n_809),
.A2(n_939),
.B1(n_910),
.B2(n_866),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_809),
.B(n_753),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_886),
.A2(n_749),
.B1(n_726),
.B2(n_744),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_879),
.A2(n_758),
.B(n_743),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_826),
.A2(n_667),
.B(n_673),
.C(n_662),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_921),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_832),
.B(n_570),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_820),
.A2(n_714),
.B(n_739),
.C(n_755),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_822),
.A2(n_746),
.B(n_742),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_875),
.A2(n_747),
.B(n_732),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_875),
.A2(n_747),
.B(n_732),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_868),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_815),
.B(n_678),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_822),
.A2(n_747),
.B(n_708),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_886),
.B(n_678),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_939),
.A2(n_751),
.B1(n_738),
.B2(n_731),
.Y(n_987)
);

OAI221xp5_ASAP7_75t_L g988 ( 
.A1(n_807),
.A2(n_319),
.B1(n_320),
.B2(n_329),
.C(n_342),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_944),
.A2(n_708),
.B(n_711),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_830),
.A2(n_808),
.B(n_807),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_919),
.B(n_776),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_921),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_908),
.A2(n_756),
.B(n_711),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_918),
.B(n_723),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_918),
.B(n_930),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_930),
.B(n_723),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_937),
.Y(n_998)
);

BUFx4f_ASAP7_75t_L g999 ( 
.A(n_962),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_956),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_933),
.A2(n_756),
.B(n_790),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_936),
.A2(n_790),
.B(n_769),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_905),
.A2(n_780),
.B(n_735),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_949),
.A2(n_721),
.B(n_729),
.C(n_745),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_921),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_921),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_829),
.A2(n_724),
.B(n_789),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_836),
.A2(n_842),
.B(n_816),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_957),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_816),
.B(n_789),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_912),
.B(n_587),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_938),
.A2(n_790),
.B(n_769),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_913),
.A2(n_769),
.B(n_734),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_868),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_883),
.B(n_736),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_922),
.B(n_591),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_817),
.B(n_736),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_901),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_916),
.B(n_776),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_892),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_813),
.A2(n_834),
.B(n_827),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_852),
.A2(n_734),
.B(n_775),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_897),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_945),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_835),
.B(n_736),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_838),
.B(n_781),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_945),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_945),
.A2(n_905),
.B(n_896),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_902),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_949),
.A2(n_783),
.B1(n_781),
.B2(n_729),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_840),
.B(n_781),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_966),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_855),
.B(n_666),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_951),
.A2(n_783),
.B1(n_721),
.B2(n_750),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_945),
.A2(n_779),
.B(n_713),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_850),
.A2(n_400),
.B1(n_342),
.B2(n_344),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_810),
.A2(n_942),
.B1(n_845),
.B2(n_839),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_847),
.B(n_594),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_935),
.B(n_594),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_947),
.B(n_839),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_953),
.A2(n_779),
.B(n_713),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_812),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_874),
.A2(n_888),
.B(n_881),
.C(n_811),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_871),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_919),
.B(n_697),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_928),
.B(n_792),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_853),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_955),
.A2(n_779),
.B(n_713),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_845),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_850),
.A2(n_934),
.B1(n_916),
.B2(n_967),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_920),
.A2(n_779),
.B(n_713),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_889),
.B(n_783),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_907),
.A2(n_762),
.B(n_779),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_853),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_928),
.B(n_590),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_967),
.A2(n_969),
.B1(n_810),
.B2(n_866),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_906),
.B(n_776),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_927),
.A2(n_762),
.B(n_419),
.Y(n_1058)
);

OR2x2_ASAP7_75t_SL g1059 ( 
.A(n_924),
.B(n_329),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_818),
.A2(n_762),
.B(n_419),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_963),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_844),
.B(n_762),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_959),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_914),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_821),
.A2(n_344),
.B(n_414),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_823),
.A2(n_351),
.B(n_414),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_849),
.B(n_354),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_841),
.A2(n_392),
.B(n_409),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_L g1069 ( 
.A(n_906),
.B(n_426),
.C(n_409),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_891),
.A2(n_406),
.B(n_400),
.Y(n_1070)
);

OAI321xp33_ASAP7_75t_L g1071 ( 
.A1(n_969),
.A2(n_406),
.A3(n_393),
.B1(n_392),
.B2(n_371),
.C(n_369),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_885),
.B(n_393),
.C(n_371),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_876),
.A2(n_336),
.B1(n_366),
.B2(n_364),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_859),
.B(n_369),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_925),
.A2(n_336),
.B1(n_12),
.B2(n_14),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_934),
.A2(n_10),
.B1(n_18),
.B2(n_20),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_876),
.B(n_336),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_870),
.B(n_89),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_854),
.A2(n_157),
.B(n_213),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_893),
.B(n_336),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_885),
.A2(n_18),
.B(n_20),
.C(n_22),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_882),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_L g1083 ( 
.A(n_894),
.B(n_212),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_858),
.A2(n_884),
.B(n_899),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_954),
.A2(n_208),
.B(n_205),
.C(n_204),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_917),
.A2(n_22),
.B(n_24),
.C(n_27),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_851),
.A2(n_203),
.B(n_195),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_843),
.A2(n_190),
.B(n_189),
.Y(n_1088)
);

AO22x1_ASAP7_75t_L g1089 ( 
.A1(n_917),
.A2(n_880),
.B1(n_860),
.B2(n_963),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_856),
.A2(n_857),
.B(n_958),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_887),
.A2(n_186),
.B(n_174),
.Y(n_1091)
);

INVx3_ASAP7_75t_SL g1092 ( 
.A(n_962),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_814),
.A2(n_173),
.B(n_160),
.C(n_158),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_890),
.A2(n_153),
.B(n_152),
.Y(n_1094)
);

BUFx8_ASAP7_75t_L g1095 ( 
.A(n_882),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_904),
.B(n_147),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_911),
.A2(n_141),
.B(n_134),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_915),
.B(n_131),
.Y(n_1098)
);

AO22x1_ASAP7_75t_L g1099 ( 
.A1(n_880),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_895),
.A2(n_31),
.B(n_34),
.C(n_36),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_828),
.B(n_34),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_961),
.A2(n_127),
.B(n_124),
.C(n_122),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_861),
.A2(n_116),
.B(n_115),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_863),
.A2(n_109),
.B(n_100),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_869),
.A2(n_93),
.B(n_90),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_873),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_837),
.A2(n_36),
.B(n_37),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_952),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_968),
.B(n_38),
.C(n_41),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_970),
.B(n_42),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_860),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_943),
.B(n_848),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_909),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_931),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_867),
.A2(n_46),
.B(n_49),
.C(n_51),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_960),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_819),
.A2(n_49),
.B(n_52),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_833),
.A2(n_53),
.B(n_55),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_L g1119 ( 
.A(n_831),
.B(n_55),
.Y(n_1119)
);

NOR3xp33_ASAP7_75t_L g1120 ( 
.A(n_872),
.B(n_56),
.C(n_59),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_877),
.B(n_61),
.Y(n_1121)
);

AOI22x1_ASAP7_75t_L g1122 ( 
.A1(n_924),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_877),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_864),
.A2(n_64),
.B(n_65),
.C(n_68),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_900),
.B(n_68),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_965),
.A2(n_71),
.B(n_75),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_940),
.B(n_76),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_946),
.A2(n_950),
.B(n_929),
.Y(n_1128)
);

BUFx4f_ASAP7_75t_L g1129 ( 
.A(n_962),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_909),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_824),
.B(n_77),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_941),
.A2(n_81),
.B(n_82),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_909),
.B(n_926),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_926),
.B(n_959),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_846),
.A2(n_940),
.B(n_878),
.C(n_862),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_926),
.A2(n_932),
.B1(n_959),
.B2(n_923),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_894),
.A2(n_932),
.B(n_898),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_932),
.Y(n_1138)
);

AO32x1_ASAP7_75t_L g1139 ( 
.A1(n_948),
.A2(n_964),
.A3(n_894),
.B1(n_931),
.B2(n_903),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_894),
.A2(n_826),
.B(n_875),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_894),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_912),
.B(n_951),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_809),
.B(n_825),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_879),
.A2(n_661),
.B(n_651),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_809),
.B(n_825),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_816),
.A2(n_850),
.B1(n_875),
.B2(n_809),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_820),
.A2(n_809),
.B(n_830),
.C(n_808),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_816),
.A2(n_850),
.B1(n_875),
.B2(n_809),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_816),
.A2(n_850),
.B1(n_875),
.B2(n_809),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_892),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_809),
.B(n_825),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_816),
.A2(n_850),
.B1(n_875),
.B2(n_809),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1146),
.A2(n_1148),
.A3(n_1149),
.B(n_1152),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_992),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_992),
.B(n_1005),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_980),
.A2(n_1088),
.B(n_1003),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1020),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1023),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1151),
.B(n_1033),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1029),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_996),
.B(n_973),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1123),
.B(n_1049),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1146),
.A2(n_1152),
.B(n_1149),
.C(n_1148),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1092),
.Y(n_1166)
);

INVx3_ASAP7_75t_SL g1167 ( 
.A(n_1114),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1028),
.A2(n_989),
.B(n_982),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_L g1169 ( 
.A1(n_981),
.A2(n_986),
.B(n_1001),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1064),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1040),
.B(n_991),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1090),
.A2(n_1013),
.B(n_1012),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1002),
.A2(n_975),
.B(n_971),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1077),
.A2(n_1056),
.B(n_1057),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_972),
.B(n_1061),
.Y(n_1175)
);

NAND2x1_ASAP7_75t_L g1176 ( 
.A(n_1005),
.B(n_1006),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1150),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1005),
.B(n_1006),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_990),
.A2(n_1121),
.B(n_1008),
.C(n_997),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_990),
.A2(n_1008),
.B(n_1140),
.C(n_1007),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_994),
.A2(n_985),
.B(n_1048),
.Y(n_1181)
);

INVxp67_ASAP7_75t_SL g1182 ( 
.A(n_1024),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1084),
.A2(n_1015),
.B(n_1007),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1017),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_984),
.A2(n_995),
.B(n_976),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1025),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1140),
.A2(n_1147),
.B(n_1037),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_984),
.A2(n_1128),
.B(n_1137),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1016),
.B(n_1082),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1010),
.A2(n_979),
.B(n_1043),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1050),
.B(n_1006),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1018),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1041),
.A2(n_1051),
.B(n_1035),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1078),
.A2(n_1098),
.B(n_1141),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_1110),
.A2(n_1131),
.B(n_1078),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_L g1196 ( 
.A(n_1050),
.B(n_1024),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1106),
.B(n_1142),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1011),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1044),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1026),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1116),
.B(n_1108),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1010),
.A2(n_1004),
.B(n_1031),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1044),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1086),
.A2(n_1081),
.A3(n_1110),
.B(n_1076),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1024),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_1132),
.A2(n_1126),
.B(n_1117),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1083),
.A2(n_1135),
.B(n_1034),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_974),
.A2(n_1106),
.B1(n_1030),
.B2(n_1045),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1089),
.B(n_1142),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1046),
.A2(n_1112),
.B1(n_977),
.B2(n_1019),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_977),
.B(n_1098),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1101),
.A2(n_1069),
.B(n_988),
.C(n_1071),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1076),
.A2(n_1118),
.A3(n_1036),
.B(n_1111),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1062),
.A2(n_1052),
.B(n_1096),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1055),
.B(n_1038),
.Y(n_1215)
);

NOR2x1_ASAP7_75t_L g1216 ( 
.A(n_1082),
.B(n_978),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_983),
.B(n_1014),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1058),
.A2(n_1027),
.B(n_1060),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_998),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1011),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1027),
.A2(n_1000),
.B(n_1009),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1042),
.B(n_1080),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1032),
.A2(n_1079),
.B(n_1125),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1039),
.B(n_1047),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_987),
.A2(n_1093),
.B(n_1087),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1044),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1054),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1107),
.A2(n_1102),
.B(n_1085),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1074),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1104),
.B(n_1105),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1068),
.A2(n_1070),
.B(n_1075),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1067),
.B(n_1113),
.Y(n_1232)
);

AOI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_1133),
.A2(n_1073),
.B(n_1134),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1091),
.A2(n_1094),
.B(n_1097),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_SL g1236 ( 
.A(n_1095),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1124),
.A2(n_1071),
.B(n_1119),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1127),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_999),
.B(n_1129),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1036),
.A2(n_1111),
.A3(n_1065),
.B(n_1066),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1130),
.A2(n_1068),
.B(n_1100),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1120),
.A2(n_1138),
.B(n_1115),
.Y(n_1242)
);

BUFx8_ASAP7_75t_SL g1243 ( 
.A(n_999),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1127),
.B(n_1136),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1063),
.B(n_1136),
.Y(n_1245)
);

AOI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1122),
.A2(n_1129),
.B(n_993),
.Y(n_1246)
);

NAND2x1_ASAP7_75t_L g1247 ( 
.A(n_1114),
.B(n_1139),
.Y(n_1247)
);

BUFx8_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1059),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1099),
.B(n_1095),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1139),
.A2(n_661),
.B(n_651),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1139),
.B(n_809),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1146),
.A2(n_1149),
.B(n_1152),
.C(n_1148),
.Y(n_1253)
);

AOI221x1_ASAP7_75t_L g1254 ( 
.A1(n_1077),
.A2(n_996),
.B1(n_990),
.B2(n_1121),
.C(n_1050),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1092),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1022),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_992),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1020),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1146),
.A2(n_820),
.A3(n_1149),
.B(n_1148),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1024),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1022),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1106),
.B(n_1142),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1095),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1056),
.A2(n_996),
.B1(n_1145),
.B2(n_1143),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1020),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_996),
.A2(n_990),
.B(n_1140),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1106),
.B(n_1142),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1056),
.A2(n_809),
.B(n_996),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1021),
.A2(n_980),
.B(n_1088),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1021),
.A2(n_980),
.B(n_1088),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1021),
.A2(n_980),
.B(n_1088),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1021),
.Y(n_1280)
);

AO21x1_ASAP7_75t_L g1281 ( 
.A1(n_996),
.A2(n_990),
.B(n_1077),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1007),
.A2(n_1140),
.B(n_1008),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1021),
.A2(n_980),
.B(n_1088),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1018),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1146),
.A2(n_1149),
.B(n_1152),
.C(n_1148),
.Y(n_1286)
);

BUFx4_ASAP7_75t_SL g1287 ( 
.A(n_993),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1022),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1020),
.Y(n_1290)
);

O2A1O1Ixp5_ASAP7_75t_L g1291 ( 
.A1(n_996),
.A2(n_990),
.B(n_1077),
.C(n_1121),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1146),
.A2(n_1149),
.B(n_1152),
.C(n_1148),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_996),
.A2(n_990),
.B(n_1140),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1022),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1144),
.A2(n_661),
.B(n_651),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1020),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1024),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1022),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1020),
.Y(n_1301)
);

AO21x1_ASAP7_75t_L g1302 ( 
.A1(n_996),
.A2(n_990),
.B(n_1077),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1021),
.A2(n_980),
.B(n_1088),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1092),
.Y(n_1305)
);

INVx3_ASAP7_75t_SL g1306 ( 
.A(n_1166),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1158),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1199),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1171),
.B(n_1285),
.Y(n_1309)
);

OAI321xp33_ASAP7_75t_L g1310 ( 
.A1(n_1268),
.A2(n_1272),
.A3(n_1294),
.B1(n_1187),
.B2(n_1212),
.C(n_1237),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1248),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1304),
.B(n_1161),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1155),
.B(n_1260),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1174),
.A2(n_1274),
.B(n_1212),
.C(n_1291),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1248),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1265),
.B(n_1270),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1255),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1192),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1248),
.Y(n_1319)
);

O2A1O1Ixp5_ASAP7_75t_L g1320 ( 
.A1(n_1291),
.A2(n_1302),
.B(n_1281),
.C(n_1179),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1199),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1160),
.Y(n_1323)
);

INVx5_ASAP7_75t_L g1324 ( 
.A(n_1243),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1284),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1203),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1162),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1197),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1287),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1166),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1271),
.B(n_1293),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1215),
.B(n_1295),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1167),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1243),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1163),
.B(n_1229),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1201),
.B(n_1198),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1207),
.A2(n_1183),
.B(n_1185),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1250),
.A2(n_1222),
.B1(n_1220),
.B2(n_1175),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1249),
.A2(n_1175),
.B1(n_1244),
.B2(n_1252),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1252),
.A2(n_1233),
.B1(n_1209),
.B2(n_1242),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1287),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1257),
.B(n_1176),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1164),
.B(n_1192),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1267),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1170),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1179),
.A2(n_1180),
.B(n_1253),
.C(n_1165),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1165),
.A2(n_1253),
.B1(n_1292),
.B2(n_1286),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1232),
.B(n_1224),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1235),
.B(n_1210),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1254),
.B(n_1286),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1255),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1305),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1263),
.B(n_1273),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_1273),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1167),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1292),
.B(n_1184),
.Y(n_1357)
);

AND2x2_ASAP7_75t_SL g1358 ( 
.A(n_1196),
.B(n_1231),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1245),
.B(n_1227),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1230),
.A2(n_1225),
.B(n_1190),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1203),
.B(n_1226),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1226),
.B(n_1217),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1177),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1217),
.B(n_1216),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1258),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1217),
.Y(n_1366)
);

INVx6_ASAP7_75t_SL g1367 ( 
.A(n_1236),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1189),
.B(n_1305),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1269),
.B(n_1290),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1186),
.B(n_1200),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1298),
.B(n_1301),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1251),
.A2(n_1169),
.B(n_1168),
.Y(n_1372)
);

NOR3xp33_ASAP7_75t_L g1373 ( 
.A(n_1246),
.B(n_1208),
.C(n_1180),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1191),
.A2(n_1231),
.B1(n_1282),
.B2(n_1241),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1196),
.A2(n_1191),
.B(n_1206),
.C(n_1247),
.Y(n_1375)
);

CKINVDCx16_ASAP7_75t_R g1376 ( 
.A(n_1267),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1219),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1154),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1223),
.A2(n_1172),
.B(n_1214),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1153),
.B(n_1259),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1231),
.A2(n_1282),
.B1(n_1202),
.B2(n_1182),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1259),
.B(n_1153),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1156),
.Y(n_1383)
);

OR2x6_ASAP7_75t_SL g1384 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1211),
.A2(n_1239),
.B(n_1221),
.C(n_1154),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1282),
.B(n_1280),
.C(n_1257),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1159),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1159),
.B(n_1205),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1259),
.B(n_1153),
.Y(n_1389)
);

INVx3_ASAP7_75t_SL g1390 ( 
.A(n_1261),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1264),
.A2(n_1289),
.B(n_1279),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1261),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1261),
.B(n_1299),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1156),
.B(n_1178),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1205),
.B(n_1182),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1153),
.B(n_1259),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1261),
.B(n_1299),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1299),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1204),
.B(n_1240),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1299),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1213),
.A2(n_1178),
.B1(n_1234),
.B2(n_1204),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1240),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1204),
.B(n_1240),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1204),
.B(n_1240),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1213),
.B(n_1194),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1218),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1193),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1228),
.A2(n_1168),
.B(n_1181),
.C(n_1173),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1157),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_1275),
.B(n_1297),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1157),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1276),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1276),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1256),
.B(n_1300),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1277),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1277),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1262),
.B(n_1296),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1195),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1288),
.B(n_1278),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1278),
.B(n_1303),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1283),
.B(n_1303),
.Y(n_1421)
);

O2A1O1Ixp5_ASAP7_75t_L g1422 ( 
.A1(n_1195),
.A2(n_996),
.B(n_1174),
.C(n_1077),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1283),
.A2(n_1146),
.B1(n_1149),
.B2(n_1148),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1161),
.B(n_1155),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1188),
.A2(n_1185),
.B(n_1207),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1171),
.B(n_1285),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1199),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1199),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1215),
.A2(n_809),
.B1(n_996),
.B2(n_1077),
.Y(n_1431)
);

AND2x2_ASAP7_75t_SL g1432 ( 
.A(n_1215),
.B(n_1077),
.Y(n_1432)
);

OAI21xp33_ASAP7_75t_L g1433 ( 
.A1(n_1274),
.A2(n_809),
.B(n_1056),
.Y(n_1433)
);

AOI221x1_ASAP7_75t_L g1434 ( 
.A1(n_1174),
.A2(n_1252),
.B1(n_1077),
.B2(n_996),
.C(n_1165),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1243),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1158),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1199),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_1166),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1171),
.B(n_1285),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1188),
.A2(n_1207),
.B(n_1183),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1192),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1248),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1174),
.A2(n_996),
.B(n_809),
.C(n_1056),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1171),
.B(n_1285),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1155),
.A2(n_1146),
.B1(n_1149),
.B2(n_1148),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1284),
.B(n_832),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1188),
.A2(n_1207),
.B(n_1183),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1215),
.A2(n_809),
.B1(n_773),
.B2(n_754),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1155),
.A2(n_1146),
.B1(n_1149),
.B2(n_1148),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1192),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1174),
.A2(n_809),
.B1(n_996),
.B2(n_1077),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1284),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1284),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1192),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1284),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1171),
.B(n_1285),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1161),
.B(n_1155),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_1166),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1291),
.A2(n_1180),
.B(n_1272),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1207),
.A2(n_1148),
.B(n_1146),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1155),
.A2(n_1146),
.B1(n_1149),
.B2(n_1148),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1376),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1398),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1358),
.B(n_1411),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_SL g1472 ( 
.A(n_1438),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1396),
.B(n_1309),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1457),
.A2(n_1433),
.B1(n_1432),
.B2(n_1454),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1359),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1363),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1307),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1398),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1323),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1327),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1318),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1346),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1365),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1444),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1334),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1431),
.A2(n_1348),
.B1(n_1350),
.B2(n_1468),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1426),
.B(n_1439),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1313),
.A2(n_1331),
.B1(n_1316),
.B2(n_1333),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1418),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1463),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1313),
.B(n_1331),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1348),
.A2(n_1468),
.B1(n_1449),
.B2(n_1455),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1398),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1449),
.A2(n_1455),
.B1(n_1423),
.B2(n_1312),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1328),
.B(n_1322),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1436),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1377),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1410),
.A2(n_1391),
.B(n_1379),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1456),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1446),
.A2(n_1429),
.B1(n_1443),
.B2(n_1450),
.Y(n_1501)
);

AOI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1314),
.A2(n_1422),
.B(n_1310),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1402),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1409),
.B(n_1415),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1341),
.A2(n_1339),
.B1(n_1340),
.B2(n_1373),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1399),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1418),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1403),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1412),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1370),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1428),
.B(n_1441),
.Y(n_1511)
);

BUFx2_ASAP7_75t_R g1512 ( 
.A(n_1329),
.Y(n_1512)
);

BUFx2_ASAP7_75t_R g1513 ( 
.A(n_1342),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1452),
.A2(n_1423),
.B1(n_1349),
.B2(n_1351),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_SL g1515 ( 
.A(n_1438),
.Y(n_1515)
);

BUFx2_ASAP7_75t_R g1516 ( 
.A(n_1384),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1404),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1405),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_SL g1519 ( 
.A(n_1465),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1434),
.A2(n_1360),
.B(n_1310),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1356),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1311),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1441),
.A2(n_1450),
.B1(n_1443),
.B2(n_1459),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1308),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1369),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1409),
.B(n_1415),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1351),
.A2(n_1357),
.B1(n_1440),
.B2(n_1448),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1367),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1390),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1418),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1408),
.A2(n_1442),
.B(n_1453),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1369),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1357),
.A2(n_1332),
.B1(n_1322),
.B2(n_1451),
.Y(n_1533)
);

BUFx4f_ASAP7_75t_SL g1534 ( 
.A(n_1367),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1461),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1344),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1328),
.B(n_1332),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_SL g1538 ( 
.A(n_1315),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1371),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1406),
.B(n_1419),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1440),
.Y(n_1541)
);

AO21x1_ASAP7_75t_SL g1542 ( 
.A1(n_1382),
.A2(n_1389),
.B(n_1466),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1317),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1319),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1406),
.B(n_1421),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1467),
.B(n_1375),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1459),
.A2(n_1336),
.B1(n_1464),
.B2(n_1424),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1366),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1336),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1372),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1448),
.A2(n_1451),
.B1(n_1354),
.B2(n_1355),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1308),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1394),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1337),
.A2(n_1462),
.B1(n_1325),
.B2(n_1460),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1389),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1354),
.B(n_1355),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1458),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1387),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1383),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1392),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1394),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1445),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1362),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1324),
.A2(n_1435),
.B1(n_1335),
.B2(n_1306),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1321),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1364),
.A2(n_1368),
.B1(n_1401),
.B2(n_1326),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1413),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1416),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1393),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1414),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1352),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1361),
.B(n_1395),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1321),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1414),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1324),
.A2(n_1435),
.B1(n_1335),
.B2(n_1374),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1394),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1380),
.A2(n_1374),
.B1(n_1466),
.B2(n_1435),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1397),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1324),
.A2(n_1335),
.B1(n_1368),
.B2(n_1338),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1388),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1345),
.Y(n_1582)
);

BUFx10_ASAP7_75t_L g1583 ( 
.A(n_1361),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1330),
.A2(n_1353),
.B1(n_1465),
.B2(n_1338),
.Y(n_1584)
);

INVx5_ASAP7_75t_L g1585 ( 
.A(n_1417),
.Y(n_1585)
);

BUFx4f_ASAP7_75t_SL g1586 ( 
.A(n_1430),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1430),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1388),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1427),
.A2(n_1347),
.B1(n_1378),
.B2(n_1343),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1430),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1381),
.A2(n_1437),
.B1(n_1386),
.B2(n_1343),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1437),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1437),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1386),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1400),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1417),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1417),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1385),
.B(n_1420),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1457),
.A2(n_1174),
.B1(n_809),
.B2(n_1077),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1363),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1380),
.B(n_1382),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1396),
.B(n_1309),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1359),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1396),
.B(n_1309),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1359),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1363),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1457),
.A2(n_1174),
.B1(n_809),
.B2(n_1077),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1432),
.A2(n_809),
.B1(n_1055),
.B2(n_1215),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_SL g1609 ( 
.A(n_1431),
.B(n_809),
.C(n_1056),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1418),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1432),
.A2(n_1077),
.B1(n_809),
.B2(n_1057),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1363),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1334),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1318),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1359),
.Y(n_1615)
);

AO21x1_ASAP7_75t_SL g1616 ( 
.A1(n_1351),
.A2(n_1405),
.B(n_1174),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1457),
.A2(n_809),
.B(n_996),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1457),
.A2(n_1174),
.B1(n_809),
.B2(n_1077),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1431),
.A2(n_1056),
.B1(n_809),
.B2(n_1457),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1363),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1320),
.A2(n_1360),
.B(n_1425),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1432),
.A2(n_1077),
.B1(n_809),
.B2(n_1057),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1431),
.A2(n_1056),
.B1(n_809),
.B2(n_1457),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1520),
.A2(n_1502),
.B(n_1499),
.Y(n_1624)
);

INVx6_ASAP7_75t_L g1625 ( 
.A(n_1583),
.Y(n_1625)
);

BUFx2_ASAP7_75t_SL g1626 ( 
.A(n_1472),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1577),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1473),
.B(n_1602),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1509),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1473),
.B(n_1602),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1577),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1582),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1481),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1475),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1503),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1604),
.B(n_1506),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1510),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1611),
.B(n_1622),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1518),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1604),
.B(n_1506),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1475),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1609),
.A2(n_1623),
.B1(n_1619),
.B2(n_1618),
.Y(n_1642)
);

OR2x6_ASAP7_75t_L g1643 ( 
.A(n_1546),
.B(n_1471),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1599),
.A2(n_1607),
.B(n_1617),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

AND2x4_ASAP7_75t_SL g1647 ( 
.A(n_1553),
.B(n_1561),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1487),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1508),
.B(n_1517),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1492),
.B(n_1488),
.Y(n_1650)
);

BUFx4f_ASAP7_75t_SL g1651 ( 
.A(n_1562),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1503),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1597),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1550),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1542),
.B(n_1555),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1511),
.B(n_1547),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1567),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1585),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1567),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1569),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1569),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1542),
.B(n_1616),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1549),
.B(n_1536),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1605),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1571),
.B(n_1575),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1571),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1504),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1601),
.B(n_1495),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_SL g1670 ( 
.A(n_1478),
.B(n_1494),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1546),
.B(n_1471),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1575),
.B(n_1596),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1521),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1596),
.B(n_1489),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1598),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1594),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1504),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1605),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1526),
.Y(n_1679)
);

INVxp33_ASAP7_75t_L g1680 ( 
.A(n_1487),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1486),
.A2(n_1474),
.B1(n_1505),
.B2(n_1493),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1526),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1615),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1615),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1489),
.B(n_1507),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1471),
.B(n_1578),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1489),
.B(n_1507),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1585),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1585),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1585),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1585),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1545),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1545),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1540),
.A2(n_1490),
.B(n_1621),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1477),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1597),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1479),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1491),
.B(n_1563),
.Y(n_1698)
);

AND2x2_ASAP7_75t_SL g1699 ( 
.A(n_1621),
.B(n_1580),
.Y(n_1699)
);

AO31x2_ASAP7_75t_L g1700 ( 
.A1(n_1501),
.A2(n_1523),
.A3(n_1589),
.B(n_1566),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1546),
.A2(n_1531),
.B(n_1591),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1491),
.B(n_1514),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1546),
.B(n_1498),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1480),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1527),
.A2(n_1497),
.B(n_1483),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1482),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1484),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1570),
.A2(n_1620),
.B(n_1606),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1557),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1500),
.Y(n_1710)
);

AO21x2_ASAP7_75t_L g1711 ( 
.A1(n_1476),
.A2(n_1612),
.B(n_1600),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1530),
.A2(n_1610),
.B(n_1561),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1530),
.A2(n_1610),
.B(n_1561),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1535),
.B(n_1614),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1553),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1478),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1548),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1548),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1525),
.B(n_1539),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1553),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1525),
.B(n_1539),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1559),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1558),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1568),
.B(n_1541),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1533),
.A2(n_1560),
.B(n_1532),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1554),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1636),
.B(n_1640),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1647),
.Y(n_1728)
);

AOI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1645),
.A2(n_1584),
.B(n_1576),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1637),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1680),
.B(n_1582),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1707),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1629),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1676),
.B(n_1573),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1629),
.Y(n_1735)
);

NAND2x1_ASAP7_75t_L g1736 ( 
.A(n_1643),
.B(n_1521),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1541),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1632),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1640),
.B(n_1541),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1647),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1664),
.B(n_1592),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1658),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1714),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1694),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1668),
.Y(n_1745)
);

AND2x4_ASAP7_75t_SL g1746 ( 
.A(n_1643),
.B(n_1671),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1656),
.B(n_1574),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1628),
.B(n_1568),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1654),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1650),
.B(n_1537),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1664),
.B(n_1496),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1655),
.B(n_1496),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1655),
.B(n_1496),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1649),
.B(n_1537),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1718),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1635),
.B(n_1592),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1668),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1666),
.B(n_1672),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1666),
.B(n_1587),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1666),
.B(n_1581),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1710),
.B(n_1587),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1635),
.B(n_1590),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1679),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1652),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1638),
.B(n_1588),
.C(n_1551),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1663),
.B(n_1595),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1652),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1708),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1642),
.A2(n_1562),
.B1(n_1469),
.B2(n_1472),
.Y(n_1772)
);

INVx3_ASAP7_75t_SL g1773 ( 
.A(n_1625),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1672),
.B(n_1593),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1708),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1681),
.A2(n_1516),
.B1(n_1469),
.B2(n_1564),
.Y(n_1776)
);

NAND2x1_ASAP7_75t_L g1777 ( 
.A(n_1643),
.B(n_1494),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1672),
.B(n_1524),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1672),
.B(n_1524),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1634),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1708),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1648),
.A2(n_1613),
.B1(n_1485),
.B2(n_1572),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1708),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1667),
.B(n_1552),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1639),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1641),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1639),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1644),
.B(n_1613),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1646),
.B(n_1485),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1667),
.B(n_1552),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1698),
.B(n_1552),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1653),
.A2(n_1543),
.B1(n_1572),
.B2(n_1472),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1665),
.B(n_1556),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1698),
.B(n_1583),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1678),
.B(n_1543),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1674),
.B(n_1529),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1683),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1772),
.A2(n_1701),
.B1(n_1653),
.B2(n_1696),
.C(n_1626),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1743),
.B(n_1684),
.Y(n_1799)
);

NOR3xp33_ASAP7_75t_SL g1800 ( 
.A(n_1792),
.B(n_1528),
.C(n_1689),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1767),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1768),
.A2(n_1669),
.B1(n_1702),
.B2(n_1633),
.C(n_1709),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1747),
.A2(n_1669),
.B1(n_1702),
.B2(n_1686),
.C(n_1653),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1733),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1729),
.B(n_1782),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1737),
.B(n_1703),
.C(n_1725),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_L g1807 ( 
.A(n_1776),
.B(n_1529),
.C(n_1716),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1796),
.B(n_1703),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1732),
.B(n_1723),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1780),
.B(n_1786),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1697),
.B1(n_1695),
.B2(n_1706),
.C(n_1704),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1751),
.B(n_1696),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1761),
.B(n_1686),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1727),
.B(n_1699),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1657),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1752),
.B(n_1657),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1727),
.B(n_1699),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1748),
.B(n_1662),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1726),
.A2(n_1696),
.B1(n_1643),
.B2(n_1671),
.C(n_1662),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1748),
.B(n_1624),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1758),
.B(n_1624),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1762),
.B(n_1624),
.Y(n_1822)
);

XNOR2xp5_ASAP7_75t_L g1823 ( 
.A(n_1738),
.B(n_1528),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1793),
.B(n_1734),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1746),
.A2(n_1687),
.B(n_1685),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1762),
.B(n_1671),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1659),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1745),
.B(n_1671),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1745),
.B(n_1671),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1760),
.B(n_1715),
.Y(n_1830)
);

NOR3xp33_ASAP7_75t_L g1831 ( 
.A(n_1788),
.B(n_1529),
.C(n_1716),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1726),
.B(n_1725),
.C(n_1705),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1760),
.B(n_1715),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1734),
.B(n_1659),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1766),
.B(n_1720),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1730),
.B(n_1660),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1774),
.B(n_1765),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1789),
.A2(n_1700),
.B1(n_1627),
.B2(n_1631),
.C(n_1704),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1796),
.A2(n_1626),
.B1(n_1519),
.B2(n_1515),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1731),
.B(n_1515),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1774),
.B(n_1660),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1765),
.B(n_1661),
.Y(n_1842)
);

AND2x2_ASAP7_75t_SL g1843 ( 
.A(n_1746),
.B(n_1658),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1766),
.B(n_1720),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1764),
.B(n_1661),
.Y(n_1845)
);

OAI21xp33_ASAP7_75t_L g1846 ( 
.A1(n_1746),
.A2(n_1627),
.B(n_1721),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1795),
.B(n_1725),
.C(n_1705),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1728),
.B(n_1740),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1791),
.B(n_1739),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1791),
.B(n_1679),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1736),
.A2(n_1712),
.B(n_1713),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1749),
.B(n_1515),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_R g1853 ( 
.A(n_1795),
.B(n_1534),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1767),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1771),
.A2(n_1781),
.B(n_1775),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1763),
.B(n_1697),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1741),
.A2(n_1519),
.B1(n_1631),
.B2(n_1651),
.Y(n_1857)
);

NAND3xp33_ASAP7_75t_L g1858 ( 
.A(n_1741),
.B(n_1725),
.C(n_1705),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1728),
.B(n_1689),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1763),
.A2(n_1724),
.B1(n_1631),
.B2(n_1674),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1753),
.A2(n_1721),
.B1(n_1719),
.B2(n_1722),
.C(n_1519),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1763),
.B(n_1711),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1863)
);

NAND3xp33_ASAP7_75t_L g1864 ( 
.A(n_1784),
.B(n_1705),
.C(n_1690),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_SL g1865 ( 
.A1(n_1796),
.A2(n_1688),
.B(n_1673),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1784),
.B(n_1690),
.C(n_1691),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1736),
.A2(n_1685),
.B1(n_1687),
.B2(n_1625),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1790),
.B(n_1691),
.C(n_1719),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1790),
.B(n_1677),
.C(n_1682),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1755),
.B(n_1693),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1778),
.B(n_1779),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1770),
.Y(n_1872)
);

NAND3xp33_ASAP7_75t_L g1873 ( 
.A(n_1759),
.B(n_1677),
.C(n_1682),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1801),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1820),
.B(n_1771),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1820),
.B(n_1775),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1824),
.B(n_1770),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1830),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1855),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1814),
.B(n_1817),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1851),
.B(n_1742),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1840),
.B(n_1852),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1831),
.B(n_1796),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1862),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1814),
.B(n_1755),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1854),
.Y(n_1886)
);

NAND2x1p5_ASAP7_75t_L g1887 ( 
.A(n_1843),
.B(n_1777),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1855),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1817),
.B(n_1756),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1849),
.B(n_1756),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1855),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1830),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1859),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1821),
.B(n_1837),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1859),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1872),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1804),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1810),
.B(n_1783),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1843),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.B(n_1822),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1808),
.B(n_1742),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1804),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1865),
.B(n_1873),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1822),
.B(n_1754),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1856),
.B(n_1759),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1808),
.B(n_1828),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1833),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1799),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1813),
.B(n_1754),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1806),
.B(n_1750),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1833),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1865),
.B(n_1847),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1845),
.B(n_1778),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1834),
.B(n_1785),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1818),
.B(n_1779),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1835),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1850),
.B(n_1744),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1842),
.B(n_1827),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1835),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1870),
.B(n_1744),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1870),
.B(n_1744),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1863),
.B(n_1787),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1815),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1874),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1924),
.B(n_1812),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1924),
.B(n_1871),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1899),
.B(n_1848),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1911),
.B(n_1841),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1899),
.B(n_1880),
.Y(n_1930)
);

OAI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1913),
.A2(n_1802),
.B(n_1805),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1879),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1874),
.Y(n_1933)
);

OAI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1913),
.A2(n_1805),
.B(n_1803),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1906),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1886),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1911),
.B(n_1832),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1909),
.B(n_1823),
.Y(n_1938)
);

NOR4xp75_ASAP7_75t_L g1939 ( 
.A(n_1883),
.B(n_1798),
.C(n_1857),
.D(n_1777),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1886),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1896),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1877),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1896),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1919),
.B(n_1809),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1880),
.B(n_1848),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1907),
.B(n_1848),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1904),
.A2(n_1838),
.B(n_1819),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1907),
.B(n_1844),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1919),
.B(n_1816),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1844),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1903),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1884),
.B(n_1811),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1898),
.Y(n_1953)
);

AND2x6_ASAP7_75t_SL g1954 ( 
.A(n_1882),
.B(n_1522),
.Y(n_1954)
);

NOR2x1p5_ASAP7_75t_SL g1955 ( 
.A(n_1879),
.B(n_1888),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1907),
.B(n_1901),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1875),
.B(n_1864),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1875),
.B(n_1858),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1877),
.B(n_1868),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1915),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1901),
.B(n_1826),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1921),
.B(n_1826),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1903),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1921),
.B(n_1828),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1906),
.B(n_1836),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1904),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1900),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1898),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1878),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1923),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1914),
.B(n_1861),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1923),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1892),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1897),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1922),
.B(n_1829),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1905),
.B(n_1757),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1897),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1918),
.B(n_1825),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1918),
.B(n_1867),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1932),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1925),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1925),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1933),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1935),
.B(n_1894),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1954),
.B(n_1885),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1933),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1931),
.A2(n_1934),
.B1(n_1947),
.B2(n_1966),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1932),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1934),
.B(n_1905),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1954),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1936),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1956),
.B(n_1881),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1931),
.B(n_1910),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1965),
.B(n_1894),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1971),
.B(n_1910),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1974),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1956),
.B(n_1881),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1936),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1940),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1940),
.Y(n_2000)
);

INVx3_ASAP7_75t_SL g2001 ( 
.A(n_1967),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1952),
.B(n_1890),
.Y(n_2002)
);

NOR2x1p5_ASAP7_75t_L g2003 ( 
.A(n_1930),
.B(n_1900),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1941),
.Y(n_2004)
);

NAND2x1p5_ASAP7_75t_L g2005 ( 
.A(n_1969),
.B(n_1928),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1941),
.Y(n_2006)
);

AOI322xp5_ASAP7_75t_L g2007 ( 
.A1(n_1938),
.A2(n_1807),
.A3(n_1878),
.B1(n_1917),
.B2(n_1912),
.C1(n_1920),
.C2(n_1908),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1943),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1928),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1943),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1944),
.B(n_1885),
.Y(n_2011)
);

A2O1A1Ixp33_ASAP7_75t_L g2012 ( 
.A1(n_1939),
.A2(n_1800),
.B(n_1839),
.C(n_1881),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1949),
.B(n_1889),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1951),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1951),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1926),
.B(n_1889),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1959),
.B(n_1890),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1963),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1929),
.B(n_1917),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1963),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1942),
.B(n_1916),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1974),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1930),
.B(n_1881),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1937),
.B(n_1866),
.C(n_1869),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1946),
.B(n_1978),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1973),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1937),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1977),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1960),
.B(n_1916),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1946),
.B(n_1900),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1969),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_1958),
.A2(n_1853),
.B1(n_1724),
.B2(n_1794),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1958),
.B(n_1953),
.Y(n_2033)
);

NOR3xp33_ASAP7_75t_SL g2034 ( 
.A(n_1939),
.B(n_1823),
.C(n_1927),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2005),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2005),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_2033),
.B(n_1957),
.Y(n_2037)
);

INVx4_ASAP7_75t_L g2038 ( 
.A(n_2001),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2003),
.B(n_1978),
.Y(n_2039)
);

CKINVDCx16_ASAP7_75t_R g2040 ( 
.A(n_1990),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2025),
.B(n_1968),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1981),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1980),
.Y(n_2043)
);

CKINVDCx16_ASAP7_75t_R g2044 ( 
.A(n_1987),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2027),
.B(n_1970),
.Y(n_2045)
);

BUFx3_ASAP7_75t_L g2046 ( 
.A(n_2001),
.Y(n_2046)
);

AND2x2_ASAP7_75t_SL g2047 ( 
.A(n_1985),
.B(n_1957),
.Y(n_2047)
);

AND4x1_ASAP7_75t_L g2048 ( 
.A(n_2034),
.B(n_1670),
.C(n_1544),
.D(n_1522),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2025),
.B(n_1948),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1982),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2026),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_2031),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1983),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1995),
.B(n_1970),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2023),
.B(n_1948),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1985),
.A2(n_1887),
.B1(n_1902),
.B2(n_1967),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1986),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_2033),
.Y(n_2058)
);

INVxp67_ASAP7_75t_L g2059 ( 
.A(n_1993),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1991),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2023),
.B(n_1950),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_2009),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1998),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1989),
.A2(n_1887),
.B1(n_1902),
.B2(n_1979),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_2009),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1999),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2002),
.B(n_1972),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2000),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2004),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_2012),
.B(n_2007),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2030),
.B(n_1950),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_2009),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_2012),
.B(n_2024),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_2006),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_2030),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1984),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_1980),
.Y(n_2077)
);

O2A1O1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_2073),
.A2(n_2010),
.B(n_2008),
.C(n_2032),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2058),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_2070),
.A2(n_2032),
.B(n_2017),
.C(n_2015),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2044),
.B(n_2016),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_2058),
.Y(n_2082)
);

INVxp67_ASAP7_75t_SL g2083 ( 
.A(n_2051),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2044),
.A2(n_2059),
.B1(n_2052),
.B2(n_2051),
.C(n_2040),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_2072),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2042),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2047),
.A2(n_2016),
.B1(n_1992),
.B2(n_1997),
.Y(n_2087)
);

OAI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2048),
.A2(n_2019),
.B1(n_1887),
.B2(n_1994),
.C(n_2011),
.Y(n_2088)
);

AOI32xp33_ASAP7_75t_L g2089 ( 
.A1(n_2075),
.A2(n_1992),
.A3(n_1997),
.B1(n_2011),
.B2(n_2013),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_2040),
.Y(n_2090)
);

OAI32xp33_ASAP7_75t_L g2091 ( 
.A1(n_2075),
.A2(n_2021),
.A3(n_2029),
.B1(n_2014),
.B2(n_2020),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2042),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2052),
.B(n_2013),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2047),
.B(n_1972),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2072),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2037),
.B(n_2018),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_2047),
.A2(n_2059),
.B1(n_2076),
.B2(n_2046),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2062),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2056),
.A2(n_1902),
.B1(n_1929),
.B2(n_1979),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2049),
.B(n_1945),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2050),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2046),
.A2(n_1895),
.B1(n_1893),
.B2(n_1876),
.Y(n_2102)
);

OAI21xp33_ASAP7_75t_L g2103 ( 
.A1(n_2076),
.A2(n_1955),
.B(n_1846),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2062),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_2046),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2049),
.B(n_1945),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2041),
.B(n_1961),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2039),
.A2(n_1902),
.B1(n_1988),
.B2(n_1996),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2090),
.B(n_2049),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_2105),
.B(n_2038),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_2082),
.B(n_2038),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_2081),
.B(n_2093),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2095),
.B(n_2038),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2100),
.B(n_2039),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2083),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2084),
.B(n_2038),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2079),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2096),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2095),
.Y(n_2119)
);

INVx1_ASAP7_75t_SL g2120 ( 
.A(n_2096),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2086),
.Y(n_2121)
);

NAND2x1_ASAP7_75t_L g2122 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2097),
.B(n_2041),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_2094),
.Y(n_2124)
);

AOI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2097),
.A2(n_2037),
.B1(n_2035),
.B2(n_2036),
.C(n_2065),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2085),
.B(n_2041),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_2098),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2087),
.B(n_2071),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2104),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2100),
.B(n_2039),
.Y(n_2130)
);

OAI21xp33_ASAP7_75t_L g2131 ( 
.A1(n_2087),
.A2(n_2048),
.B(n_2064),
.Y(n_2131)
);

INVx1_ASAP7_75t_SL g2132 ( 
.A(n_2104),
.Y(n_2132)
);

OAI211xp5_ASAP7_75t_SL g2133 ( 
.A1(n_2116),
.A2(n_2088),
.B(n_2078),
.C(n_2080),
.Y(n_2133)
);

AOI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2125),
.A2(n_2091),
.B1(n_2089),
.B2(n_2103),
.C(n_2101),
.Y(n_2134)
);

AOI211xp5_ASAP7_75t_L g2135 ( 
.A1(n_2131),
.A2(n_2099),
.B(n_2102),
.C(n_2065),
.Y(n_2135)
);

OAI211xp5_ASAP7_75t_L g2136 ( 
.A1(n_2123),
.A2(n_2065),
.B(n_2108),
.C(n_2092),
.Y(n_2136)
);

O2A1O1Ixp5_ASAP7_75t_SL g2137 ( 
.A1(n_2119),
.A2(n_2050),
.B(n_2057),
.C(n_2053),
.Y(n_2137)
);

OAI21xp33_ASAP7_75t_L g2138 ( 
.A1(n_2128),
.A2(n_2107),
.B(n_2036),
.Y(n_2138)
);

OAI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_2112),
.A2(n_2045),
.B1(n_2036),
.B2(n_2035),
.C(n_2067),
.Y(n_2139)
);

AOI211xp5_ASAP7_75t_L g2140 ( 
.A1(n_2112),
.A2(n_2035),
.B(n_2045),
.C(n_2074),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_2115),
.A2(n_2074),
.B(n_2067),
.C(n_2071),
.Y(n_2141)
);

AOI211x1_ASAP7_75t_L g2142 ( 
.A1(n_2109),
.A2(n_2054),
.B(n_2106),
.C(n_2057),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_2124),
.A2(n_2074),
.B(n_2060),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2114),
.A2(n_2106),
.B1(n_2055),
.B2(n_2061),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2126),
.B(n_2054),
.Y(n_2145)
);

AOI211xp5_ASAP7_75t_L g2146 ( 
.A1(n_2110),
.A2(n_2060),
.B(n_2063),
.C(n_2053),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2122),
.A2(n_2066),
.B(n_2063),
.Y(n_2147)
);

AOI211xp5_ASAP7_75t_L g2148 ( 
.A1(n_2133),
.A2(n_2110),
.B(n_2111),
.C(n_2118),
.Y(n_2148)
);

NAND4xp25_ASAP7_75t_L g2149 ( 
.A(n_2135),
.B(n_2111),
.C(n_2117),
.D(n_2120),
.Y(n_2149)
);

NOR3xp33_ASAP7_75t_L g2150 ( 
.A(n_2136),
.B(n_2113),
.C(n_2127),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2140),
.B(n_2113),
.C(n_2121),
.Y(n_2151)
);

NOR2xp67_ASAP7_75t_SL g2152 ( 
.A(n_2143),
.B(n_1544),
.Y(n_2152)
);

NOR2x1_ASAP7_75t_L g2153 ( 
.A(n_2147),
.B(n_2113),
.Y(n_2153)
);

HB1xp67_ASAP7_75t_L g2154 ( 
.A(n_2141),
.Y(n_2154)
);

NOR3xp33_ASAP7_75t_SL g2155 ( 
.A(n_2138),
.B(n_2132),
.C(n_2129),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2146),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2145),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2142),
.B(n_2130),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2134),
.B(n_2055),
.Y(n_2159)
);

NOR3x1_ASAP7_75t_L g2160 ( 
.A(n_2149),
.B(n_2139),
.C(n_2077),
.Y(n_2160)
);

INVx1_ASAP7_75t_SL g2161 ( 
.A(n_2153),
.Y(n_2161)
);

AOI211xp5_ASAP7_75t_L g2162 ( 
.A1(n_2150),
.A2(n_2137),
.B(n_2144),
.C(n_2068),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2151),
.B(n_2066),
.Y(n_2163)
);

AND4x1_ASAP7_75t_L g2164 ( 
.A(n_2148),
.B(n_1538),
.C(n_1513),
.D(n_1512),
.Y(n_2164)
);

NAND3xp33_ASAP7_75t_L g2165 ( 
.A(n_2155),
.B(n_2154),
.C(n_2156),
.Y(n_2165)
);

NAND4xp25_ASAP7_75t_L g2166 ( 
.A(n_2159),
.B(n_2068),
.C(n_2069),
.D(n_2043),
.Y(n_2166)
);

OAI211xp5_ASAP7_75t_SL g2167 ( 
.A1(n_2157),
.A2(n_2069),
.B(n_2043),
.C(n_2077),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_L g2168 ( 
.A(n_2158),
.B(n_2077),
.C(n_2043),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2163),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2165),
.A2(n_2152),
.B1(n_2061),
.B2(n_1988),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2161),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_2164),
.B(n_1996),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2167),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2168),
.B(n_2022),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2166),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2160),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2162),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_2177),
.A2(n_2028),
.B1(n_2022),
.B2(n_1893),
.Y(n_2178)
);

NOR3xp33_ASAP7_75t_L g2179 ( 
.A(n_2176),
.B(n_2028),
.C(n_1470),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2170),
.A2(n_1977),
.B1(n_1895),
.B2(n_1876),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2169),
.B(n_1586),
.Y(n_2181)
);

NOR3xp33_ASAP7_75t_L g2182 ( 
.A(n_2171),
.B(n_1470),
.C(n_1716),
.Y(n_2182)
);

OAI211xp5_ASAP7_75t_SL g2183 ( 
.A1(n_2175),
.A2(n_1976),
.B(n_1891),
.C(n_1879),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2173),
.B(n_1961),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2184),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2181),
.Y(n_2186)
);

NOR2xp67_ASAP7_75t_L g2187 ( 
.A(n_2178),
.B(n_2174),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2179),
.Y(n_2188)
);

OAI22xp5_ASAP7_75t_SL g2189 ( 
.A1(n_2185),
.A2(n_2172),
.B1(n_2180),
.B2(n_2182),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2186),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2189),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2191),
.A2(n_2190),
.B1(n_2187),
.B2(n_2188),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2191),
.A2(n_2183),
.B1(n_2187),
.B2(n_1565),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2193),
.B(n_1955),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_2192),
.B(n_1964),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2195),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2194),
.A2(n_1891),
.B(n_1888),
.Y(n_2197)
);

OAI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_2196),
.A2(n_1962),
.B(n_1975),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_2198),
.A2(n_2197),
.B1(n_1891),
.B2(n_1888),
.Y(n_2199)
);

OAI221xp5_ASAP7_75t_R g2200 ( 
.A1(n_2199),
.A2(n_1860),
.B1(n_1565),
.B2(n_1670),
.C(n_1478),
.Y(n_2200)
);

AOI211xp5_ASAP7_75t_L g2201 ( 
.A1(n_2200),
.A2(n_1478),
.B(n_1494),
.C(n_1773),
.Y(n_2201)
);


endmodule