module fake_jpeg_25985_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_44),
.B1(n_36),
.B2(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_27),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_24),
.B1(n_25),
.B2(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_20),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AO21x1_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_14),
.B(n_22),
.Y(n_56)
);

OAI22x1_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_31),
.B(n_25),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_28),
.C(n_31),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_22),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_28),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_70),
.B(n_83),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_45),
.B1(n_32),
.B2(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_40),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_60),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_87),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_16),
.CI(n_33),
.CON(n_86),
.SN(n_86)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_91),
.B(n_18),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_12),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_89),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_84),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_67),
.B(n_1),
.C(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_76),
.B1(n_70),
.B2(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_80),
.B1(n_55),
.B2(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_86),
.B1(n_6),
.B2(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_89),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_73),
.B(n_52),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_94),
.B(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_119),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_86),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_106),
.B(n_108),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_11),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_99),
.C(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_3),
.C(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_114),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_117),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_125),
.C(n_2),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_64),
.B(n_133),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_135),
.B(n_132),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_64),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);


endmodule