module real_aes_8829_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_0), .A2(n_7), .B1(n_440), .B2(n_712), .C1(n_717), .C2(n_718), .Y(n_439) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_1), .B(n_85), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g433 ( .A(n_1), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_2), .A2(n_140), .B(n_145), .C(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_3), .A2(n_135), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g452 ( .A(n_4), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_5), .B(n_159), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_6), .B(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_7), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_8), .A2(n_135), .B(n_470), .Y(n_469) );
AND2x6_ASAP7_75t_L g140 ( .A(n_9), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g169 ( .A(n_10), .Y(n_169) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_11), .B(n_43), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_12), .A2(n_247), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_13), .B(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g474 ( .A(n_14), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_15), .B(n_149), .Y(n_522) );
INVx1_ASAP7_75t_L g133 ( .A(n_16), .Y(n_133) );
INVx1_ASAP7_75t_L g534 ( .A(n_17), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_18), .A2(n_170), .B(n_195), .C(n_197), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_19), .B(n_159), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_20), .B(n_463), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_21), .B(n_135), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_22), .B(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_23), .A2(n_149), .B(n_151), .C(n_155), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_24), .B(n_159), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_25), .B(n_150), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_26), .A2(n_153), .B(n_197), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_27), .B(n_150), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_28), .Y(n_215) );
INVx1_ASAP7_75t_L g229 ( .A(n_29), .Y(n_229) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_30), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_31), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_32), .B(n_150), .Y(n_453) );
INVx1_ASAP7_75t_L g252 ( .A(n_33), .Y(n_252) );
INVx1_ASAP7_75t_L g487 ( .A(n_34), .Y(n_487) );
INVx2_ASAP7_75t_L g138 ( .A(n_35), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_36), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_37), .A2(n_149), .B(n_208), .C(n_210), .Y(n_207) );
INVxp67_ASAP7_75t_L g253 ( .A(n_38), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_39), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_40), .A2(n_145), .B(n_228), .C(n_234), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_41), .A2(n_140), .B(n_145), .C(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_42), .A2(n_118), .B1(n_119), .B2(n_426), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_42), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_43), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g486 ( .A(n_44), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_45), .A2(n_167), .B(n_168), .C(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_46), .B(n_150), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_47), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_48), .Y(n_249) );
INVx1_ASAP7_75t_L g143 ( .A(n_49), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_50), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_51), .B(n_135), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_52), .A2(n_145), .B1(n_155), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_53), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_54), .Y(n_449) );
CKINVDCx14_ASAP7_75t_R g165 ( .A(n_55), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_56), .A2(n_167), .B(n_210), .C(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_57), .Y(n_515) );
INVx1_ASAP7_75t_L g471 ( .A(n_58), .Y(n_471) );
INVx1_ASAP7_75t_L g141 ( .A(n_59), .Y(n_141) );
INVx1_ASAP7_75t_L g132 ( .A(n_60), .Y(n_132) );
INVx1_ASAP7_75t_SL g209 ( .A(n_61), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_62), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_63), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g218 ( .A(n_64), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_SL g462 ( .A1(n_65), .A2(n_210), .B(n_463), .C(n_464), .Y(n_462) );
INVxp67_ASAP7_75t_L g465 ( .A(n_66), .Y(n_465) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_68), .A2(n_135), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_69), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_70), .A2(n_135), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_71), .Y(n_490) );
INVx1_ASAP7_75t_L g509 ( .A(n_72), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_73), .A2(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g193 ( .A(n_74), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_75), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_76), .A2(n_140), .B(n_145), .C(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_77), .A2(n_100), .B1(n_111), .B2(n_723), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_78), .A2(n_135), .B(n_142), .Y(n_134) );
INVx1_ASAP7_75t_L g196 ( .A(n_79), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_80), .B(n_230), .Y(n_503) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g183 ( .A(n_82), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_83), .B(n_463), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_84), .A2(n_140), .B(n_145), .C(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g430 ( .A(n_85), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g710 ( .A(n_85), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_85), .B(n_432), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_86), .A2(n_145), .B(n_217), .C(n_220), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_87), .B(n_162), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_88), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_89), .A2(n_140), .B(n_145), .C(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_90), .Y(n_526) );
INVx1_ASAP7_75t_L g461 ( .A(n_91), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_92), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_93), .B(n_230), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_94), .B(n_128), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_95), .B(n_128), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_98), .A2(n_135), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_SL g723 ( .A(n_102), .Y(n_723) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_438), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g722 ( .A(n_115), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_427), .B(n_435), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_120), .A2(n_441), .B1(n_709), .B2(n_711), .Y(n_440) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g716 ( .A(n_121), .Y(n_716) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_352), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_294), .C(n_324), .D(n_334), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_199), .B(n_257), .C(n_284), .Y(n_123) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_124), .A2(n_299), .B1(n_380), .B2(n_381), .C1(n_382), .C2(n_383), .Y(n_379) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_174), .Y(n_124) );
AOI33xp33_ASAP7_75t_L g305 ( .A1(n_125), .A2(n_292), .A3(n_293), .B1(n_306), .B2(n_311), .B3(n_313), .Y(n_305) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_125), .A2(n_363), .B(n_365), .C(n_367), .Y(n_362) );
OR2x2_ASAP7_75t_L g378 ( .A(n_125), .B(n_364), .Y(n_378) );
INVx1_ASAP7_75t_L g411 ( .A(n_125), .Y(n_411) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
INVx2_ASAP7_75t_L g288 ( .A(n_126), .Y(n_288) );
AND2x2_ASAP7_75t_L g304 ( .A(n_126), .B(n_190), .Y(n_304) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_126), .Y(n_339) );
AND2x2_ASAP7_75t_L g368 ( .A(n_126), .B(n_161), .Y(n_368) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_158), .Y(n_126) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_127), .A2(n_191), .B(n_198), .Y(n_190) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_127), .A2(n_204), .B(n_212), .Y(n_203) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_128), .A2(n_459), .B(n_466), .Y(n_458) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g245 ( .A(n_129), .Y(n_245) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_130), .B(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g247 ( .A(n_135), .Y(n_247) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_136), .B(n_140), .Y(n_180) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g233 ( .A(n_137), .Y(n_233) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx3_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
INVx1_ASAP7_75t_L g463 ( .A(n_139), .Y(n_463) );
INVx4_ASAP7_75t_SL g157 ( .A(n_140), .Y(n_157) );
BUFx3_ASAP7_75t_L g234 ( .A(n_140), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_157), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_144), .A2(n_157), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_144), .A2(n_157), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_144), .A2(n_157), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_144), .A2(n_157), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_144), .A2(n_157), .B(n_461), .C(n_462), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_144), .A2(n_157), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_144), .A2(n_157), .B(n_531), .C(n_532), .Y(n_530) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_149), .B(n_209), .Y(n_208) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_153), .B(n_196), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_153), .A2(n_230), .B1(n_252), .B2(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_153), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g485 ( .A1(n_154), .A2(n_185), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g454 ( .A(n_155), .Y(n_454) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_157), .A2(n_180), .B1(n_484), .B2(n_488), .Y(n_483) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_159), .A2(n_469), .B(n_475), .Y(n_468) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_160), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_214), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_160), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_160), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g268 ( .A(n_161), .Y(n_268) );
BUFx3_ASAP7_75t_L g276 ( .A(n_161), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_161), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_161), .B(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_161), .B(n_175), .Y(n_316) );
AND2x2_ASAP7_75t_L g385 ( .A(n_161), .B(n_319), .Y(n_385) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_173), .Y(n_161) );
INVx1_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx2_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_162), .A2(n_180), .B(n_226), .C(n_227), .Y(n_225) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_162), .A2(n_529), .B(n_535), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx5_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_170), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_170), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVx2_ASAP7_75t_SL g279 ( .A(n_174), .Y(n_279) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_175), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g321 ( .A(n_175), .Y(n_321) );
AND2x2_ASAP7_75t_L g332 ( .A(n_175), .B(n_288), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_175), .B(n_317), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_175), .B(n_319), .Y(n_364) );
AND2x2_ASAP7_75t_L g423 ( .A(n_175), .B(n_368), .Y(n_423) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g293 ( .A(n_176), .B(n_190), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g325 ( .A(n_176), .Y(n_325) );
AND3x2_ASAP7_75t_L g384 ( .A(n_176), .B(n_385), .C(n_386), .Y(n_384) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_177), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_177), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_177), .B(n_526), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_180), .A2(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_180), .A2(n_449), .B(n_450), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_180), .A2(n_509), .B(n_510), .Y(n_508) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_187), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_187), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_187), .A2(n_512), .B(n_513), .Y(n_511) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_190), .Y(n_275) );
INVx1_ASAP7_75t_SL g319 ( .A(n_190), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_190), .B(n_268), .C(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_237), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_200), .A2(n_303), .B(n_355), .C(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_202), .B(n_224), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_202), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g371 ( .A(n_202), .Y(n_371) );
AND2x2_ASAP7_75t_L g392 ( .A(n_202), .B(n_239), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_202), .B(n_301), .Y(n_420) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AND2x2_ASAP7_75t_L g265 ( .A(n_203), .B(n_256), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_203), .Y(n_272) );
AND2x2_ASAP7_75t_L g292 ( .A(n_203), .B(n_239), .Y(n_292) );
AND2x2_ASAP7_75t_L g342 ( .A(n_203), .B(n_224), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_203), .Y(n_346) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_211), .Y(n_523) );
INVx2_ASAP7_75t_SL g256 ( .A(n_213), .Y(n_256) );
BUFx2_ASAP7_75t_L g282 ( .A(n_213), .Y(n_282) );
AND2x2_ASAP7_75t_L g409 ( .A(n_213), .B(n_224), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_223), .A2(n_518), .B(n_525), .Y(n_517) );
INVx3_ASAP7_75t_SL g239 ( .A(n_224), .Y(n_239) );
AND2x2_ASAP7_75t_L g264 ( .A(n_224), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g271 ( .A(n_224), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g301 ( .A(n_224), .B(n_261), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_224), .B(n_256), .Y(n_310) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_224), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_224), .B(n_286), .Y(n_333) );
AND2x2_ASAP7_75t_L g361 ( .A(n_224), .B(n_241), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_224), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g399 ( .A(n_224), .B(n_240), .Y(n_399) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .C(n_232), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_230), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_233), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g323 ( .A(n_239), .B(n_272), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_239), .B(n_265), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_286), .Y(n_369) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_256), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_241), .B(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
OR2x2_ASAP7_75t_L g356 ( .A(n_241), .B(n_276), .Y(n_356) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_246), .B(n_254), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_262), .B(n_263), .Y(n_261) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_243), .A2(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g499 ( .A1(n_244), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_245), .A2(n_448), .B(n_455), .Y(n_447) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_245), .A2(n_483), .B(n_489), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_245), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_254), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_256), .B(n_261), .Y(n_291) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
AND2x2_ASAP7_75t_L g394 ( .A(n_256), .B(n_272), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_266), .B1(n_269), .B2(n_273), .C1(n_277), .C2(n_280), .Y(n_257) );
INVx1_ASAP7_75t_L g389 ( .A(n_258), .Y(n_389) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_259), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g296 ( .A(n_259), .B(n_265), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_259), .B(n_287), .Y(n_312) );
OAI222xp33_ASAP7_75t_L g334 ( .A1(n_259), .A2(n_335), .B1(n_340), .B2(n_341), .C1(n_349), .C2(n_351), .Y(n_334) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g322 ( .A(n_261), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_261), .B(n_342), .Y(n_382) );
AND2x2_ASAP7_75t_L g393 ( .A(n_261), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_264), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_266), .B(n_317), .Y(n_380) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_268), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_268), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx3_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_271), .A2(n_374), .B(n_377), .C(n_379), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_271), .B(n_308), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_271), .B(n_291), .Y(n_413) );
AND2x2_ASAP7_75t_L g286 ( .A(n_272), .B(n_282), .Y(n_286) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_276), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g365 ( .A(n_276), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_304), .Y(n_404) );
INVx1_ASAP7_75t_L g416 ( .A(n_276), .Y(n_416) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_279), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g397 ( .A(n_282), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_287), .B(n_289), .C(n_293), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_315), .B1(n_330), .B2(n_333), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_286), .B(n_300), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_286), .B(n_308), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_287), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g350 ( .A(n_287), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_287), .B(n_337), .Y(n_357) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NOR4xp25_ASAP7_75t_L g295 ( .A(n_292), .B(n_296), .C(n_297), .D(n_300), .Y(n_295) );
INVx1_ASAP7_75t_SL g366 ( .A(n_293), .Y(n_366) );
AND2x2_ASAP7_75t_L g410 ( .A(n_293), .B(n_411), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_302), .B(n_305), .C(n_314), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_301), .B(n_371), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_303), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
INVx1_ASAP7_75t_SL g376 ( .A(n_304), .Y(n_376) );
AND2x2_ASAP7_75t_L g415 ( .A(n_304), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_308), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_313), .B(n_338), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_320), .B(n_322), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g390 ( .A(n_317), .Y(n_390) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g418 ( .A(n_318), .Y(n_418) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B(n_329), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_325), .Y(n_337) );
OR2x2_ASAP7_75t_L g375 ( .A(n_325), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_328), .A2(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_332), .A2(n_359), .B1(n_362), .B2(n_369), .C(n_370), .Y(n_358) );
INVx1_ASAP7_75t_SL g402 ( .A(n_333), .Y(n_402) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g349 ( .A(n_337), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_346), .B2(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g381 ( .A(n_342), .Y(n_381) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_345), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_387), .C(n_400), .D(n_412), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_358), .C(n_373), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_356), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_363), .B(n_368), .Y(n_372) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_375), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_405), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_377), .A2(n_392), .B(n_393), .C(n_395), .Y(n_391) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_395) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_390), .C(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g406 ( .A(n_399), .Y(n_406) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_417), .B2(n_419), .C(n_421), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_431), .B(n_710), .Y(n_720) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g709 ( .A(n_432), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_435), .A2(n_439), .B(n_721), .Y(n_438) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g713 ( .A(n_441), .Y(n_713) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_625), .Y(n_441) );
NOR5xp2_ASAP7_75t_L g442 ( .A(n_443), .B(n_548), .C(n_580), .D(n_595), .E(n_612), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_476), .B(n_495), .C(n_536), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_445), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_445), .B(n_600), .Y(n_663) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_446), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_446), .B(n_492), .Y(n_549) );
AND2x2_ASAP7_75t_L g590 ( .A(n_446), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_446), .B(n_559), .Y(n_594) );
OR2x2_ASAP7_75t_L g631 ( .A(n_446), .B(n_482), .Y(n_631) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g481 ( .A(n_447), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g539 ( .A(n_447), .Y(n_539) );
OR2x2_ASAP7_75t_L g702 ( .A(n_447), .B(n_542), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_457), .A2(n_605), .B1(n_606), .B2(n_609), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_457), .B(n_539), .Y(n_688) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
AND2x2_ASAP7_75t_L g494 ( .A(n_458), .B(n_482), .Y(n_494) );
AND2x2_ASAP7_75t_L g541 ( .A(n_458), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
INVx3_ASAP7_75t_L g559 ( .A(n_458), .Y(n_559) );
OR2x2_ASAP7_75t_L g579 ( .A(n_458), .B(n_542), .Y(n_579) );
AND2x2_ASAP7_75t_L g598 ( .A(n_458), .B(n_468), .Y(n_598) );
BUFx2_ASAP7_75t_L g630 ( .A(n_458), .Y(n_630) );
AND2x4_ASAP7_75t_L g545 ( .A(n_467), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g480 ( .A(n_468), .Y(n_480) );
INVx2_ASAP7_75t_L g493 ( .A(n_468), .Y(n_493) );
OR2x2_ASAP7_75t_L g561 ( .A(n_468), .B(n_542), .Y(n_561) );
AND2x2_ASAP7_75t_L g591 ( .A(n_468), .B(n_482), .Y(n_591) );
AND2x2_ASAP7_75t_L g608 ( .A(n_468), .B(n_539), .Y(n_608) );
AND2x2_ASAP7_75t_L g648 ( .A(n_468), .B(n_559), .Y(n_648) );
AND2x2_ASAP7_75t_SL g684 ( .A(n_468), .B(n_494), .Y(n_684) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_478), .B(n_491), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_479), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_480), .A2(n_494), .B(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_480), .B(n_482), .Y(n_678) );
AND2x2_ASAP7_75t_L g614 ( .A(n_481), .B(n_615), .Y(n_614) );
INVx3_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_482), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_491), .B(n_539), .Y(n_707) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_492), .A2(n_650), .B1(n_651), .B2(n_656), .Y(n_649) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g540 ( .A(n_493), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g578 ( .A(n_493), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g615 ( .A(n_493), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_494), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g669 ( .A(n_494), .Y(n_669) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_516), .Y(n_496) );
INVx4_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
AND2x2_ASAP7_75t_L g633 ( .A(n_497), .B(n_600), .Y(n_633) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx3_ASAP7_75t_L g552 ( .A(n_498), .Y(n_552) );
AND2x2_ASAP7_75t_L g566 ( .A(n_498), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_498), .Y(n_570) );
INVx2_ASAP7_75t_L g584 ( .A(n_498), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_498), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g641 ( .A(n_498), .B(n_636), .Y(n_641) );
AND2x2_ASAP7_75t_L g706 ( .A(n_498), .B(n_676), .Y(n_706) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
AND2x2_ASAP7_75t_L g547 ( .A(n_507), .B(n_528), .Y(n_547) );
INVx2_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
INVx1_ASAP7_75t_L g572 ( .A(n_516), .Y(n_572) );
AND2x2_ASAP7_75t_L g618 ( .A(n_516), .B(n_566), .Y(n_618) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx2_ASAP7_75t_L g557 ( .A(n_517), .Y(n_557) );
INVx1_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_517), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_517), .B(n_567), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_557), .Y(n_600) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g553 ( .A(n_528), .Y(n_553) );
AND2x2_ASAP7_75t_L g636 ( .A(n_528), .B(n_567), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_543), .B(n_547), .Y(n_536) );
INVx1_ASAP7_75t_SL g581 ( .A(n_537), .Y(n_581) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_538), .B(n_545), .Y(n_638) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g587 ( .A(n_539), .B(n_542), .Y(n_587) );
AND2x2_ASAP7_75t_L g616 ( .A(n_539), .B(n_560), .Y(n_616) );
OR2x2_ASAP7_75t_L g619 ( .A(n_539), .B(n_579), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_540), .A2(n_632), .B1(n_684), .B2(n_685), .C1(n_687), .C2(n_689), .Y(n_683) );
BUFx2_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g586 ( .A(n_545), .B(n_587), .Y(n_586) );
INVx3_ASAP7_75t_SL g603 ( .A(n_545), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_545), .B(n_597), .Y(n_657) );
AND2x2_ASAP7_75t_L g592 ( .A(n_547), .B(n_552), .Y(n_592) );
INVx1_ASAP7_75t_L g611 ( .A(n_547), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_550), .B1(n_554), .B2(n_558), .C(n_562), .Y(n_548) );
OR2x2_ASAP7_75t_L g620 ( .A(n_550), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g605 ( .A(n_552), .B(n_575), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_552), .B(n_565), .Y(n_645) );
AND2x2_ASAP7_75t_L g650 ( .A(n_552), .B(n_600), .Y(n_650) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_552), .Y(n_660) );
NAND2x1_ASAP7_75t_SL g671 ( .A(n_552), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g556 ( .A(n_553), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g576 ( .A(n_553), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_553), .B(n_571), .Y(n_602) );
INVx1_ASAP7_75t_L g668 ( .A(n_553), .Y(n_668) );
INVx1_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g655 ( .A(n_555), .Y(n_655) );
NOR2xp67_ASAP7_75t_L g667 ( .A(n_555), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_556), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g575 ( .A(n_557), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_557), .B(n_567), .Y(n_588) );
INVx1_ASAP7_75t_L g654 ( .A(n_557), .Y(n_654) );
INVx1_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_568), .B(n_577), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x2_ASAP7_75t_L g708 ( .A(n_564), .B(n_641), .Y(n_708) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g676 ( .A(n_565), .B(n_636), .Y(n_676) );
AOI32xp33_ASAP7_75t_L g589 ( .A1(n_566), .A2(n_572), .A3(n_590), .B1(n_592), .B2(n_593), .Y(n_589) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_566), .A2(n_598), .A3(n_681), .B1(n_692), .B2(n_693), .C1(n_694), .C2(n_696), .Y(n_691) );
INVx2_ASAP7_75t_L g571 ( .A(n_567), .Y(n_571) );
INVx1_ASAP7_75t_L g681 ( .A(n_567), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B1(n_573), .B2(n_574), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_569), .B(n_575), .Y(n_624) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_570), .B(n_636), .Y(n_686) );
INVx1_ASAP7_75t_L g573 ( .A(n_571), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_571), .B(n_600), .Y(n_690) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_579), .B(n_674), .Y(n_673) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B1(n_585), .B2(n_588), .C(n_589), .Y(n_580) );
OR2x2_ASAP7_75t_L g601 ( .A(n_582), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g610 ( .A(n_582), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g635 ( .A(n_583), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g639 ( .A(n_593), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_599), .B1(n_601), .B2(n_603), .C(n_604), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_597), .A2(n_628), .B1(n_632), .B2(n_633), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_598), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_598), .Y(n_703) );
INVx1_ASAP7_75t_L g697 ( .A(n_600), .Y(n_697) );
INVx1_ASAP7_75t_SL g632 ( .A(n_601), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_603), .B(n_631), .Y(n_693) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_608), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g674 ( .A(n_608), .Y(n_674) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_617), .B1(n_619), .B2(n_620), .C(n_622), .Y(n_612) );
NOR2xp33_ASAP7_75t_SL g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_614), .A2(n_632), .B1(n_678), .B2(n_679), .Y(n_677) );
CKINVDCx14_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_619), .A2(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_658), .C(n_682), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_634), .C(n_642), .D(n_649), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g705 ( .A(n_630), .Y(n_705) );
INVx3_ASAP7_75t_SL g699 ( .A(n_631), .Y(n_699) );
OR2x2_ASAP7_75t_L g704 ( .A(n_631), .B(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_639), .B2(n_641), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_636), .B(n_654), .Y(n_695) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B(n_646), .Y(n_642) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_661), .B(n_664), .C(n_677), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g692 ( .A(n_663), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_669), .B1(n_670), .B2(n_673), .C1(n_675), .C2(n_676), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND4xp25_ASAP7_75t_SL g701 ( .A(n_674), .B(n_702), .C(n_703), .D(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_691), .C(n_700), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_711), .Y(n_715) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
endmodule