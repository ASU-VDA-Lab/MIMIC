module fake_jpeg_26358_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_8),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_47),
.Y(n_66)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_8),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_59),
.B1(n_19),
.B2(n_28),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_33),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_42),
.C(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_67),
.C(n_72),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_22),
.B1(n_45),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_17),
.B(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_23),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_19),
.B1(n_27),
.B2(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_26),
.C(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_74),
.B(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_103),
.B1(n_55),
.B2(n_49),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_92),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_24),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.C(n_68),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_64),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_95),
.B1(n_55),
.B2(n_49),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_20),
.B1(n_17),
.B2(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_20),
.B1(n_35),
.B2(n_2),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_8),
.B1(n_1),
.B2(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_100),
.Y(n_122)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_0),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_9),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_83),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_83),
.B1(n_91),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_57),
.CI(n_55),
.CON(n_123),
.SN(n_123)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_87),
.A3(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_126),
.B1(n_73),
.B2(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_0),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_79),
.B(n_88),
.Y(n_151)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_111),
.B(n_123),
.C(n_128),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_84),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_78),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_76),
.B(n_84),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_142),
.B(n_145),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_147),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_73),
.B(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_75),
.B1(n_97),
.B2(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_152),
.B1(n_142),
.B2(n_147),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_79),
.C(n_94),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_150),
.C(n_107),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_79),
.C(n_94),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_102),
.B1(n_85),
.B2(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_5),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_155),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_87),
.B1(n_102),
.B2(n_12),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_131),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_162),
.B1(n_136),
.B2(n_110),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_167),
.C(n_151),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_107),
.C(n_112),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_123),
.B(n_117),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_175),
.B(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_170),
.B(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_123),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_149),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_155),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_137),
.B(n_141),
.C(n_138),
.D(n_157),
.Y(n_180)
);

OAI322xp33_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_182),
.A3(n_191),
.B1(n_174),
.B2(n_175),
.C1(n_160),
.C2(n_179),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_153),
.Y(n_210)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_146),
.B1(n_134),
.B2(n_145),
.C(n_143),
.Y(n_182)
);

OA21x2_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_150),
.B(n_130),
.Y(n_183)
);

AOI321xp33_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_187),
.A3(n_161),
.B1(n_171),
.B2(n_167),
.C(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_135),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_171),
.C(n_108),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_176),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_192),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_110),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_161),
.B(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_159),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_196),
.A2(n_193),
.B1(n_194),
.B2(n_190),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_109),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_159),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_205),
.B(n_187),
.Y(n_217)
);

OAI321xp33_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_165),
.A3(n_161),
.B1(n_162),
.B2(n_169),
.C(n_160),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_189),
.B(n_184),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_204),
.B1(n_211),
.B2(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_170),
.B1(n_161),
.B2(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_197),
.C(n_188),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_181),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_132),
.B1(n_114),
.B2(n_106),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_214),
.B(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_222),
.C(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_195),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_203),
.B1(n_202),
.B2(n_211),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_218),
.B(n_205),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_186),
.B(n_192),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_180),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_204),
.C(n_208),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_185),
.C(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_227),
.C(n_228),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_222),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_209),
.B1(n_201),
.B2(n_132),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_129),
.C(n_114),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_106),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_221),
.B(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_225),
.C(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.C(n_129),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_115),
.B1(n_7),
.B2(n_12),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_5),
.B1(n_7),
.B2(n_13),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_237),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_242),
.C(n_5),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_234),
.B(n_14),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_14),
.C(n_15),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_15),
.Y(n_248)
);


endmodule