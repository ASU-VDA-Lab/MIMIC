module fake_ibex_556_n_1027 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_1027);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_1027;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_457;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_497;
wire n_243;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_929;
wire n_315;
wire n_604;
wire n_441;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_646;
wire n_448;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_662;
wire n_267;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_283;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_912;
wire n_890;
wire n_921;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_565;
wire n_424;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_159;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_20),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_28),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_51),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_10),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_27),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_78),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_68),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_47),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_39),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_27),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_55),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_56),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_22),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_46),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_141),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_49),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_74),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_31),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_67),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_63),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_85),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_54),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_97),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_30),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_26),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_108),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_66),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_14),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_53),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_59),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_7),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_52),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_17),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_37),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_60),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_19),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_135),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_72),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_75),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_80),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_19),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_0),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_178),
.B(n_194),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_0),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_150),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_151),
.B(n_1),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_147),
.A2(n_65),
.B(n_139),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_189),
.B(n_1),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_2),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g271 ( 
.A1(n_147),
.A2(n_69),
.B(n_131),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_3),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_4),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_4),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_6),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_179),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_162),
.B(n_7),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_145),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_148),
.B(n_9),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_145),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_156),
.B(n_9),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_148),
.B(n_169),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_164),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_157),
.A2(n_187),
.B(n_180),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_183),
.B(n_11),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_161),
.B(n_82),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_175),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_165),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_12),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_166),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_168),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_188),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_172),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_228),
.B(n_12),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_173),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_161),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_145),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_174),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_188),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_176),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_227),
.B(n_13),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g314 ( 
.A1(n_157),
.A2(n_84),
.B(n_129),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_182),
.B(n_13),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_184),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_185),
.B(n_14),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_227),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_192),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_163),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_195),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_197),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_199),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_201),
.Y(n_325)
);

XOR2x2_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_15),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_15),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_252),
.B(n_232),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

OR2x2_ASAP7_75t_SL g334 ( 
.A(n_252),
.B(n_186),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_258),
.Y(n_337)
);

BUFx4f_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_259),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_265),
.B(n_163),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_254),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_258),
.B(n_254),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_262),
.A2(n_229),
.B1(n_190),
.B2(n_245),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_258),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_275),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_258),
.B(n_152),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_262),
.B(n_263),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_280),
.A2(n_237),
.B1(n_181),
.B2(n_241),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_270),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

AO21x2_ASAP7_75t_L g361 ( 
.A1(n_266),
.A2(n_247),
.B(n_246),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_280),
.B(n_196),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_287),
.B(n_155),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_263),
.B(n_180),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_276),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_264),
.B(n_171),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_264),
.B(n_187),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_274),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_274),
.B(n_205),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_275),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_155),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_288),
.A2(n_244),
.B1(n_212),
.B2(n_219),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_277),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_288),
.B(n_206),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_207),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_274),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_250),
.B(n_224),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_296),
.B(n_208),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_278),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_277),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_299),
.B(n_210),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx4_ASAP7_75t_SL g389 ( 
.A(n_291),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_256),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_250),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_256),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

AND2x4_ASAP7_75t_SL g397 ( 
.A(n_290),
.B(n_153),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_284),
.Y(n_398)
);

OR2x6_ASAP7_75t_L g399 ( 
.A(n_290),
.B(n_209),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_299),
.B(n_213),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_284),
.B(n_297),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_301),
.B(n_302),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_297),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_301),
.B(n_214),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_319),
.Y(n_406)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_291),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_302),
.B(n_216),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_291),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_303),
.B(n_215),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_306),
.B(n_159),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_306),
.B(n_217),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

BUFx4f_ASAP7_75t_L g419 ( 
.A(n_291),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_303),
.B(n_231),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_291),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_286),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_305),
.B(n_230),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_278),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

AO22x2_ASAP7_75t_L g426 ( 
.A1(n_326),
.A2(n_154),
.B1(n_242),
.B2(n_220),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_305),
.B(n_209),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_269),
.B(n_209),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_286),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_269),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_307),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_307),
.B(n_234),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_255),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_315),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_255),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_328),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_289),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_315),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_249),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_249),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_278),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_289),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_326),
.A2(n_191),
.B1(n_241),
.B2(n_153),
.Y(n_443)
);

AO21x2_ASAP7_75t_L g444 ( 
.A1(n_266),
.A2(n_240),
.B(n_236),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_272),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_255),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_291),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_278),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_310),
.B(n_203),
.Y(n_449)
);

AO22x1_ASAP7_75t_L g450 ( 
.A1(n_401),
.A2(n_181),
.B1(n_326),
.B2(n_272),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_343),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_330),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_430),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_338),
.B(n_261),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_343),
.B(n_273),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_345),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_329),
.B(n_310),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_347),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_312),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_345),
.B(n_312),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_316),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_391),
.A2(n_225),
.B1(n_211),
.B2(n_191),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_397),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_445),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_333),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_401),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_442),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_342),
.A2(n_266),
.B(n_314),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_338),
.B(n_261),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_316),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_438),
.B(n_317),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_356),
.B(n_317),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_359),
.B(n_360),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_320),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_337),
.B(n_320),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_355),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_355),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_367),
.B(n_322),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_436),
.A2(n_211),
.B1(n_225),
.B2(n_282),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_331),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_395),
.B(n_261),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_376),
.B(n_322),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_341),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_349),
.B(n_323),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_374),
.B(n_158),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_409),
.B(n_279),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_323),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_401),
.A2(n_318),
.B1(n_325),
.B2(n_324),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_447),
.B(n_279),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_341),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_350),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_374),
.A2(n_327),
.B(n_325),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_333),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_415),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_386),
.A2(n_327),
.B1(n_324),
.B2(n_294),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_404),
.B(n_251),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_368),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_390),
.A2(n_281),
.B1(n_295),
.B2(n_292),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_358),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_398),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_392),
.A2(n_281),
.B1(n_295),
.B2(n_292),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_332),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_385),
.B(n_251),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_394),
.B(n_253),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_398),
.B(n_253),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_339),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_353),
.B(n_257),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_368),
.B(n_314),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_363),
.A2(n_158),
.B1(n_159),
.B2(n_239),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_396),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_351),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_353),
.B(n_257),
.Y(n_538)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_340),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_363),
.A2(n_203),
.B1(n_239),
.B2(n_146),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_403),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_381),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_354),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_364),
.B(n_198),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_397),
.B(n_281),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_428),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_334),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_380),
.B(n_209),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_380),
.B(n_226),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_381),
.B(n_314),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_412),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_418),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_416),
.A2(n_292),
.B1(n_279),
.B2(n_294),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_369),
.B(n_193),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_336),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_451),
.B(n_486),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_453),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_486),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

BUFx6f_ASAP7_75t_SL g564 ( 
.A(n_507),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_473),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_482),
.A2(n_383),
.B1(n_336),
.B2(n_348),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_537),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_537),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_454),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_477),
.A2(n_383),
.B1(n_348),
.B2(n_371),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_471),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_495),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_454),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_510),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_478),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_524),
.B(n_426),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_527),
.B(n_416),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_533),
.A2(n_371),
.B1(n_379),
.B2(n_426),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_524),
.B(n_426),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_527),
.B(n_416),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_466),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_416),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_472),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

BUFx8_ASAP7_75t_L g592 ( 
.A(n_549),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_507),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_507),
.B(n_379),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_483),
.B(n_457),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_489),
.B(n_369),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_357),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_473),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_548),
.B(n_378),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_465),
.B(n_488),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_511),
.A2(n_411),
.B1(n_378),
.B2(n_382),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_558),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_479),
.A2(n_342),
.B(n_372),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_488),
.B(n_382),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_491),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_459),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_452),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_463),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_532),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_498),
.B(n_387),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_497),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_463),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

BUFx12f_ASAP7_75t_L g622 ( 
.A(n_518),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_545),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_467),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_467),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_467),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_467),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_470),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_462),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_535),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_544),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_469),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_497),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_458),
.A2(n_372),
.B1(n_405),
.B2(n_377),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_479),
.A2(n_444),
.B(n_361),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_547),
.B(n_387),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_469),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_450),
.B(n_411),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_485),
.B(n_509),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_544),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_475),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_533),
.A2(n_377),
.B1(n_432),
.B2(n_405),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_552),
.A2(n_433),
.B(n_446),
.Y(n_646)
);

AOI222xp33_ASAP7_75t_L g647 ( 
.A1(n_520),
.A2(n_375),
.B1(n_346),
.B2(n_432),
.C1(n_423),
.C2(n_420),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_546),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_529),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_501),
.B(n_346),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_475),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_529),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_546),
.A2(n_400),
.B1(n_408),
.B2(n_375),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_531),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_481),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_551),
.A2(n_400),
.B1(n_408),
.B2(n_423),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_542),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_481),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_513),
.B(n_389),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_474),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_501),
.B(n_420),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_591),
.A2(n_539),
.B1(n_494),
.B2(n_476),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_637),
.A2(n_506),
.B(n_512),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_635),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_556),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_575),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_582),
.A2(n_539),
.B1(n_494),
.B2(n_519),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_654),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_586),
.B(n_513),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_562),
.B(n_556),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_592),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_662),
.B(n_538),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_581),
.B(n_538),
.C(n_555),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_579),
.A2(n_584),
.B1(n_658),
.B2(n_581),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_571),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_588),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_561),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_503),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_595),
.B(n_553),
.Y(n_685)
);

INVx4_ASAP7_75t_SL g686 ( 
.A(n_654),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_650),
.A2(n_521),
.B1(n_517),
.B2(n_484),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_602),
.B(n_365),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_492),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_605),
.A2(n_493),
.B1(n_504),
.B2(n_519),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_592),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_597),
.B(n_554),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_605),
.A2(n_484),
.B1(n_515),
.B2(n_370),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_612),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_622),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_648),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_620),
.Y(n_698)
);

NAND4xp25_ASAP7_75t_L g699 ( 
.A(n_599),
.B(n_370),
.C(n_365),
.D(n_525),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_631),
.A2(n_597),
.B1(n_564),
.B2(n_594),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_564),
.A2(n_505),
.B1(n_552),
.B2(n_515),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_611),
.A2(n_517),
.B1(n_521),
.B2(n_490),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_594),
.A2(n_534),
.B1(n_314),
.B2(n_271),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_580),
.A2(n_505),
.B1(n_534),
.B2(n_444),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_568),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_608),
.B(n_456),
.Y(n_706)
);

NOR2x1_ASAP7_75t_SL g707 ( 
.A(n_593),
.B(n_485),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_583),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_616),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_589),
.B(n_455),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_637),
.A2(n_506),
.B(n_500),
.Y(n_711)
);

OAI21x1_ASAP7_75t_SL g712 ( 
.A1(n_583),
.A2(n_522),
.B(n_525),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_594),
.A2(n_455),
.B1(n_480),
.B2(n_522),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_646),
.A2(n_512),
.B(n_500),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_589),
.B(n_480),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_621),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_623),
.Y(n_717)
);

BUFx10_ASAP7_75t_L g718 ( 
.A(n_593),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_625),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_645),
.A2(n_559),
.B1(n_485),
.B2(n_509),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_638),
.A2(n_361),
.B1(n_294),
.B2(n_295),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_603),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_655),
.B(n_559),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_640),
.A2(n_530),
.B1(n_509),
.B2(n_485),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_593),
.B(n_389),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_645),
.A2(n_509),
.B1(n_530),
.B2(n_540),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_607),
.A2(n_271),
.B(n_543),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_619),
.B(n_435),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_633),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_638),
.B(n_16),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_647),
.B(n_410),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_SL g734 ( 
.A(n_625),
.B(n_407),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_618),
.A2(n_413),
.B(n_414),
.C(n_417),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_644),
.B(n_540),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_614),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_640),
.A2(n_530),
.B1(n_540),
.B2(n_271),
.Y(n_738)
);

AOI221xp5_ASAP7_75t_L g739 ( 
.A1(n_649),
.A2(n_652),
.B1(n_580),
.B2(n_585),
.C(n_629),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_613),
.B(n_18),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_640),
.A2(n_530),
.B1(n_421),
.B2(n_407),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_565),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_648),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_585),
.A2(n_540),
.B1(n_243),
.B2(n_407),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_606),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_596),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_610),
.B(n_389),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_604),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_SL g750 ( 
.A1(n_641),
.A2(n_557),
.B(n_543),
.C(n_536),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_636),
.A2(n_268),
.B1(n_283),
.B2(n_309),
.C(n_285),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_653),
.B(n_499),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_620),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_615),
.B(n_18),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_610),
.B(n_20),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_661),
.A2(n_271),
.B1(n_407),
.B2(n_421),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_590),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_657),
.A2(n_421),
.B1(n_268),
.B2(n_283),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_632),
.A2(n_421),
.B1(n_267),
.B2(n_283),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_566),
.A2(n_557),
.B(n_536),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_565),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_577),
.B(n_21),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_566),
.A2(n_570),
.B1(n_601),
.B2(n_577),
.Y(n_763)
);

OAI21xp33_ASAP7_75t_L g764 ( 
.A1(n_570),
.A2(n_523),
.B(n_514),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_601),
.B(n_21),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_569),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_632),
.B(n_22),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_587),
.B(n_523),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_569),
.A2(n_514),
.B(n_499),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_642),
.B(n_23),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_SL g771 ( 
.A1(n_642),
.A2(n_267),
.B1(n_268),
.B2(n_283),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_573),
.A2(n_268),
.B(n_309),
.C(n_285),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_573),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_587),
.A2(n_267),
.B1(n_285),
.B2(n_309),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_660),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_578),
.Y(n_776)
);

OAI21xp33_ASAP7_75t_SL g777 ( 
.A1(n_598),
.A2(n_298),
.B(n_309),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_598),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_660),
.Y(n_779)
);

CKINVDCx6p67_ASAP7_75t_R g780 ( 
.A(n_625),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_630),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_630),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_643),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_669),
.B(n_641),
.C(n_278),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_689),
.B(n_643),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_651),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_681),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_700),
.B(n_578),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_780),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_691),
.A2(n_659),
.B1(n_656),
.B2(n_651),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_SL g791 ( 
.A1(n_775),
.A2(n_578),
.B(n_628),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_698),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_691),
.A2(n_659),
.B1(n_656),
.B2(n_625),
.Y(n_793)
);

OAI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_672),
.A2(n_285),
.B(n_298),
.C(n_626),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_753),
.Y(n_795)
);

CKINVDCx6p67_ASAP7_75t_R g796 ( 
.A(n_692),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_676),
.A2(n_578),
.B1(n_639),
.B2(n_634),
.Y(n_797)
);

O2A1O1Ixp5_ASAP7_75t_L g798 ( 
.A1(n_728),
.A2(n_626),
.B(n_298),
.C(n_600),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_684),
.A2(n_639),
.B1(n_634),
.B2(n_600),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_732),
.A2(n_639),
.B1(n_634),
.B2(n_609),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_720),
.B(n_624),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_699),
.A2(n_639),
.B1(n_634),
.B2(n_609),
.Y(n_802)
);

NOR2x1_ASAP7_75t_L g803 ( 
.A(n_696),
.B(n_628),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_679),
.A2(n_624),
.B1(n_617),
.B2(n_614),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

AOI221xp5_ASAP7_75t_L g806 ( 
.A1(n_724),
.A2(n_311),
.B1(n_293),
.B2(n_300),
.C(n_304),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_707),
.A2(n_660),
.B1(n_624),
.B2(n_617),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_677),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_680),
.A2(n_660),
.B1(n_624),
.B2(n_617),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_679),
.A2(n_660),
.B1(n_617),
.B2(n_614),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_682),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_754),
.B(n_23),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_703),
.A2(n_448),
.B(n_441),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_677),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_739),
.A2(n_267),
.B1(n_293),
.B2(n_300),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_763),
.A2(n_267),
.B1(n_293),
.B2(n_300),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_763),
.A2(n_267),
.B1(n_293),
.B2(n_300),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_720),
.B(n_24),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_685),
.A2(n_267),
.B1(n_293),
.B2(n_300),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_666),
.Y(n_820)
);

AOI221xp5_ASAP7_75t_L g821 ( 
.A1(n_695),
.A2(n_293),
.B1(n_300),
.B2(n_304),
.C(n_311),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_694),
.A2(n_701),
.B1(n_670),
.B2(n_702),
.Y(n_822)
);

CKINVDCx6p67_ASAP7_75t_R g823 ( 
.A(n_690),
.Y(n_823)
);

AOI21xp33_ASAP7_75t_L g824 ( 
.A1(n_733),
.A2(n_24),
.B(n_25),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_737),
.Y(n_825)
);

AOI21xp33_ASAP7_75t_L g826 ( 
.A1(n_664),
.A2(n_25),
.B(n_311),
.Y(n_826)
);

OR2x6_ASAP7_75t_L g827 ( 
.A(n_667),
.B(n_304),
.Y(n_827)
);

AO221x1_ASAP7_75t_L g828 ( 
.A1(n_703),
.A2(n_311),
.B1(n_304),
.B2(n_41),
.C(n_44),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_686),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_737),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_737),
.Y(n_831)
);

OAI211xp5_ASAP7_75t_L g832 ( 
.A1(n_694),
.A2(n_304),
.B(n_311),
.C(n_424),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_693),
.A2(n_304),
.B1(n_311),
.B2(n_424),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_683),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_755),
.A2(n_448),
.B1(n_441),
.B2(n_424),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_671),
.A2(n_448),
.B1(n_441),
.B2(n_388),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_741),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_674),
.A2(n_388),
.B(n_384),
.C(n_373),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_SL g839 ( 
.A1(n_705),
.A2(n_32),
.B1(n_36),
.B2(n_50),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_721),
.B(n_57),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_674),
.A2(n_777),
.B(n_735),
.C(n_668),
.Y(n_841)
);

AOI21xp33_ASAP7_75t_L g842 ( 
.A1(n_690),
.A2(n_58),
.B(n_76),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_706),
.A2(n_688),
.B1(n_704),
.B2(n_687),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_388),
.B1(n_384),
.B2(n_373),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_SL g845 ( 
.A1(n_744),
.A2(n_77),
.B1(n_86),
.B2(n_88),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_709),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_686),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_762),
.A2(n_384),
.B1(n_373),
.B2(n_366),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_673),
.B(n_89),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_716),
.A2(n_366),
.B1(n_362),
.B2(n_352),
.C(n_344),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_717),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_765),
.A2(n_366),
.B1(n_362),
.B2(n_352),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_725),
.A2(n_362),
.B1(n_352),
.B2(n_344),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_773),
.A2(n_344),
.B1(n_335),
.B2(n_93),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_719),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_725),
.B(n_90),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_746),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_767),
.A2(n_335),
.B1(n_98),
.B2(n_102),
.Y(n_858)
);

OAI221xp5_ASAP7_75t_L g859 ( 
.A1(n_713),
.A2(n_335),
.B1(n_106),
.B2(n_110),
.C(n_113),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_726),
.A2(n_91),
.B1(n_114),
.B2(n_115),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_712),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_710),
.A2(n_126),
.B1(n_127),
.B2(n_140),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_777),
.B(n_723),
.C(n_751),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_731),
.B(n_749),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_738),
.A2(n_766),
.B1(n_778),
.B2(n_782),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_729),
.A2(n_723),
.B(n_665),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_L g867 ( 
.A1(n_752),
.A2(n_764),
.B(n_770),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_727),
.B(n_708),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_747),
.A2(n_715),
.B1(n_710),
.B2(n_722),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_715),
.B1(n_718),
.B2(n_697),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_697),
.A2(n_715),
.B1(n_757),
.B2(n_708),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_730),
.B(n_718),
.Y(n_872)
);

INVx3_ASAP7_75t_SL g873 ( 
.A(n_796),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_805),
.B(n_761),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_866),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_834),
.B(n_783),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_866),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_820),
.B(n_743),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_825),
.Y(n_879)
);

OR2x2_ASAP7_75t_SL g880 ( 
.A(n_829),
.B(n_741),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_L g881 ( 
.A1(n_787),
.A2(n_771),
.B1(n_772),
.B2(n_774),
.C(n_736),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_857),
.B(n_781),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_824),
.B(n_776),
.C(n_768),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_818),
.A2(n_727),
.B1(n_743),
.B2(n_764),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_846),
.Y(n_885)
);

AOI221xp5_ASAP7_75t_L g886 ( 
.A1(n_851),
.A2(n_758),
.B1(n_760),
.B2(n_711),
.C(n_714),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_855),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_788),
.A2(n_748),
.B1(n_745),
.B2(n_756),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_822),
.A2(n_843),
.B1(n_785),
.B2(n_869),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_825),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_811),
.B(n_741),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_792),
.A2(n_748),
.B1(n_742),
.B2(n_779),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_795),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_864),
.B(n_769),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_825),
.Y(n_895)
);

OAI322xp33_ASAP7_75t_L g896 ( 
.A1(n_812),
.A2(n_734),
.A3(n_750),
.B1(n_759),
.B2(n_779),
.C1(n_786),
.C2(n_845),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_790),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_869),
.A2(n_809),
.B1(n_856),
.B2(n_871),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_872),
.Y(n_899)
);

OAI211xp5_ASAP7_75t_L g900 ( 
.A1(n_870),
.A2(n_847),
.B(n_803),
.C(n_849),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_784),
.B(n_819),
.C(n_841),
.Y(n_902)
);

OAI21xp33_ASAP7_75t_SL g903 ( 
.A1(n_828),
.A2(n_810),
.B(n_790),
.Y(n_903)
);

NAND4xp25_ASAP7_75t_L g904 ( 
.A(n_847),
.B(n_814),
.C(n_808),
.D(n_816),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_856),
.B(n_801),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_823),
.B(n_868),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_865),
.Y(n_907)
);

OA21x2_ASAP7_75t_L g908 ( 
.A1(n_813),
.A2(n_867),
.B(n_832),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_802),
.B(n_815),
.C(n_826),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_810),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_863),
.A2(n_794),
.B1(n_793),
.B2(n_814),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_807),
.A2(n_842),
.B(n_862),
.Y(n_913)
);

OAI211xp5_ASAP7_75t_SL g914 ( 
.A1(n_817),
.A2(n_799),
.B(n_833),
.C(n_861),
.Y(n_914)
);

AOI222xp33_ASAP7_75t_L g915 ( 
.A1(n_839),
.A2(n_868),
.B1(n_860),
.B2(n_867),
.C1(n_840),
.C2(n_859),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_827),
.A2(n_800),
.B1(n_858),
.B2(n_852),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_830),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_827),
.B(n_837),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_827),
.B(n_837),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_797),
.B(n_791),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_830),
.B(n_837),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_SL g922 ( 
.A1(n_836),
.A2(n_804),
.B(n_848),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_830),
.B(n_831),
.Y(n_923)
);

NAND4xp25_ASAP7_75t_L g924 ( 
.A(n_889),
.B(n_806),
.C(n_821),
.D(n_798),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_923),
.B(n_831),
.Y(n_925)
);

AOI33xp33_ASAP7_75t_L g926 ( 
.A1(n_885),
.A2(n_835),
.A3(n_853),
.B1(n_844),
.B2(n_850),
.B3(n_838),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_885),
.B(n_831),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_887),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_889),
.A2(n_854),
.B(n_903),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_893),
.B(n_899),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_887),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_909),
.Y(n_932)
);

AO221x2_ASAP7_75t_L g933 ( 
.A1(n_903),
.A2(n_913),
.B1(n_916),
.B2(n_902),
.C(n_920),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_874),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_898),
.A2(n_884),
.B1(n_905),
.B2(n_912),
.Y(n_935)
);

OAI31xp33_ASAP7_75t_L g936 ( 
.A1(n_900),
.A2(n_905),
.A3(n_904),
.B(n_914),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_882),
.B(n_894),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_875),
.Y(n_938)
);

NAND4xp75_ASAP7_75t_L g939 ( 
.A(n_898),
.B(n_906),
.C(n_873),
.D(n_894),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_SL g940 ( 
.A(n_918),
.B(n_919),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_923),
.B(n_911),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_882),
.B(n_876),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_878),
.Y(n_944)
);

AOI221xp5_ASAP7_75t_L g945 ( 
.A1(n_896),
.A2(n_901),
.B1(n_907),
.B2(n_881),
.C(n_897),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_897),
.B(n_907),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_875),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_880),
.B(n_911),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_877),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_880),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_891),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_891),
.B(n_877),
.Y(n_952)
);

AOI221xp5_ASAP7_75t_L g953 ( 
.A1(n_886),
.A2(n_909),
.B1(n_910),
.B2(n_883),
.C(n_892),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_909),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_922),
.A2(n_908),
.B(n_915),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_952),
.B(n_908),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_952),
.B(n_895),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_928),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_946),
.B(n_895),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_941),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_938),
.B(n_908),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_950),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_938),
.B(n_908),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_931),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_937),
.B(n_919),
.Y(n_965)
);

OAI31xp33_ASAP7_75t_L g966 ( 
.A1(n_936),
.A2(n_918),
.A3(n_888),
.B(n_873),
.Y(n_966)
);

AOI211xp5_ASAP7_75t_SL g967 ( 
.A1(n_955),
.A2(n_922),
.B(n_873),
.C(n_890),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_947),
.Y(n_968)
);

AOI31xp33_ASAP7_75t_L g969 ( 
.A1(n_948),
.A2(n_879),
.A3(n_890),
.B(n_917),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_941),
.B(n_879),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_960),
.B(n_941),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_960),
.B(n_947),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_969),
.B(n_932),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_957),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_957),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_965),
.B(n_944),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_965),
.B(n_951),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_968),
.Y(n_978)
);

OAI31xp33_ASAP7_75t_L g979 ( 
.A1(n_966),
.A2(n_935),
.A3(n_929),
.B(n_948),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_958),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_958),
.B(n_930),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_964),
.B(n_943),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_975),
.B(n_962),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_976),
.B(n_934),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_973),
.B(n_932),
.Y(n_986)
);

OAI211xp5_ASAP7_75t_SL g987 ( 
.A1(n_979),
.A2(n_966),
.B(n_967),
.C(n_962),
.Y(n_987)
);

XNOR2xp5_ASAP7_75t_L g988 ( 
.A(n_971),
.B(n_974),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_979),
.A2(n_967),
.B(n_939),
.Y(n_989)
);

OAI211xp5_ASAP7_75t_SL g990 ( 
.A1(n_981),
.A2(n_953),
.B(n_945),
.C(n_954),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_980),
.Y(n_991)
);

NOR2x1_ASAP7_75t_L g992 ( 
.A(n_982),
.B(n_932),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_991),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_983),
.Y(n_994)
);

AND3x4_ASAP7_75t_L g995 ( 
.A(n_992),
.B(n_933),
.C(n_970),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_985),
.Y(n_996)
);

XNOR2x1_ASAP7_75t_L g997 ( 
.A(n_988),
.B(n_971),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_980),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_986),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_989),
.A2(n_978),
.B(n_982),
.C(n_977),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_987),
.A2(n_933),
.B1(n_974),
.B2(n_972),
.Y(n_1001)
);

XOR2x2_ASAP7_75t_L g1002 ( 
.A(n_989),
.B(n_972),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_SL g1003 ( 
.A1(n_999),
.A2(n_933),
.B(n_969),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_999),
.B(n_956),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_990),
.C(n_924),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_998),
.Y(n_1006)
);

NAND4xp75_ASAP7_75t_L g1007 ( 
.A(n_1000),
.B(n_956),
.C(n_959),
.D(n_964),
.Y(n_1007)
);

NOR4xp25_ASAP7_75t_L g1008 ( 
.A(n_998),
.B(n_927),
.C(n_942),
.D(n_956),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1008),
.B(n_1001),
.Y(n_1009)
);

NAND4xp25_ASAP7_75t_L g1010 ( 
.A(n_1005),
.B(n_994),
.C(n_995),
.D(n_1002),
.Y(n_1010)
);

NAND4xp75_ASAP7_75t_L g1011 ( 
.A(n_1004),
.B(n_993),
.C(n_996),
.D(n_959),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_1003),
.A2(n_997),
.B1(n_968),
.B2(n_963),
.C(n_961),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_963),
.Y(n_1013)
);

NAND5xp2_ASAP7_75t_L g1014 ( 
.A(n_1009),
.B(n_1006),
.C(n_1007),
.D(n_961),
.E(n_963),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_961),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1011),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_1013),
.B(n_925),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_1016),
.B(n_970),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1015),
.Y(n_1019)
);

NOR4xp25_ASAP7_75t_L g1020 ( 
.A(n_1017),
.B(n_926),
.C(n_917),
.D(n_949),
.Y(n_1020)
);

OAI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_1014),
.B1(n_949),
.B2(n_940),
.C(n_926),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1018),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1018),
.A2(n_970),
.B1(n_925),
.B2(n_940),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_1022),
.A2(n_1019),
.B1(n_970),
.B2(n_925),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1024),
.Y(n_1025)
);

XNOR2xp5_ASAP7_75t_L g1026 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_1026),
.A2(n_1021),
.B(n_921),
.Y(n_1027)
);


endmodule