module fake_jpeg_19486_n_206 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_12),
.B1(n_21),
.B2(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_21),
.B1(n_12),
.B2(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_21),
.B1(n_12),
.B2(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_40),
.B1(n_28),
.B2(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_21),
.B1(n_12),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_46),
.B1(n_33),
.B2(n_25),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_31),
.C(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_30),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_53),
.B(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_14),
.B1(n_13),
.B2(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_52),
.Y(n_58)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_31),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_25),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_32),
.B1(n_24),
.B2(n_27),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_45),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_24),
.B1(n_36),
.B2(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_63),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_23),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_44),
.C(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_57),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_54),
.B1(n_41),
.B2(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_80),
.B1(n_85),
.B2(n_65),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_49),
.B1(n_42),
.B2(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_44),
.B1(n_46),
.B2(n_51),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_50),
.B(n_53),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_72),
.B(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_104),
.B1(n_51),
.B2(n_56),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_65),
.C(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_100),
.C(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_75),
.B(n_53),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_70),
.CI(n_58),
.CON(n_99),
.SN(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_70),
.C(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_59),
.B1(n_70),
.B2(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_111),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_74),
.B1(n_85),
.B2(n_76),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_116),
.B1(n_90),
.B2(n_16),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_122),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_82),
.B(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_60),
.B1(n_49),
.B2(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_49),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_29),
.B1(n_11),
.B2(n_20),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_15),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_118),
.B1(n_114),
.B2(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_9),
.C(n_10),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_9),
.C(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_84),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_103),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_56),
.B1(n_62),
.B2(n_90),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_141),
.B1(n_116),
.B2(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_16),
.B1(n_17),
.B2(n_2),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_29),
.C(n_11),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_108),
.C(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_112),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_29),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_152),
.B1(n_158),
.B2(n_136),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_106),
.B(n_120),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_20),
.B(n_19),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_112),
.C(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_126),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_29),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_129),
.B1(n_131),
.B2(n_117),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_139),
.B1(n_132),
.B2(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_165),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_140),
.B1(n_133),
.B2(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_168),
.B(n_0),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_154),
.C(n_153),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_177),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_147),
.B(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_167),
.B(n_161),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_13),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_168),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_153),
.B(n_9),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_182),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_18),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_165),
.B(n_162),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_169),
.C(n_22),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_20),
.B(n_19),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_19),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_18),
.B1(n_11),
.B2(n_10),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_1),
.C(n_4),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_22),
.B1(n_7),
.B2(n_2),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_22),
.C(n_1),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_185),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_197),
.A3(n_194),
.B1(n_22),
.B2(n_193),
.C1(n_5),
.C2(n_6),
.Y(n_200)
);

AOI321xp33_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_7),
.A3(n_22),
.B1(n_2),
.B2(n_3),
.C(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_4),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.C(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_7),
.Y(n_202)
);

OAI222xp33_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_22),
.C2(n_204),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_6),
.C(n_191),
.Y(n_206)
);


endmodule