module fake_jpeg_10216_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_48),
.B(n_71),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_59),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_34),
.B2(n_23),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_61),
.B1(n_69),
.B2(n_44),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_32),
.B1(n_34),
.B2(n_23),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_34),
.B1(n_26),
.B2(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_38),
.B1(n_44),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_83),
.B1(n_20),
.B2(n_16),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_44),
.B1(n_40),
.B2(n_35),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_82),
.B1(n_88),
.B2(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_22),
.B1(n_33),
.B2(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_29),
.B1(n_35),
.B2(n_31),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_90),
.B(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_40),
.B1(n_31),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_94),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_19),
.B1(n_27),
.B2(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_37),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_21),
.B1(n_17),
.B2(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_33),
.B1(n_22),
.B2(n_17),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_104),
.B1(n_45),
.B2(n_16),
.Y(n_141)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_109),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_56),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_41),
.B1(n_17),
.B2(n_24),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_119),
.Y(n_149)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_16),
.B1(n_20),
.B2(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_62),
.C(n_58),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_126),
.C(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_102),
.B1(n_108),
.B2(n_101),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_141),
.B1(n_16),
.B2(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_62),
.C(n_58),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_62),
.C(n_45),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_56),
.B1(n_65),
.B2(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_76),
.B1(n_98),
.B2(n_109),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_45),
.C(n_53),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_53),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_110),
.B(n_82),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_144),
.B(n_159),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_74),
.Y(n_144)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_111),
.Y(n_145)
);

OR2x2_ASAP7_75t_SL g187 ( 
.A(n_145),
.B(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_147),
.B(n_148),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_97),
.B1(n_103),
.B2(n_85),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_155),
.B1(n_162),
.B2(n_131),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_164),
.B1(n_167),
.B2(n_0),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_74),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_165),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_87),
.B1(n_74),
.B2(n_95),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_173),
.B1(n_141),
.B2(n_128),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_45),
.B(n_106),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_106),
.B(n_91),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_163),
.B(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_128),
.C(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_108),
.B1(n_104),
.B2(n_56),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_86),
.B1(n_52),
.B2(n_55),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_18),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_52),
.B1(n_16),
.B2(n_53),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_127),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_0),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_120),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_179),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_184),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_136),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_127),
.A3(n_119),
.B1(n_118),
.B2(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_117),
.B1(n_114),
.B2(n_140),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_144),
.B1(n_166),
.B2(n_161),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_145),
.B(n_152),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_133),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_193),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_205),
.B1(n_167),
.B2(n_153),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_200),
.B1(n_162),
.B2(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_165),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_137),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_204),
.C(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_0),
.C(n_2),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_3),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_220),
.B(n_209),
.C(n_183),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_199),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_223),
.B(n_225),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_158),
.C(n_149),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_217),
.C(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_149),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_156),
.B1(n_169),
.B2(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_163),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_163),
.B(n_4),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_8),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_200),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_176),
.A2(n_3),
.B(n_4),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_9),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_181),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_188),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_194),
.C(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_241),
.C(n_243),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_226),
.B(n_223),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_179),
.C(n_197),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_228),
.C(n_213),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_222),
.B(n_203),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_206),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_224),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_243),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.C(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_273),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_217),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_268),
.C(n_270),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_236),
.B1(n_254),
.B2(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_277),
.B(n_246),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_242),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_242),
.A2(n_230),
.B1(n_212),
.B2(n_181),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_247),
.B1(n_250),
.B2(n_249),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_210),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.C(n_248),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_230),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_177),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_186),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_222),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_248),
.B(n_187),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_284),
.B(n_287),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_215),
.C(n_246),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_220),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_220),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_270),
.C(n_263),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_225),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_252),
.B1(n_227),
.B2(n_231),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_267),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

OAI211xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_262),
.B(n_271),
.C(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_301),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_288),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_296),
.B(n_178),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_266),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_290),
.B(n_292),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_276),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_282),
.C(n_285),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_259),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_312),
.C(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_291),
.B(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_307),
.B(n_299),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_233),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_195),
.B1(n_186),
.B2(n_234),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_10),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_307),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_235),
.B(n_195),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_298),
.C(n_14),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_324),
.Y(n_325)
);

AOI31xp67_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_298),
.A3(n_13),
.B(n_14),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_10),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_312),
.B(n_315),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_319),
.B(n_14),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_325),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_321),
.B(n_13),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.Y(n_334)
);


endmodule