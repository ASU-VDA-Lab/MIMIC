module real_aes_16512_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_725, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_725;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_171;
wire n_87;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_0), .Y(n_173) );
INVx1_ASAP7_75t_L g700 ( .A(n_1), .Y(n_700) );
INVx1_ASAP7_75t_L g580 ( .A(n_2), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_2), .B(n_533), .Y(n_664) );
BUFx3_ASAP7_75t_L g217 ( .A(n_3), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_4), .A2(n_48), .B1(n_641), .B2(n_642), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_4), .A2(n_29), .B1(n_666), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_5), .A2(n_29), .B1(n_641), .B2(n_642), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_5), .A2(n_48), .B1(n_673), .B2(n_676), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_8), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_10), .A2(n_64), .B1(n_131), .B2(n_143), .Y(n_226) );
INVx1_ASAP7_75t_L g597 ( .A(n_11), .Y(n_597) );
INVx1_ASAP7_75t_L g616 ( .A(n_11), .Y(n_616) );
INVx2_ASAP7_75t_L g501 ( .A(n_12), .Y(n_501) );
OAI21x1_ASAP7_75t_L g112 ( .A1(n_13), .A2(n_32), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_14), .B(n_120), .Y(n_119) );
AO32x1_ASAP7_75t_L g223 ( .A1(n_15), .A2(n_111), .A3(n_153), .B1(n_195), .B2(n_224), .Y(n_223) );
AO32x2_ASAP7_75t_L g258 ( .A1(n_15), .A2(n_111), .A3(n_153), .B1(n_195), .B2(n_224), .Y(n_258) );
INVx1_ASAP7_75t_L g555 ( .A(n_16), .Y(n_555) );
INVx1_ASAP7_75t_L g566 ( .A(n_17), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_17), .A2(n_71), .B1(n_599), .B2(n_604), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_18), .A2(n_36), .B1(n_120), .B2(n_129), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_19), .B(n_147), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_20), .A2(n_70), .B1(n_143), .B2(n_148), .Y(n_225) );
BUFx3_ASAP7_75t_L g521 ( .A(n_21), .Y(n_521) );
INVx1_ASAP7_75t_L g569 ( .A(n_22), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_23), .B(n_188), .Y(n_192) );
INVx2_ASAP7_75t_L g503 ( .A(n_24), .Y(n_503) );
INVx1_ASAP7_75t_L g652 ( .A(n_24), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_25), .A2(n_50), .B1(n_148), .B2(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g540 ( .A(n_26), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_27), .A2(n_34), .B1(n_635), .B2(n_639), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_27), .A2(n_58), .B1(n_673), .B2(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g504 ( .A(n_28), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_30), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g704 ( .A(n_31), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_33), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_34), .A2(n_75), .B1(n_666), .B2(n_668), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_35), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_37), .A2(n_57), .B1(n_174), .B2(n_188), .Y(n_202) );
BUFx3_ASAP7_75t_L g518 ( .A(n_38), .Y(n_518) );
BUFx3_ASAP7_75t_L g498 ( .A(n_39), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_40), .A2(n_60), .B1(n_131), .B2(n_143), .Y(n_213) );
AND2x4_ASAP7_75t_L g96 ( .A(n_41), .B(n_97), .Y(n_96) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_41), .Y(n_514) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_43), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_44), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g97 ( .A(n_45), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_46), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_47), .A2(n_171), .B(n_172), .C(n_175), .Y(n_170) );
NAND3xp33_ASAP7_75t_L g151 ( .A(n_49), .B(n_143), .C(n_150), .Y(n_151) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_51), .Y(n_537) );
AND2x2_ASAP7_75t_L g177 ( .A(n_52), .B(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_53), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_54), .A2(n_73), .B1(n_131), .B2(n_174), .Y(n_204) );
INVx2_ASAP7_75t_L g93 ( .A(n_55), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_56), .B(n_125), .Y(n_124) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_58), .A2(n_75), .B1(n_654), .B2(n_656), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_59), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_61), .A2(n_525), .B1(n_693), .B2(n_707), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_61), .Y(n_707) );
INVx1_ASAP7_75t_L g530 ( .A(n_62), .Y(n_530) );
BUFx3_ASAP7_75t_L g533 ( .A(n_63), .Y(n_533) );
INVx1_ASAP7_75t_L g558 ( .A(n_63), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_65), .B(n_150), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_65), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_65), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_66), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_66), .Y(n_522) );
INVx1_ASAP7_75t_L g584 ( .A(n_67), .Y(n_584) );
INVx2_ASAP7_75t_L g633 ( .A(n_67), .Y(n_633) );
INVx1_ASAP7_75t_L g651 ( .A(n_67), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_68), .A2(n_77), .B1(n_129), .B2(n_148), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_69), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g695 ( .A(n_70), .Y(n_695) );
INVx1_ASAP7_75t_L g562 ( .A(n_71), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_72), .B(n_134), .Y(n_197) );
INVx1_ASAP7_75t_L g547 ( .A(n_74), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_76), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_98), .B(n_487), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
INVx4_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_94), .Y(n_83) );
AO21x2_ASAP7_75t_L g722 ( .A1(n_84), .A2(n_712), .B(n_723), .Y(n_722) );
NAND2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_91), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx2_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
INVx1_ASAP7_75t_L g171 ( .A(n_90), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_90), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_91), .A2(n_192), .B(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_91), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_91), .A2(n_92), .B1(n_213), .B2(n_214), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_91), .A2(n_190), .B1(n_238), .B2(n_240), .Y(n_237) );
INVx6_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_92), .A2(n_142), .B(n_144), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_92), .A2(n_121), .B1(n_225), .B2(n_226), .Y(n_224) );
BUFx8_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx2_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
INVx1_ASAP7_75t_L g169 ( .A(n_93), .Y(n_169) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
BUFx10_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
BUFx10_ASAP7_75t_L g132 ( .A(n_96), .Y(n_132) );
INVx1_ASAP7_75t_L g176 ( .A(n_96), .Y(n_176) );
INVx1_ASAP7_75t_L g196 ( .A(n_96), .Y(n_196) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_96), .A2(n_200), .A3(n_237), .B(n_241), .Y(n_236) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_97), .Y(n_512) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_103), .B(n_361), .Y(n_102) );
AND5x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_287), .C(n_307), .D(n_323), .E(n_343), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_247), .Y(n_104) );
OAI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_154), .B(n_218), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g355 ( .A(n_107), .Y(n_355) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g341 ( .A(n_108), .Y(n_341) );
OR2x2_ASAP7_75t_L g378 ( .A(n_108), .B(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g444 ( .A(n_108), .B(n_198), .Y(n_444) );
OR2x2_ASAP7_75t_L g453 ( .A(n_108), .B(n_272), .Y(n_453) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_137), .Y(n_108) );
BUFx2_ASAP7_75t_L g230 ( .A(n_109), .Y(n_230) );
INVx1_ASAP7_75t_L g246 ( .A(n_109), .Y(n_246) );
INVx2_ASAP7_75t_SL g305 ( .A(n_109), .Y(n_305) );
AND2x2_ASAP7_75t_L g326 ( .A(n_109), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g430 ( .A(n_109), .B(n_199), .Y(n_430) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_133), .Y(n_109) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_110), .A2(n_114), .B(n_133), .Y(n_270) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx4_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
INVx2_ASAP7_75t_SL g184 ( .A(n_111), .Y(n_184) );
BUFx3_ASAP7_75t_L g200 ( .A(n_111), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_111), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_111), .B(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
OAI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_123), .B(n_132), .Y(n_114) );
O2A1O1Ixp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_119), .C(n_121), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_120), .A2(n_129), .B1(n_166), .B2(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g239 ( .A(n_120), .Y(n_239) );
BUFx4f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B1(n_128), .B2(n_130), .Y(n_123) );
INVx2_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g175 ( .A(n_127), .Y(n_175) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g194 ( .A(n_131), .Y(n_194) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_132), .A2(n_141), .B(n_146), .Y(n_140) );
AOI31xp67_ASAP7_75t_L g210 ( .A1(n_132), .A2(n_211), .A3(n_212), .B(n_215), .Y(n_210) );
INVx2_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g139 ( .A(n_136), .Y(n_139) );
INVx2_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
AND2x2_ASAP7_75t_L g286 ( .A(n_137), .B(n_270), .Y(n_286) );
AND2x2_ASAP7_75t_L g396 ( .A(n_137), .B(n_254), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_152), .Y(n_137) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_138), .A2(n_140), .B(n_152), .Y(n_233) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_SL g188 ( .A(n_143), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_151), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2x1_ASAP7_75t_L g155 ( .A(n_156), .B(n_180), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_158), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g330 ( .A(n_159), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_160), .Y(n_228) );
AND2x2_ASAP7_75t_L g260 ( .A(n_160), .B(n_236), .Y(n_260) );
INVx1_ASAP7_75t_L g264 ( .A(n_160), .Y(n_264) );
INVx1_ASAP7_75t_L g302 ( .A(n_160), .Y(n_302) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g243 ( .A(n_161), .Y(n_243) );
AOI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_177), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_170), .B(n_176), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_165), .B(n_168), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_167), .A2(n_525), .B1(n_693), .B2(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_167), .Y(n_720) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_SL g203 ( .A(n_169), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g721 ( .A(n_173), .Y(n_721) );
INVx2_ASAP7_75t_L g190 ( .A(n_175), .Y(n_190) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_179), .B(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_198), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_181), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g227 ( .A(n_182), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g256 ( .A(n_182), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g265 ( .A(n_182), .Y(n_265) );
INVx3_ASAP7_75t_L g277 ( .A(n_182), .Y(n_277) );
BUFx2_ASAP7_75t_L g315 ( .A(n_182), .Y(n_315) );
INVxp67_ASAP7_75t_L g335 ( .A(n_182), .Y(n_335) );
AND2x2_ASAP7_75t_L g358 ( .A(n_182), .B(n_258), .Y(n_358) );
INVx1_ASAP7_75t_L g372 ( .A(n_182), .Y(n_372) );
OR2x2_ASAP7_75t_L g393 ( .A(n_182), .B(n_257), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_182), .B(n_236), .Y(n_449) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_197), .Y(n_183) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_191), .B(n_195), .Y(n_185) );
AOI21x1_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_190), .Y(n_186) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_SL g205 ( .A(n_196), .Y(n_205) );
INVx1_ASAP7_75t_L g360 ( .A(n_198), .Y(n_360) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
AND2x2_ASAP7_75t_L g245 ( .A(n_199), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
INVx2_ASAP7_75t_L g291 ( .A(n_199), .Y(n_291) );
AND2x2_ASAP7_75t_L g306 ( .A(n_199), .B(n_254), .Y(n_306) );
INVx1_ASAP7_75t_L g327 ( .A(n_199), .Y(n_327) );
AND2x2_ASAP7_75t_L g385 ( .A(n_199), .B(n_208), .Y(n_385) );
AND2x2_ASAP7_75t_L g395 ( .A(n_199), .B(n_270), .Y(n_395) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .A3(n_205), .B(n_206), .Y(n_199) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g232 ( .A(n_209), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g254 ( .A(n_210), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_217), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_229), .B1(n_234), .B2(n_244), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_219), .A2(n_447), .B1(n_451), .B2(n_452), .Y(n_446) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_227), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_220), .B(n_260), .Y(n_351) );
NAND2xp5_ASAP7_75t_R g370 ( .A(n_220), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g382 ( .A(n_222), .B(n_277), .Y(n_382) );
INVx1_ASAP7_75t_L g450 ( .A(n_222), .Y(n_450) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g278 ( .A(n_223), .B(n_236), .Y(n_278) );
OR2x2_ASAP7_75t_L g319 ( .A(n_223), .B(n_236), .Y(n_319) );
INVx1_ASAP7_75t_L g331 ( .A(n_223), .Y(n_331) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_227), .Y(n_473) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g288 ( .A(n_230), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_230), .B(n_306), .Y(n_322) );
INVx1_ASAP7_75t_L g384 ( .A(n_230), .Y(n_384) );
AND2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_231), .B(n_326), .Y(n_475) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
INVx1_ASAP7_75t_L g368 ( .A(n_232), .Y(n_368) );
OR2x2_ASAP7_75t_L g421 ( .A(n_232), .B(n_290), .Y(n_421) );
INVx2_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_234), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_234), .B(n_335), .Y(n_356) );
INVx1_ASAP7_75t_L g416 ( .A(n_234), .Y(n_416) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_234), .A2(n_388), .A3(n_473), .B(n_474), .Y(n_472) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_243), .Y(n_234) );
AND2x4_ASAP7_75t_L g263 ( .A(n_235), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g338 ( .A(n_235), .B(n_258), .Y(n_338) );
INVx1_ASAP7_75t_L g373 ( .A(n_235), .Y(n_373) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g301 ( .A(n_236), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g281 ( .A(n_243), .Y(n_281) );
INVx1_ASAP7_75t_L g337 ( .A(n_243), .Y(n_337) );
OR2x2_ASAP7_75t_L g411 ( .A(n_243), .B(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_243), .B(n_277), .Y(n_469) );
AND2x4_ASAP7_75t_L g249 ( .A(n_245), .B(n_250), .Y(n_249) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_255), .B1(n_261), .B2(n_266), .C(n_275), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_251), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g390 ( .A(n_251), .B(n_291), .Y(n_390) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g274 ( .A(n_252), .Y(n_274) );
INVx1_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
INVx1_ASAP7_75t_L g342 ( .A(n_253), .Y(n_342) );
AND2x2_ASAP7_75t_L g406 ( .A(n_253), .B(n_327), .Y(n_406) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g269 ( .A(n_254), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
AND2x2_ASAP7_75t_L g311 ( .A(n_256), .B(n_301), .Y(n_311) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g298 ( .A(n_258), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_259), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g294 ( .A(n_260), .Y(n_294) );
AND2x4_ASAP7_75t_L g381 ( .A(n_260), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g460 ( .A(n_260), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_262), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx2_ASAP7_75t_L g401 ( .A(n_263), .Y(n_401) );
INVx1_ASAP7_75t_L g317 ( .A(n_264), .Y(n_317) );
AND2x2_ASAP7_75t_L g300 ( .A(n_265), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g375 ( .A(n_265), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_265), .Y(n_410) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_265), .Y(n_461) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_269), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_269), .B(n_325), .Y(n_456) );
INVx1_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_282), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g426 ( .A(n_277), .B(n_338), .Y(n_426) );
AND2x2_ASAP7_75t_L g279 ( .A(n_278), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g376 ( .A(n_278), .Y(n_376) );
INVx1_ASAP7_75t_L g309 ( .A(n_279), .Y(n_309) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g346 ( .A(n_284), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g403 ( .A(n_284), .B(n_348), .Y(n_403) );
OR2x2_ASAP7_75t_L g485 ( .A(n_285), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI32xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_293), .A3(n_295), .B1(n_299), .B2(n_303), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_289), .A2(n_394), .B1(n_426), .B2(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_290), .B(n_294), .C(n_365), .D(n_366), .Y(n_364) );
INVx2_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g419 ( .A(n_291), .B(n_372), .Y(n_419) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g299 ( .A(n_296), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g479 ( .A(n_298), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_300), .A2(n_406), .B(n_434), .C(n_435), .Y(n_433) );
BUFx2_ASAP7_75t_L g388 ( .A(n_301), .Y(n_388) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_305), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g442 ( .A(n_305), .Y(n_442) );
INVx2_ASAP7_75t_L g379 ( .A(n_306), .Y(n_379) );
AND2x4_ASAP7_75t_L g435 ( .A(n_306), .B(n_347), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_320), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_314), .A2(n_414), .A3(n_416), .B1(n_417), .B2(n_418), .C1(n_420), .C2(n_422), .Y(n_413) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g432 ( .A(n_315), .B(n_319), .Y(n_432) );
INVx1_ASAP7_75t_L g443 ( .A(n_316), .Y(n_443) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g437 ( .A(n_317), .B(n_358), .Y(n_437) );
AND2x2_ASAP7_75t_L g458 ( .A(n_318), .B(n_337), .Y(n_458) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g468 ( .A(n_319), .B(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_332), .B2(n_336), .C1(n_339), .C2(n_725), .Y(n_323) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_324), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g366 ( .A(n_325), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_326), .B(n_396), .Y(n_415) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g400 ( .A(n_335), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_335), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_336), .Y(n_465) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx3_ASAP7_75t_L g412 ( .A(n_338), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_339), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_350), .B(n_352), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_347), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .A3(n_356), .B1(n_357), .B2(n_359), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g455 ( .A(n_354), .B(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g365 ( .A(n_358), .Y(n_365) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_438), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_397), .C(n_424), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .C(n_380), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_366), .B(n_384), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B1(n_374), .B2(n_377), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g486 ( .A(n_385), .Y(n_486) );
OAI21xp33_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_391), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g470 ( .A(n_390), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx2_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g428 ( .A(n_396), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_413), .Y(n_397) );
AOI22xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_402), .B1(n_404), .B2(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_401), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g441 ( .A(n_406), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1p5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND4xp25_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .C(n_433), .D(n_436), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_435), .B(n_437), .Y(n_436) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_454), .C(n_462), .D(n_471), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_444), .B2(n_445), .C(n_446), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g451 ( .A(n_444), .Y(n_451) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g480 ( .A(n_448), .Y(n_480) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g483 ( .A(n_450), .Y(n_483) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_457), .B(n_459), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_466), .C(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI31xp33_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_480), .A3(n_481), .B(n_484), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_515), .B1(n_706), .B2(n_708), .C(n_713), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx12f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx8_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_504), .B(n_505), .C(n_511), .Y(n_492) );
AND2x2_ASAP7_75t_L g718 ( .A(n_493), .B(n_505), .Y(n_718) );
INVx4_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_495), .B(n_506), .C(n_509), .Y(n_505) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g603 ( .A(n_497), .Y(n_603) );
AND2x4_ASAP7_75t_L g644 ( .A(n_497), .B(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g595 ( .A(n_498), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_498), .B(n_597), .Y(n_620) );
INVx2_ASAP7_75t_L g628 ( .A(n_498), .Y(n_628) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
AND2x4_ASAP7_75t_L g608 ( .A(n_500), .B(n_595), .Y(n_608) );
INVx1_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
OR2x6_ASAP7_75t_L g618 ( .A(n_500), .B(n_619), .Y(n_618) );
OR2x4_ASAP7_75t_L g623 ( .A(n_500), .B(n_614), .Y(n_623) );
NAND3x1_ASAP7_75t_L g649 ( .A(n_500), .B(n_650), .C(n_652), .Y(n_649) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g510 ( .A(n_501), .B(n_503), .Y(n_510) );
BUFx3_ASAP7_75t_L g602 ( .A(n_501), .Y(n_602) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_503), .Y(n_587) );
AND3x4_ASAP7_75t_L g631 ( .A(n_503), .B(n_602), .C(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g508 ( .A(n_504), .Y(n_508) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g717 ( .A(n_511), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
BUFx2_ASAP7_75t_L g712 ( .A(n_512), .Y(n_712) );
AND2x2_ASAP7_75t_L g723 ( .A(n_512), .B(n_513), .Y(n_723) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g711 ( .A(n_514), .B(n_712), .Y(n_711) );
XNOR2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_694), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_525), .B1(n_692), .B2(n_693), .Y(n_516) );
CKINVDCx14_ASAP7_75t_R g692 ( .A(n_517), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_520), .B2(n_524), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_518), .Y(n_524) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_521), .Y(n_523) );
INVx1_ASAP7_75t_L g693 ( .A(n_525), .Y(n_693) );
BUFx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
NAND3x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_629), .C(n_658), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_578), .B1(n_585), .B2(n_591), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_546), .C(n_561), .D(n_575), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_540), .B2(n_541), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_530), .A2(n_540), .B1(n_610), .B2(n_617), .Y(n_609) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
OR2x2_ASAP7_75t_L g542 ( .A(n_532), .B(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g567 ( .A(n_532), .B(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g554 ( .A(n_533), .Y(n_554) );
AND2x4_ASAP7_75t_L g572 ( .A(n_533), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g686 ( .A(n_533), .B(n_580), .Y(n_686) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g667 ( .A(n_535), .Y(n_667) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g545 ( .A(n_537), .Y(n_545) );
OR2x2_ASAP7_75t_L g552 ( .A(n_537), .B(n_539), .Y(n_552) );
AND2x2_ASAP7_75t_L g559 ( .A(n_537), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g565 ( .A(n_537), .B(n_539), .Y(n_565) );
INVx1_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_539), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g560 ( .A(n_539), .Y(n_560) );
BUFx2_ASAP7_75t_L g568 ( .A(n_539), .Y(n_568) );
AND2x2_ASAP7_75t_L g671 ( .A(n_539), .B(n_545), .Y(n_671) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_555), .B2(n_556), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_547), .A2(n_555), .B1(n_622), .B2(n_624), .Y(n_621) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x6_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g577 ( .A(n_554), .Y(n_577) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_559), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_566), .B2(n_567), .C1(n_569), .C2(n_570), .Y(n_561) );
BUFx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g576 ( .A(n_564), .B(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g680 ( .A(n_565), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g592 ( .A1(n_569), .A2(n_593), .B(n_598), .C(n_608), .Y(n_592) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g590 ( .A(n_583), .Y(n_590) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g688 ( .A(n_590), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_609), .C(n_621), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g639 ( .A(n_595), .Y(n_639) );
BUFx2_ASAP7_75t_L g657 ( .A(n_595), .Y(n_657) );
INVx1_ASAP7_75t_L g645 ( .A(n_596), .Y(n_645) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g607 ( .A(n_597), .Y(n_607) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x4_ASAP7_75t_L g605 ( .A(n_601), .B(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x4_ASAP7_75t_L g624 ( .A(n_613), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g638 ( .A(n_615), .Y(n_638) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g627 ( .A(n_616), .Y(n_627) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_625), .Y(n_641) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x4_ASAP7_75t_L g637 ( .A(n_628), .B(n_638), .Y(n_637) );
AOI33xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .A3(n_640), .B1(n_646), .B2(n_647), .B3(n_653), .Y(n_629) );
BUFx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g663 ( .A(n_633), .Y(n_663) );
BUFx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx8_ASAP7_75t_L g655 ( .A(n_637), .Y(n_655) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx5_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx8_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI33xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_665), .A3(n_672), .B1(n_681), .B2(n_685), .B3(n_689), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_671), .Y(n_691) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g684 ( .A(n_680), .Y(n_684) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_705), .Y(n_694) );
INVx1_ASAP7_75t_L g705 ( .A(n_695), .Y(n_705) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_703), .B2(n_704), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_709), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_710), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_719), .B1(n_721), .B2(n_722), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x6_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
endmodule