module real_aes_11420_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_571;
wire n_1328;
wire n_549;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_2006;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1994;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1931;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_1969;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g1318 ( .A(n_0), .B(n_1319), .Y(n_1318) );
AO221x1_ASAP7_75t_L g1710 ( .A1(n_0), .A2(n_150), .B1(n_1662), .B2(n_1711), .C(n_1713), .Y(n_1710) );
AOI22xp5_ASAP7_75t_L g1687 ( .A1(n_1), .A2(n_134), .B1(n_1662), .B2(n_1668), .Y(n_1687) );
INVx1_ASAP7_75t_L g1468 ( .A(n_2), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_3), .Y(n_1537) );
CKINVDCx5p33_ASAP7_75t_R g1563 ( .A(n_4), .Y(n_1563) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_5), .A2(n_271), .B1(n_850), .B2(n_917), .C(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1137 ( .A(n_5), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_6), .A2(n_108), .B1(n_465), .B2(n_473), .Y(n_464) );
INVx1_ASAP7_75t_L g566 ( .A(n_6), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_7), .A2(n_333), .B1(n_692), .B2(n_695), .Y(n_1064) );
INVx1_ASAP7_75t_L g1086 ( .A(n_7), .Y(n_1086) );
INVx1_ASAP7_75t_L g1184 ( .A(n_8), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_8), .A2(n_155), .B1(n_1160), .B2(n_1214), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_9), .A2(n_228), .B1(n_916), .B2(n_917), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_9), .A2(n_228), .B1(n_932), .B2(n_934), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g1643 ( .A1(n_10), .A2(n_220), .B1(n_727), .B2(n_728), .C(n_850), .Y(n_1643) );
OAI22xp33_ASAP7_75t_L g1648 ( .A1(n_10), .A2(n_335), .B1(n_695), .B2(n_1367), .Y(n_1648) );
INVx1_ASAP7_75t_L g1953 ( .A(n_11), .Y(n_1953) );
INVx1_ASAP7_75t_L g714 ( .A(n_12), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_12), .A2(n_117), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g1339 ( .A(n_13), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_13), .A2(n_214), .B1(n_622), .B2(n_628), .Y(n_1348) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_14), .A2(n_106), .B1(n_633), .B2(n_635), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_14), .A2(n_106), .B1(n_642), .B2(n_654), .C(n_656), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_15), .A2(n_297), .B1(n_607), .B2(n_610), .C(n_1235), .Y(n_1449) );
OAI22xp33_ASAP7_75t_L g1455 ( .A1(n_15), .A2(n_114), .B1(n_1369), .B2(n_1371), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_16), .A2(n_120), .B1(n_730), .B2(n_732), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_16), .A2(n_120), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g1714 ( .A(n_17), .Y(n_1714) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_18), .A2(n_318), .B1(n_544), .B2(n_610), .C(n_717), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_18), .A2(n_318), .B1(n_747), .B2(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g1059 ( .A(n_19), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_20), .A2(n_75), .B1(n_465), .B2(n_473), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_20), .A2(n_205), .B1(n_390), .B2(n_712), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1584 ( .A(n_21), .Y(n_1584) );
AO22x2_ASAP7_75t_L g894 ( .A1(n_22), .A2(n_895), .B1(n_955), .B2(n_956), .Y(n_894) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_22), .Y(n_955) );
CKINVDCx16_ASAP7_75t_R g1112 ( .A(n_23), .Y(n_1112) );
AOI21xp5_ASAP7_75t_L g1195 ( .A1(n_24), .A2(n_606), .B(n_607), .Y(n_1195) );
INVx1_ASAP7_75t_L g1198 ( .A(n_24), .Y(n_1198) );
XNOR2xp5_ASAP7_75t_L g1566 ( .A(n_25), .B(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1257 ( .A(n_26), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_26), .A2(n_128), .B1(n_816), .B2(n_939), .Y(n_1303) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_27), .A2(n_98), .B1(n_730), .B2(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_27), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_28), .A2(n_374), .B1(n_941), .B2(n_1043), .Y(n_1620) );
INVxp67_ASAP7_75t_SL g1637 ( .A(n_28), .Y(n_1637) );
INVx1_ASAP7_75t_L g1016 ( .A(n_29), .Y(n_1016) );
OAI222xp33_ASAP7_75t_L g1022 ( .A1(n_29), .A2(n_259), .B1(n_348), .B2(n_604), .C1(n_948), .C2(n_1023), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g977 ( .A1(n_30), .A2(n_140), .B1(n_978), .B2(n_979), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_30), .A2(n_140), .B1(n_986), .B2(n_987), .Y(n_985) );
INVx1_ASAP7_75t_L g1127 ( .A(n_31), .Y(n_1127) );
AOI22xp33_ASAP7_75t_SL g1161 ( .A1(n_31), .A2(n_323), .B1(n_937), .B2(n_1036), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_32), .A2(n_76), .B1(n_986), .B2(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1140 ( .A(n_32), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_33), .A2(n_222), .B1(n_847), .B2(n_848), .C(n_850), .Y(n_846) );
INVx1_ASAP7_75t_L g882 ( .A(n_33), .Y(n_882) );
INVx1_ASAP7_75t_L g964 ( .A(n_34), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_34), .A2(n_349), .B1(n_717), .B2(n_727), .Y(n_983) );
INVx1_ASAP7_75t_L g1123 ( .A(n_35), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_35), .A2(n_183), .B1(n_1156), .B2(n_1160), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_36), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g564 ( .A(n_36), .Y(n_564) );
INVx1_ASAP7_75t_L g1514 ( .A(n_37), .Y(n_1514) );
AOI221xp5_ASAP7_75t_L g1544 ( .A1(n_37), .A2(n_170), .B1(n_1545), .B2(n_1546), .C(n_1547), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_38), .A2(n_286), .B1(n_919), .B2(n_920), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_38), .A2(n_286), .B1(n_816), .B2(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g381 ( .A(n_39), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_40), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_41), .A2(n_119), .B1(n_854), .B2(n_858), .Y(n_1124) );
INVx1_ASAP7_75t_L g1150 ( .A(n_41), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_42), .A2(n_121), .B1(n_455), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_42), .A2(n_121), .B1(n_982), .B2(n_986), .Y(n_1031) );
AOI21xp33_ASAP7_75t_L g1181 ( .A1(n_43), .A2(n_544), .B(n_610), .Y(n_1181) );
INVx1_ASAP7_75t_L g1211 ( .A(n_43), .Y(n_1211) );
INVx1_ASAP7_75t_L g1471 ( .A(n_44), .Y(n_1471) );
OAI211xp5_ASAP7_75t_SL g1494 ( .A1(n_44), .A2(n_635), .B(n_1495), .C(n_1500), .Y(n_1494) );
INVx1_ASAP7_75t_L g1977 ( .A(n_45), .Y(n_1977) );
OAI221xp5_ASAP7_75t_L g1994 ( .A1(n_45), .A2(n_633), .B1(n_1493), .B2(n_1995), .C(n_1996), .Y(n_1994) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_46), .A2(n_169), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g883 ( .A(n_46), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1683 ( .A1(n_47), .A2(n_158), .B1(n_1662), .B2(n_1668), .Y(n_1683) );
XOR2xp5_ASAP7_75t_L g1054 ( .A(n_48), .B(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1985 ( .A(n_49), .Y(n_1985) );
OAI22xp5_ASAP7_75t_L g2005 ( .A1(n_49), .A2(n_266), .B1(n_1369), .B2(n_1371), .Y(n_2005) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_50), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_50), .A2(n_195), .B1(n_757), .B2(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_51), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_51), .A2(n_238), .B1(n_727), .B2(n_807), .Y(n_812) );
INVx1_ASAP7_75t_L g1026 ( .A(n_52), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_52), .A2(n_256), .B1(n_941), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_53), .A2(n_159), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_53), .A2(n_159), .B1(n_642), .B2(n_744), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_54), .Y(n_1189) );
INVx1_ASAP7_75t_L g1523 ( .A(n_55), .Y(n_1523) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_55), .A2(n_138), .B1(n_751), .B2(n_939), .Y(n_1561) );
CKINVDCx5p33_ASAP7_75t_R g1268 ( .A(n_56), .Y(n_1268) );
AOI22x1_ASAP7_75t_SL g1006 ( .A1(n_57), .A2(n_1007), .B1(n_1044), .B2(n_1045), .Y(n_1006) );
INVx1_ASAP7_75t_L g1044 ( .A(n_57), .Y(n_1044) );
INVx1_ASAP7_75t_L g1930 ( .A(n_58), .Y(n_1930) );
INVx1_ASAP7_75t_L g1428 ( .A(n_59), .Y(n_1428) );
OAI221xp5_ASAP7_75t_L g1436 ( .A1(n_59), .A2(n_633), .B1(n_868), .B2(n_1437), .C(n_1442), .Y(n_1436) );
AO221x2_ASAP7_75t_L g1810 ( .A1(n_60), .A2(n_305), .B1(n_1711), .B2(n_1811), .C(n_1813), .Y(n_1810) );
OAI22xp33_ASAP7_75t_L g1477 ( .A1(n_61), .A2(n_272), .B1(n_692), .B2(n_695), .Y(n_1477) );
INVx1_ASAP7_75t_L g1498 ( .A(n_61), .Y(n_1498) );
INVx1_ASAP7_75t_L g1075 ( .A(n_62), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_62), .A2(n_257), .B1(n_932), .B2(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1619 ( .A(n_63), .Y(n_1619) );
INVx1_ASAP7_75t_L g1393 ( .A(n_64), .Y(n_1393) );
INVx1_ASAP7_75t_L g972 ( .A(n_65), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_65), .A2(n_202), .B1(n_730), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_66), .A2(n_262), .B1(n_919), .B2(n_920), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_66), .A2(n_262), .B1(n_816), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1602 ( .A(n_67), .Y(n_1602) );
OAI22xp33_ASAP7_75t_L g1608 ( .A1(n_67), .A2(n_141), .B1(n_695), .B2(n_1367), .Y(n_1608) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_68), .A2(n_375), .B1(n_941), .B2(n_1102), .Y(n_1575) );
INVx1_ASAP7_75t_L g1589 ( .A(n_68), .Y(n_1589) );
INVx1_ASAP7_75t_L g1070 ( .A(n_69), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_69), .A2(n_218), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
INVx1_ASAP7_75t_L g593 ( .A(n_70), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_70), .A2(n_281), .B1(n_642), .B2(n_644), .C(n_647), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_71), .B(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_72), .A2(n_327), .B1(n_1662), .B2(n_1668), .Y(n_1661) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_73), .A2(n_217), .B1(n_730), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_73), .A2(n_217), .B1(n_741), .B2(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1686 ( .A1(n_74), .A2(n_354), .B1(n_1670), .B2(n_1676), .Y(n_1686) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_75), .A2(n_153), .B1(n_807), .B2(n_916), .Y(n_1032) );
INVx1_ASAP7_75t_L g1138 ( .A(n_76), .Y(n_1138) );
INVxp33_ASAP7_75t_SL g1912 ( .A(n_77), .Y(n_1912) );
AOI22xp33_ASAP7_75t_L g1941 ( .A1(n_77), .A2(n_367), .B1(n_1942), .B2(n_1944), .Y(n_1941) );
INVx1_ASAP7_75t_L g1066 ( .A(n_78), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_79), .A2(n_162), .B1(n_610), .B2(n_807), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_79), .A2(n_162), .B1(n_939), .B2(n_1038), .Y(n_1037) );
AO22x1_ASAP7_75t_L g1702 ( .A1(n_80), .A2(n_290), .B1(n_1668), .B2(n_1703), .Y(n_1702) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_81), .Y(n_1383) );
INVx1_ASAP7_75t_L g1474 ( .A(n_82), .Y(n_1474) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_82), .A2(n_255), .B1(n_622), .B2(n_628), .Y(n_1482) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_83), .Y(n_1279) );
INVx1_ASAP7_75t_L g777 ( .A(n_84), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_84), .A2(n_185), .B1(n_730), .B2(n_811), .Y(n_810) );
AO22x1_ASAP7_75t_L g1704 ( .A1(n_85), .A2(n_288), .B1(n_1670), .B2(n_1676), .Y(n_1704) );
INVx1_ASAP7_75t_L g1512 ( .A(n_86), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_86), .A2(n_246), .B1(n_937), .B2(n_1550), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_87), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1573 ( .A(n_88), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_89), .A2(n_283), .B1(n_816), .B2(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g950 ( .A(n_89), .Y(n_950) );
INVxp67_ASAP7_75t_SL g1924 ( .A(n_90), .Y(n_1924) );
AOI221xp5_ASAP7_75t_L g1948 ( .A1(n_90), .A2(n_370), .B1(n_1101), .B2(n_1949), .C(n_1950), .Y(n_1948) );
INVx1_ASAP7_75t_L g1386 ( .A(n_91), .Y(n_1386) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_91), .A2(n_633), .B1(n_868), .B2(n_1397), .C(n_1398), .Y(n_1396) );
INVx1_ASAP7_75t_L g904 ( .A(n_92), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_92), .A2(n_215), .B1(n_947), .B2(n_948), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g1614 ( .A(n_93), .Y(n_1614) );
XNOR2x2_ASAP7_75t_L g581 ( .A(n_94), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_95), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_95), .A2(n_287), .B1(n_741), .B2(n_751), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g1519 ( .A1(n_96), .A2(n_127), .B1(n_1242), .B2(n_1247), .C(n_1520), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_96), .A2(n_127), .B1(n_1288), .B2(n_1552), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_97), .Y(n_609) );
INVxp33_ASAP7_75t_L g767 ( .A(n_98), .Y(n_767) );
BUFx2_ASAP7_75t_L g407 ( .A(n_99), .Y(n_407) );
BUFx2_ASAP7_75t_L g505 ( .A(n_99), .Y(n_505) );
INVx1_ASAP7_75t_L g576 ( .A(n_99), .Y(n_576) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_99), .B(n_620), .Y(n_1246) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_100), .A2(n_268), .B1(n_919), .B2(n_982), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_100), .A2(n_268), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1174 ( .A(n_101), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_101), .A2(n_145), .B1(n_942), .B2(n_1036), .Y(n_1218) );
INVx1_ASAP7_75t_L g1974 ( .A(n_102), .Y(n_1974) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_103), .A2(n_111), .B1(n_662), .B2(n_671), .Y(n_1391) );
INVx1_ASAP7_75t_L g1410 ( .A(n_103), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_104), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_105), .A2(n_362), .B1(n_642), .B2(n_744), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_105), .A2(n_362), .B1(n_727), .B2(n_989), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_107), .Y(n_1233) );
INVx1_ASAP7_75t_L g444 ( .A(n_108), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_109), .A2(n_172), .B1(n_760), .B2(n_967), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_109), .A2(n_172), .B1(n_720), .B2(n_1000), .Y(n_999) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_110), .Y(n_591) );
INVx1_ASAP7_75t_L g1409 ( .A(n_111), .Y(n_1409) );
OAI221xp5_ASAP7_75t_L g1913 ( .A1(n_112), .A2(n_204), .B1(n_1242), .B2(n_1520), .C(n_1914), .Y(n_1913) );
OAI22xp5_ASAP7_75t_L g1945 ( .A1(n_112), .A2(n_204), .B1(n_1552), .B2(n_1946), .Y(n_1945) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_113), .A2(n_206), .B1(n_544), .B2(n_715), .C(n_1130), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_113), .A2(n_206), .B1(n_1012), .B2(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1447 ( .A(n_114), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_115), .A2(n_223), .B1(n_727), .B2(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_115), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g2002 ( .A(n_116), .Y(n_2002) );
INVxp33_ASAP7_75t_L g709 ( .A(n_117), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g1068 ( .A1(n_118), .A2(n_633), .B1(n_868), .B2(n_1069), .C(n_1073), .Y(n_1068) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_118), .A2(n_295), .B1(n_939), .B2(n_1038), .Y(n_1104) );
INVx1_ASAP7_75t_L g1149 ( .A(n_119), .Y(n_1149) );
AO221x1_ASAP7_75t_L g1697 ( .A1(n_122), .A2(n_136), .B1(n_1662), .B2(n_1668), .C(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_L g1390 ( .A(n_123), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_123), .A2(n_251), .B1(n_622), .B2(n_628), .Y(n_1395) );
AO221x1_ASAP7_75t_L g1689 ( .A1(n_124), .A2(n_342), .B1(n_1662), .B2(n_1668), .C(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1694 ( .A(n_125), .Y(n_1694) );
AOI22xp33_ASAP7_75t_L g1979 ( .A1(n_126), .A2(n_142), .B1(n_816), .B2(n_937), .Y(n_1979) );
OAI22xp5_ASAP7_75t_L g2000 ( .A1(n_126), .A2(n_142), .B1(n_1092), .B2(n_1093), .Y(n_2000) );
INVx1_ASAP7_75t_L g1264 ( .A(n_128), .Y(n_1264) );
INVx1_ASAP7_75t_L g1470 ( .A(n_129), .Y(n_1470) );
OAI221xp5_ASAP7_75t_L g1483 ( .A1(n_129), .A2(n_633), .B1(n_1484), .B2(n_1487), .C(n_1493), .Y(n_1483) );
XNOR2xp5_ASAP7_75t_L g1373 ( .A(n_130), .B(n_1374), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1581 ( .A1(n_131), .A2(n_216), .B1(n_671), .B2(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1606 ( .A(n_131), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_132), .Y(n_1425) );
INVx1_ASAP7_75t_L g1700 ( .A(n_133), .Y(n_1700) );
OA22x2_ASAP7_75t_L g404 ( .A1(n_134), .A2(n_405), .B1(n_579), .B2(n_580), .Y(n_404) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_134), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g1682 ( .A1(n_135), .A2(n_163), .B1(n_1670), .B2(n_1676), .Y(n_1682) );
AOI22xp5_ASAP7_75t_L g1960 ( .A1(n_135), .A2(n_1961), .B1(n_1966), .B2(n_2006), .Y(n_1960) );
XOR2x2_ASAP7_75t_L g1968 ( .A(n_135), .B(n_1969), .Y(n_1968) );
INVx1_ASAP7_75t_L g1640 ( .A(n_137), .Y(n_1640) );
OAI22xp33_ASAP7_75t_L g1649 ( .A1(n_137), .A2(n_220), .B1(n_1369), .B2(n_1371), .Y(n_1649) );
INVx1_ASAP7_75t_L g1531 ( .A(n_138), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_139), .A2(n_180), .B1(n_934), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g953 ( .A(n_139), .Y(n_953) );
AOI221xp5_ASAP7_75t_L g1603 ( .A1(n_141), .A2(n_324), .B1(n_607), .B2(n_727), .C(n_728), .Y(n_1603) );
INVx1_ASAP7_75t_L g1622 ( .A(n_143), .Y(n_1622) );
OAI221xp5_ASAP7_75t_L g1630 ( .A1(n_143), .A2(n_633), .B1(n_1493), .B2(n_1631), .C(n_1635), .Y(n_1630) );
INVx1_ASAP7_75t_L g1814 ( .A(n_144), .Y(n_1814) );
INVx1_ASAP7_75t_L g1175 ( .A(n_145), .Y(n_1175) );
INVx1_ASAP7_75t_L g1063 ( .A(n_146), .Y(n_1063) );
INVx1_ASAP7_75t_L g795 ( .A(n_147), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_147), .A2(n_334), .B1(n_642), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_148), .A2(n_174), .B1(n_994), .B2(n_995), .Y(n_993) );
INVx1_ASAP7_75t_L g1002 ( .A(n_148), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_149), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_151), .A2(n_311), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_151), .A2(n_311), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_L g1598 ( .A(n_152), .Y(n_1598) );
OAI22xp33_ASAP7_75t_L g1609 ( .A1(n_152), .A2(n_324), .B1(n_1369), .B2(n_1371), .Y(n_1609) );
INVx1_ASAP7_75t_L g1011 ( .A(n_153), .Y(n_1011) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_154), .Y(n_445) );
INVx1_ASAP7_75t_L g1179 ( .A(n_155), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_156), .Y(n_1194) );
INVx1_ASAP7_75t_L g1989 ( .A(n_157), .Y(n_1989) );
OAI22xp5_ASAP7_75t_L g2004 ( .A1(n_157), .A2(n_247), .B1(n_695), .B2(n_1367), .Y(n_2004) );
INVx1_ASAP7_75t_L g1667 ( .A(n_160), .Y(n_1667) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_161), .A2(n_350), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
INVx1_ASAP7_75t_L g1451 ( .A(n_161), .Y(n_1451) );
INVx1_ASAP7_75t_L g1691 ( .A(n_164), .Y(n_1691) );
INVx1_ASAP7_75t_L g790 ( .A(n_165), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_165), .A2(n_213), .B1(n_687), .B2(n_816), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_166), .A2(n_373), .B1(n_1154), .B2(n_1341), .Y(n_1426) );
INVx1_ASAP7_75t_L g1439 ( .A(n_166), .Y(n_1439) );
INVx1_ASAP7_75t_L g1973 ( .A(n_167), .Y(n_1973) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_168), .A2(n_328), .B1(n_844), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_168), .A2(n_328), .B1(n_649), .B2(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g879 ( .A(n_169), .Y(n_879) );
INVx1_ASAP7_75t_L g1516 ( .A(n_170), .Y(n_1516) );
INVx1_ASAP7_75t_L g710 ( .A(n_171), .Y(n_710) );
INVx1_ASAP7_75t_L g1258 ( .A(n_173), .Y(n_1258) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_173), .A2(n_229), .B1(n_649), .B2(n_1299), .C(n_1301), .Y(n_1298) );
INVx1_ASAP7_75t_L g1003 ( .A(n_174), .Y(n_1003) );
INVx1_ASAP7_75t_L g1465 ( .A(n_175), .Y(n_1465) );
INVx1_ASAP7_75t_L g1665 ( .A(n_176), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_176), .B(n_1673), .Y(n_1678) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_177), .A2(n_325), .B1(n_986), .B2(n_1192), .C(n_1193), .Y(n_1191) );
INVx1_ASAP7_75t_L g1201 ( .A(n_177), .Y(n_1201) );
INVx1_ASAP7_75t_L g1429 ( .A(n_178), .Y(n_1429) );
OAI211xp5_ASAP7_75t_SL g1444 ( .A1(n_178), .A2(n_635), .B(n_1445), .C(n_1450), .Y(n_1444) );
INVx1_ASAP7_75t_L g900 ( .A(n_179), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_179), .A2(n_208), .B1(n_924), .B2(n_927), .Y(n_923) );
INVx1_ASAP7_75t_L g945 ( .A(n_180), .Y(n_945) );
INVx1_ASAP7_75t_L g1237 ( .A(n_181), .Y(n_1237) );
AOI21xp33_ASAP7_75t_L g1294 ( .A1(n_181), .A2(n_1295), .B(n_1296), .Y(n_1294) );
INVx2_ASAP7_75t_L g393 ( .A(n_182), .Y(n_393) );
INVx1_ASAP7_75t_L g1132 ( .A(n_183), .Y(n_1132) );
INVx1_ASAP7_75t_L g1239 ( .A(n_184), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_184), .A2(n_250), .B1(n_817), .B2(n_1154), .Y(n_1293) );
INVx1_ASAP7_75t_L g780 ( .A(n_185), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g1626 ( .A1(n_186), .A2(n_226), .B1(n_1433), .B2(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1645 ( .A(n_186), .Y(n_1645) );
AOI22xp5_ASAP7_75t_L g1900 ( .A1(n_187), .A2(n_1901), .B1(n_1902), .B2(n_1954), .Y(n_1900) );
CKINVDCx5p33_ASAP7_75t_R g1954 ( .A(n_187), .Y(n_1954) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_188), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_189), .A2(n_369), .B1(n_816), .B2(n_1580), .Y(n_1579) );
OAI22xp5_ASAP7_75t_L g1586 ( .A1(n_189), .A2(n_369), .B1(n_1092), .B2(n_1093), .Y(n_1586) );
INVx1_ASAP7_75t_L g463 ( .A(n_190), .Y(n_463) );
BUFx3_ASAP7_75t_L g479 ( .A(n_190), .Y(n_479) );
INVx1_ASAP7_75t_L g1448 ( .A(n_191), .Y(n_1448) );
OAI22xp33_ASAP7_75t_L g1454 ( .A1(n_191), .A2(n_297), .B1(n_695), .B2(n_1367), .Y(n_1454) );
INVx1_ASAP7_75t_L g863 ( .A(n_192), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_192), .A2(n_291), .B1(n_675), .B2(n_680), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_193), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g1344 ( .A1(n_194), .A2(n_347), .B1(n_662), .B2(n_671), .Y(n_1344) );
INVx1_ASAP7_75t_L g1362 ( .A(n_194), .Y(n_1362) );
INVx1_ASAP7_75t_L g721 ( .A(n_195), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_196), .Y(n_452) );
INVxp33_ASAP7_75t_SL g1909 ( .A(n_197), .Y(n_1909) );
AOI221xp5_ASAP7_75t_L g1937 ( .A1(n_197), .A2(n_319), .B1(n_939), .B2(n_1299), .C(n_1938), .Y(n_1937) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_198), .A2(n_361), .B1(n_606), .B2(n_607), .C(n_1235), .Y(n_1360) );
OAI22xp33_ASAP7_75t_L g1368 ( .A1(n_198), .A2(n_221), .B1(n_1369), .B2(n_1371), .Y(n_1368) );
INVx1_ASAP7_75t_L g1404 ( .A(n_199), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g1413 ( .A1(n_199), .A2(n_201), .B1(n_1369), .B2(n_1371), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_200), .A2(n_341), .B1(n_622), .B2(n_628), .Y(n_621) );
INVx1_ASAP7_75t_L g660 ( .A(n_200), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g1407 ( .A1(n_201), .A2(n_240), .B1(n_606), .B2(n_607), .C(n_717), .Y(n_1407) );
INVx1_ASAP7_75t_L g973 ( .A(n_202), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_203), .A2(n_280), .B1(n_760), .B2(n_782), .C(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g793 ( .A(n_203), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_205), .A2(n_259), .B1(n_1040), .B2(n_1041), .Y(n_1039) );
INVx1_ASAP7_75t_L g1623 ( .A(n_207), .Y(n_1623) );
OAI211xp5_ASAP7_75t_SL g1638 ( .A1(n_207), .A2(n_635), .B(n_1639), .C(n_1644), .Y(n_1638) );
INVx1_ASAP7_75t_L g910 ( .A(n_208), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_209), .Y(n_1539) );
AOI22xp5_ASAP7_75t_L g1669 ( .A1(n_210), .A2(n_242), .B1(n_1670), .B2(n_1676), .Y(n_1669) );
AOI22xp33_ASAP7_75t_L g1975 ( .A1(n_211), .A2(n_351), .B1(n_941), .B2(n_1043), .Y(n_1975) );
INVxp67_ASAP7_75t_SL g1999 ( .A(n_211), .Y(n_1999) );
INVx1_ASAP7_75t_L g1715 ( .A(n_212), .Y(n_1715) );
INVx1_ASAP7_75t_L g791 ( .A(n_213), .Y(n_791) );
INVx1_ASAP7_75t_L g1342 ( .A(n_214), .Y(n_1342) );
INVx1_ASAP7_75t_L g907 ( .A(n_215), .Y(n_907) );
INVx1_ASAP7_75t_L g1605 ( .A(n_216), .Y(n_1605) );
INVx1_ASAP7_75t_L g1072 ( .A(n_218), .Y(n_1072) );
INVx1_ASAP7_75t_L g1816 ( .A(n_219), .Y(n_1816) );
INVx1_ASAP7_75t_L g1357 ( .A(n_221), .Y(n_1357) );
INVx1_ASAP7_75t_L g880 ( .A(n_222), .Y(n_880) );
INVxp33_ASAP7_75t_L g762 ( .A(n_223), .Y(n_762) );
INVx1_ASAP7_75t_L g503 ( .A(n_224), .Y(n_503) );
INVx1_ASAP7_75t_L g669 ( .A(n_224), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g1478 ( .A1(n_225), .A2(n_303), .B1(n_1369), .B2(n_1371), .Y(n_1478) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_225), .A2(n_272), .B1(n_607), .B2(n_1122), .C(n_1235), .Y(n_1499) );
INVx1_ASAP7_75t_L g1646 ( .A(n_226), .Y(n_1646) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_227), .Y(n_522) );
INVx1_ASAP7_75t_L g1260 ( .A(n_229), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1536 ( .A(n_230), .Y(n_1536) );
INVx1_ASAP7_75t_L g860 ( .A(n_231), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_231), .A2(n_284), .B1(n_649), .B2(n_817), .Y(n_877) );
INVx1_ASAP7_75t_L g1932 ( .A(n_232), .Y(n_1932) );
CKINVDCx5p33_ASAP7_75t_R g1540 ( .A(n_233), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_234), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_235), .Y(n_899) );
INVx1_ASAP7_75t_L g1699 ( .A(n_236), .Y(n_1699) );
XOR2xp5_ASAP7_75t_L g1507 ( .A(n_237), .B(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g784 ( .A(n_238), .Y(n_784) );
INVxp67_ASAP7_75t_SL g1925 ( .A(n_239), .Y(n_1925) );
AOI22xp33_ASAP7_75t_L g1951 ( .A1(n_239), .A2(n_320), .B1(n_1040), .B2(n_1043), .Y(n_1951) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_240), .A2(n_338), .B1(n_695), .B2(n_1367), .Y(n_1412) );
INVx1_ASAP7_75t_L g1525 ( .A(n_241), .Y(n_1525) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_241), .A2(n_260), .B1(n_1556), .B2(n_1557), .C(n_1558), .Y(n_1555) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_243), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_244), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_244), .A2(n_662), .B1(n_670), .B2(n_671), .C(n_674), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g1266 ( .A(n_245), .Y(n_1266) );
INVx1_ASAP7_75t_L g1517 ( .A(n_246), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g1990 ( .A1(n_247), .A2(n_266), .B1(n_607), .B2(n_727), .C(n_736), .Y(n_1990) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_248), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_249), .A2(n_275), .B1(n_854), .B2(n_858), .Y(n_853) );
INVx1_ASAP7_75t_L g888 ( .A(n_249), .Y(n_888) );
INVx1_ASAP7_75t_L g1229 ( .A(n_250), .Y(n_1229) );
INVx1_ASAP7_75t_L g1389 ( .A(n_251), .Y(n_1389) );
INVx1_ASAP7_75t_L g1062 ( .A(n_252), .Y(n_1062) );
INVx1_ASAP7_75t_L g892 ( .A(n_253), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g1467 ( .A(n_254), .Y(n_1467) );
INVx1_ASAP7_75t_L g1473 ( .A(n_255), .Y(n_1473) );
INVx1_ASAP7_75t_L g1027 ( .A(n_256), .Y(n_1027) );
INVx1_ASAP7_75t_L g1074 ( .A(n_257), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g1325 ( .A(n_258), .Y(n_1325) );
INVx1_ASAP7_75t_L g1528 ( .A(n_260), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_261), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_263), .Y(n_1187) );
INVx1_ASAP7_75t_L g1578 ( .A(n_264), .Y(n_1578) );
OAI211xp5_ASAP7_75t_SL g1595 ( .A1(n_264), .A2(n_635), .B(n_1596), .C(n_1604), .Y(n_1595) );
CKINVDCx16_ASAP7_75t_R g698 ( .A(n_265), .Y(n_698) );
INVx1_ASAP7_75t_L g1334 ( .A(n_267), .Y(n_1334) );
OAI221xp5_ASAP7_75t_L g1349 ( .A1(n_267), .A2(n_633), .B1(n_868), .B2(n_1350), .C(n_1351), .Y(n_1349) );
INVx1_ASAP7_75t_L g1418 ( .A(n_269), .Y(n_1418) );
INVx1_ASAP7_75t_L g1577 ( .A(n_270), .Y(n_1577) );
OAI221xp5_ASAP7_75t_L g1587 ( .A1(n_270), .A2(n_633), .B1(n_868), .B2(n_1588), .C(n_1594), .Y(n_1587) );
INVx1_ASAP7_75t_L g1141 ( .A(n_271), .Y(n_1141) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_273), .Y(n_1329) );
INVx1_ASAP7_75t_L g1463 ( .A(n_274), .Y(n_1463) );
INVx1_ASAP7_75t_L g886 ( .A(n_275), .Y(n_886) );
INVx1_ASAP7_75t_L g909 ( .A(n_276), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_276), .A2(n_363), .B1(n_916), .B2(n_917), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_277), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_278), .A2(n_300), .B1(n_412), .B2(n_420), .Y(n_411) );
INVx1_ASAP7_75t_L g536 ( .A(n_278), .Y(n_536) );
INVx1_ASAP7_75t_L g1423 ( .A(n_279), .Y(n_1423) );
AOI21xp33_ASAP7_75t_L g1443 ( .A1(n_279), .A2(n_544), .B(n_1122), .Y(n_1443) );
INVx1_ASAP7_75t_L g794 ( .A(n_280), .Y(n_794) );
AOI21xp33_ASAP7_75t_L g595 ( .A1(n_281), .A2(n_544), .B(n_596), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g1572 ( .A(n_282), .Y(n_1572) );
INVx1_ASAP7_75t_L g951 ( .A(n_283), .Y(n_951) );
INVx1_ASAP7_75t_L g861 ( .A(n_284), .Y(n_861) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_285), .A2(n_427), .B(n_432), .C(n_439), .Y(n_426) );
INVx1_ASAP7_75t_L g532 ( .A(n_285), .Y(n_532) );
INVx1_ASAP7_75t_L g704 ( .A(n_287), .Y(n_704) );
INVx1_ASAP7_75t_L g1978 ( .A(n_289), .Y(n_1978) );
OAI211xp5_ASAP7_75t_SL g1982 ( .A1(n_289), .A2(n_635), .B(n_1983), .C(n_1991), .Y(n_1982) );
XNOR2xp5_ASAP7_75t_L g1415 ( .A(n_290), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g852 ( .A(n_291), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g1430 ( .A1(n_292), .A2(n_315), .B1(n_751), .B2(n_1324), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_292), .A2(n_315), .B1(n_1092), .B2(n_1093), .Y(n_1435) );
BUFx3_ASAP7_75t_L g462 ( .A(n_293), .Y(n_462) );
INVx1_ASAP7_75t_L g472 ( .A(n_293), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_294), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_295), .A2(n_635), .B1(n_1078), .B2(n_1081), .C(n_1087), .Y(n_1077) );
INVx1_ASAP7_75t_L g1480 ( .A(n_296), .Y(n_1480) );
INVx1_ASAP7_75t_L g1336 ( .A(n_298), .Y(n_1336) );
OAI211xp5_ASAP7_75t_L g1354 ( .A1(n_298), .A2(n_635), .B(n_1355), .C(n_1361), .Y(n_1354) );
AO22x2_ASAP7_75t_L g771 ( .A1(n_299), .A2(n_772), .B1(n_826), .B2(n_827), .Y(n_771) );
INVxp67_ASAP7_75t_L g826 ( .A(n_299), .Y(n_826) );
INVx1_ASAP7_75t_L g534 ( .A(n_300), .Y(n_534) );
XNOR2xp5_ASAP7_75t_L g1457 ( .A(n_301), .B(n_1458), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_302), .Y(n_389) );
INVx1_ASAP7_75t_L g578 ( .A(n_302), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_302), .B(n_353), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_302), .B(n_416), .Y(n_624) );
INVx1_ASAP7_75t_L g1497 ( .A(n_303), .Y(n_1497) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_304), .A2(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g685 ( .A(n_304), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g960 ( .A(n_306), .B(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g459 ( .A(n_307), .Y(n_459) );
OR2x2_ASAP7_75t_L g684 ( .A(n_307), .B(n_669), .Y(n_684) );
INVx1_ASAP7_75t_L g1359 ( .A(n_308), .Y(n_1359) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_308), .A2(n_361), .B1(n_695), .B2(n_1367), .Y(n_1366) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_309), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_310), .Y(n_513) );
INVx1_ASAP7_75t_L g1346 ( .A(n_312), .Y(n_1346) );
INVx1_ASAP7_75t_L g1387 ( .A(n_313), .Y(n_1387) );
OAI211xp5_ASAP7_75t_L g1402 ( .A1(n_313), .A2(n_635), .B(n_1403), .C(n_1408), .Y(n_1402) );
INVx1_ASAP7_75t_L g1927 ( .A(n_314), .Y(n_1927) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_316), .Y(n_599) );
INVx1_ASAP7_75t_L g1224 ( .A(n_317), .Y(n_1224) );
INVxp33_ASAP7_75t_L g1911 ( .A(n_319), .Y(n_1911) );
INVxp33_ASAP7_75t_L g1917 ( .A(n_320), .Y(n_1917) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_321), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_322), .A2(n_340), .B1(n_642), .B2(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g1005 ( .A(n_322), .Y(n_1005) );
INVx1_ASAP7_75t_L g1126 ( .A(n_323), .Y(n_1126) );
INVx1_ASAP7_75t_L g1199 ( .A(n_325), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1624 ( .A1(n_326), .A2(n_355), .B1(n_1107), .B2(n_1625), .Y(n_1624) );
OAI22xp5_ASAP7_75t_L g1629 ( .A1(n_326), .A2(n_355), .B1(n_622), .B2(n_628), .Y(n_1629) );
INVx1_ASAP7_75t_L g1611 ( .A(n_327), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_329), .A2(n_371), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_329), .A2(n_371), .B1(n_484), .B2(n_744), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g1980 ( .A1(n_330), .A2(n_366), .B1(n_671), .B2(n_1582), .Y(n_1980) );
INVx1_ASAP7_75t_L g1993 ( .A(n_330), .Y(n_1993) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_331), .Y(n_1271) );
CKINVDCx5p33_ASAP7_75t_R g1379 ( .A(n_332), .Y(n_1379) );
INVx1_ASAP7_75t_L g1079 ( .A(n_333), .Y(n_1079) );
INVx1_ASAP7_75t_L g800 ( .A(n_334), .Y(n_800) );
INVx1_ASAP7_75t_L g1642 ( .A(n_335), .Y(n_1642) );
INVx1_ASAP7_75t_L g1060 ( .A(n_336), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1475 ( .A1(n_337), .A2(n_360), .B1(n_1432), .B2(n_1433), .Y(n_1475) );
INVx1_ASAP7_75t_L g1502 ( .A(n_337), .Y(n_1502) );
INVx1_ASAP7_75t_L g1406 ( .A(n_338), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_339), .Y(n_1380) );
INVx1_ASAP7_75t_L g998 ( .A(n_340), .Y(n_998) );
INVx1_ASAP7_75t_L g657 ( .A(n_341), .Y(n_657) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
AND3x2_ASAP7_75t_L g1666 ( .A(n_343), .B(n_381), .C(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_343), .B(n_381), .Y(n_1675) );
INVx2_ASAP7_75t_L g394 ( .A(n_344), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g1327 ( .A(n_345), .Y(n_1327) );
INVx1_ASAP7_75t_L g1382 ( .A(n_346), .Y(n_1382) );
AOI21xp33_ASAP7_75t_L g1400 ( .A1(n_346), .A2(n_544), .B(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1364 ( .A(n_347), .Y(n_1364) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_348), .Y(n_1015) );
INVx1_ASAP7_75t_L g969 ( .A(n_349), .Y(n_969) );
INVx1_ASAP7_75t_L g1452 ( .A(n_350), .Y(n_1452) );
INVxp67_ASAP7_75t_SL g1997 ( .A(n_351), .Y(n_1997) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_352), .A2(n_356), .B1(n_1242), .B2(n_1247), .C(n_1249), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1284 ( .A1(n_352), .A2(n_356), .B1(n_1285), .B2(n_1288), .C(n_1290), .Y(n_1284) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
INVx2_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
AO22x2_ASAP7_75t_L g1165 ( .A1(n_357), .A2(n_1166), .B1(n_1220), .B2(n_1221), .Y(n_1165) );
INVxp67_ASAP7_75t_SL g1220 ( .A(n_357), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_358), .Y(n_410) );
INVx1_ASAP7_75t_L g1933 ( .A(n_359), .Y(n_1933) );
INVx1_ASAP7_75t_L g1501 ( .A(n_360), .Y(n_1501) );
INVx1_ASAP7_75t_L g902 ( .A(n_363), .Y(n_902) );
INVx1_ASAP7_75t_L g613 ( .A(n_364), .Y(n_613) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_364), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_365), .A2(n_482), .B(n_487), .C(n_498), .Y(n_481) );
INVx1_ASAP7_75t_L g571 ( .A(n_365), .Y(n_571) );
INVx1_ASAP7_75t_L g1992 ( .A(n_366), .Y(n_1992) );
INVxp33_ASAP7_75t_SL g1907 ( .A(n_367), .Y(n_1907) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_368), .B(n_1143), .Y(n_1142) );
INVxp33_ASAP7_75t_SL g1921 ( .A(n_370), .Y(n_1921) );
INVx1_ASAP7_75t_L g1618 ( .A(n_372), .Y(n_1618) );
INVx1_ASAP7_75t_L g1441 ( .A(n_373), .Y(n_1441) );
INVxp33_ASAP7_75t_SL g1636 ( .A(n_374), .Y(n_1636) );
INVx1_ASAP7_75t_L g1593 ( .A(n_375), .Y(n_1593) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_397), .B(n_1653), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1965 ( .A(n_379), .B(n_385), .Y(n_1965) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1959 ( .A(n_380), .Y(n_1959) );
NAND2xp5_ASAP7_75t_L g2008 ( .A(n_380), .B(n_382), .Y(n_2008) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1958 ( .A(n_382), .B(n_1959), .Y(n_1958) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g406 ( .A(n_387), .B(n_407), .Y(n_406) );
OR2x6_ASAP7_75t_L g701 ( .A(n_387), .B(n_407), .Y(n_701) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g725 ( .A(n_388), .B(n_396), .Y(n_725) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g544 ( .A(n_389), .B(n_415), .Y(n_544) );
INVx8_ASAP7_75t_L g409 ( .A(n_390), .Y(n_409) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_391), .Y(n_546) );
OR2x6_ASAP7_75t_L g712 ( .A(n_391), .B(n_414), .Y(n_712) );
INVx2_ASAP7_75t_SL g1256 ( .A(n_391), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_391), .B(n_1246), .Y(n_1277) );
INVx1_ASAP7_75t_L g1353 ( .A(n_391), .Y(n_1353) );
BUFx2_ASAP7_75t_L g1490 ( .A(n_391), .Y(n_1490) );
INVx2_ASAP7_75t_SL g1920 ( .A(n_391), .Y(n_1920) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_L g419 ( .A(n_393), .Y(n_419) );
AND2x4_ASAP7_75t_L g424 ( .A(n_393), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_393), .B(n_394), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_394), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
INVx1_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g627 ( .A(n_394), .Y(n_627) );
AND2x4_ASAP7_75t_L g446 ( .A(n_395), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g948 ( .A(n_396), .B(n_450), .Y(n_948) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_396), .B(n_450), .Y(n_1000) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_1047), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_829), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_696), .Y(n_402) );
XNOR2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_581), .Y(n_403) );
INVx1_ASAP7_75t_L g579 ( .A(n_405), .Y(n_579) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_453), .C(n_506), .Y(n_405) );
AOI31xp33_ASAP7_75t_L g943 ( .A1(n_406), .A2(n_944), .A3(n_949), .B(n_952), .Y(n_943) );
AND2x4_ASAP7_75t_L g539 ( .A(n_407), .B(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g688 ( .A(n_407), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g752 ( .A(n_407), .B(n_540), .Y(n_752) );
AOI211xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_411), .C(n_426), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_409), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_409), .A2(n_711), .B1(n_779), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_409), .A2(n_899), .B1(n_953), .B2(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_409), .A2(n_954), .B1(n_970), .B2(n_1005), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_410), .A2(n_523), .B1(n_530), .B2(n_532), .Y(n_529) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_417), .Y(n_412) );
AOI322xp5_ASAP7_75t_L g439 ( .A1(n_413), .A2(n_440), .A3(n_444), .B1(n_445), .B2(n_446), .C1(n_448), .C2(n_452), .Y(n_439) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g421 ( .A(n_414), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g705 ( .A(n_414), .B(n_625), .Y(n_705) );
AND2x4_ASAP7_75t_L g707 ( .A(n_414), .B(n_422), .Y(n_707) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g436 ( .A(n_416), .Y(n_436) );
INVx2_ASAP7_75t_L g552 ( .A(n_417), .Y(n_552) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_417), .Y(n_1183) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g559 ( .A(n_418), .Y(n_559) );
INVx1_ASAP7_75t_L g587 ( .A(n_418), .Y(n_587) );
INVx1_ASAP7_75t_L g616 ( .A(n_419), .Y(n_616) );
AND2x4_ASAP7_75t_L g625 ( .A(n_419), .B(n_626), .Y(n_625) );
INVx5_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_421), .A2(n_705), .B1(n_950), .B2(n_951), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_421), .A2(n_705), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_421), .A2(n_705), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g1534 ( .A(n_423), .Y(n_1534) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g555 ( .A(n_424), .Y(n_555) );
INVx3_ASAP7_75t_L g563 ( .A(n_424), .Y(n_563) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_424), .Y(n_922) );
AND2x4_ASAP7_75t_L g437 ( .A(n_425), .B(n_438), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g1254 ( .A1(n_427), .A2(n_1255), .B1(n_1257), .B2(n_1258), .Y(n_1254) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_427), .A2(n_1270), .B1(n_1271), .B2(n_1272), .Y(n_1269) );
OAI221xp5_ASAP7_75t_L g1995 ( .A1(n_427), .A2(n_1076), .B1(n_1919), .B2(n_1973), .C(n_1974), .Y(n_1995) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g1632 ( .A(n_428), .Y(n_1632) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g549 ( .A(n_429), .Y(n_549) );
INVx3_ASAP7_75t_L g594 ( .A(n_429), .Y(n_594) );
INVx2_ASAP7_75t_L g604 ( .A(n_429), .Y(n_604) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_430), .B(n_431), .Y(n_570) );
INVx1_ASAP7_75t_L g450 ( .A(n_431), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_432), .B(n_703), .C(n_708), .D(n_713), .Y(n_702) );
NAND4xp25_ASAP7_75t_SL g788 ( .A(n_432), .B(n_789), .C(n_792), .D(n_799), .Y(n_788) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
AOI211xp5_ASAP7_75t_L g944 ( .A1(n_433), .A2(n_848), .B(n_945), .C(n_946), .Y(n_944) );
AOI211xp5_ASAP7_75t_L g997 ( .A1(n_433), .A2(n_917), .B(n_998), .C(n_999), .Y(n_997) );
NOR3xp33_ASAP7_75t_L g1021 ( .A(n_433), .B(n_1022), .C(n_1024), .Y(n_1021) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_436), .B(n_578), .Y(n_577) );
BUFx3_ASAP7_75t_L g637 ( .A(n_437), .Y(n_637) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_437), .Y(n_717) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_437), .Y(n_737) );
BUFx2_ASAP7_75t_L g798 ( .A(n_437), .Y(n_798) );
BUFx3_ASAP7_75t_L g1235 ( .A(n_437), .Y(n_1235) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g806 ( .A(n_441), .Y(n_806) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_441), .Y(n_1401) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_442), .Y(n_610) );
AND2x4_ASAP7_75t_L g634 ( .A(n_442), .B(n_624), .Y(n_634) );
BUFx2_ASAP7_75t_L g847 ( .A(n_442), .Y(n_847) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g597 ( .A(n_443), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g487 ( .A1(n_445), .A2(n_452), .A3(n_488), .B1(n_490), .B2(n_491), .C1(n_492), .C2(n_496), .Y(n_487) );
INVx2_ASAP7_75t_L g720 ( .A(n_446), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g792 ( .A1(n_446), .A2(n_448), .B1(n_793), .B2(n_794), .C1(n_795), .C2(n_796), .Y(n_792) );
INVx2_ASAP7_75t_L g947 ( .A(n_446), .Y(n_947) );
INVx2_ASAP7_75t_L g1023 ( .A(n_446), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_447), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g856 ( .A(n_447), .Y(n_856) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_447), .Y(n_1089) );
AOI222xp33_ASAP7_75t_L g713 ( .A1(n_448), .A2(n_714), .B1(n_715), .B2(n_718), .C1(n_719), .C2(n_721), .Y(n_713) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI31xp33_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_464), .A3(n_481), .B(n_501), .Y(n_453) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_456), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_456), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_456), .A2(n_474), .B1(n_899), .B2(n_900), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_456), .A2(n_766), .B1(n_972), .B2(n_973), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_456), .A2(n_474), .B1(n_1169), .B2(n_1201), .Y(n_1200) );
AND2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .Y(n_456) );
AND2x4_ASAP7_75t_L g763 ( .A(n_457), .B(n_764), .Y(n_763) );
AND2x4_ASAP7_75t_L g775 ( .A(n_457), .B(n_764), .Y(n_775) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g758 ( .A(n_458), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g468 ( .A(n_459), .Y(n_468) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_459), .Y(n_476) );
AND2x2_ASAP7_75t_L g510 ( .A(n_459), .B(n_503), .Y(n_510) );
INVx2_ASAP7_75t_L g541 ( .A(n_459), .Y(n_541) );
INVx1_ASAP7_75t_L g537 ( .A(n_460), .Y(n_537) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_460), .Y(n_742) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_460), .Y(n_751) );
INVx2_ASAP7_75t_L g1108 ( .A(n_460), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g1341 ( .A(n_460), .Y(n_1341) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
INVx1_ASAP7_75t_L g650 ( .A(n_461), .Y(n_650) );
INVx1_ASAP7_75t_L g693 ( .A(n_461), .Y(n_693) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_461), .Y(n_817) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g480 ( .A(n_462), .Y(n_480) );
AND2x2_ASAP7_75t_L g486 ( .A(n_462), .B(n_479), .Y(n_486) );
INVx1_ASAP7_75t_L g470 ( .A(n_463), .Y(n_470) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
INVx1_ASAP7_75t_L g490 ( .A(n_466), .Y(n_490) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g483 ( .A(n_467), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
AND2x6_ASAP7_75t_L g766 ( .A(n_467), .B(n_489), .Y(n_766) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g496 ( .A(n_468), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g524 ( .A(n_469), .Y(n_524) );
INVx1_ASAP7_75t_L g1210 ( .A(n_469), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_469), .B(n_684), .Y(n_1311) );
BUFx2_ASAP7_75t_L g1422 ( .A(n_469), .Y(n_1422) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g528 ( .A(n_470), .B(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g489 ( .A(n_472), .B(n_479), .Y(n_489) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_474), .A2(n_710), .B1(n_762), .B2(n_763), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_474), .A2(n_766), .B1(n_779), .B2(n_780), .C(n_781), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_474), .A2(n_775), .B1(n_969), .B2(n_970), .Y(n_968) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_475), .B(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g906 ( .A(n_475), .B(n_493), .Y(n_906) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx6_ASAP7_75t_L g646 ( .A(n_477), .Y(n_646) );
INVx2_ASAP7_75t_L g681 ( .A(n_477), .Y(n_681) );
AND2x2_ASAP7_75t_L g689 ( .A(n_477), .B(n_667), .Y(n_689) );
BUFx2_ASAP7_75t_L g747 ( .A(n_477), .Y(n_747) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g497 ( .A(n_478), .Y(n_497) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g495 ( .A(n_480), .Y(n_495) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g754 ( .A1(n_483), .A2(n_499), .B(n_755), .C(n_756), .Y(n_754) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_484), .Y(n_903) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_484), .Y(n_965) );
HB1xp67_ASAP7_75t_L g1546 ( .A(n_484), .Y(n_1546) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g499 ( .A(n_485), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g643 ( .A(n_485), .Y(n_643) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_485), .Y(n_785) );
INVx1_ASAP7_75t_L g891 ( .A(n_485), .Y(n_891) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_486), .Y(n_676) );
INVx2_ASAP7_75t_L g516 ( .A(n_488), .Y(n_516) );
INVx1_ASAP7_75t_L g1338 ( .A(n_488), .Y(n_1338) );
INVx2_ASAP7_75t_SL g1378 ( .A(n_488), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g535 ( .A(n_489), .Y(n_535) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_489), .Y(n_649) );
BUFx2_ASAP7_75t_L g741 ( .A(n_489), .Y(n_741) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_489), .Y(n_942) );
BUFx6f_ASAP7_75t_L g1154 ( .A(n_489), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1324 ( .A(n_489), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_491), .A2(n_557), .B1(n_560), .B2(n_564), .Y(n_556) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g759 ( .A(n_494), .Y(n_759) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g664 ( .A(n_495), .Y(n_664) );
INVx3_ASAP7_75t_L g760 ( .A(n_496), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_496), .A2(n_902), .B1(n_903), .B2(n_904), .C1(n_905), .C2(n_907), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_496), .A2(n_906), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI222xp33_ASAP7_75t_L g1202 ( .A1(n_496), .A2(n_905), .B1(n_1189), .B2(n_1190), .C1(n_1194), .C2(n_1203), .Y(n_1202) );
BUFx3_ASAP7_75t_L g673 ( .A(n_497), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_498), .B(n_1010), .C(n_1014), .Y(n_1009) );
CKINVDCx8_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g897 ( .A(n_499), .Y(n_897) );
AOI211xp5_ASAP7_75t_L g963 ( .A1(n_499), .A2(n_964), .B(n_965), .C(n_966), .Y(n_963) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_500), .A2(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_SL g769 ( .A(n_501), .Y(n_769) );
OAI31xp33_ASAP7_75t_L g1008 ( .A1(n_501), .A2(n_1009), .A3(n_1017), .B(n_1019), .Y(n_1008) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
AND2x4_ASAP7_75t_L g787 ( .A(n_502), .B(n_504), .Y(n_787) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g540 ( .A(n_503), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g1095 ( .A(n_504), .Y(n_1095) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g511 ( .A(n_505), .Y(n_511) );
OR2x6_ASAP7_75t_L g543 ( .A(n_505), .B(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_542), .Y(n_506) );
OAI33xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_512), .A3(n_521), .B1(n_529), .B2(n_533), .B3(n_538), .Y(n_507) );
INVx1_ASAP7_75t_SL g739 ( .A(n_508), .Y(n_739) );
OAI33xp33_ASAP7_75t_L g1321 ( .A1(n_508), .A2(n_1322), .A3(n_1328), .B1(n_1333), .B2(n_1337), .B3(n_1343), .Y(n_1321) );
OAI33xp33_ASAP7_75t_L g1376 ( .A1(n_508), .A2(n_1343), .A3(n_1377), .B1(n_1381), .B2(n_1384), .B3(n_1388), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_508), .A2(n_1219), .B1(n_1421), .B2(n_1427), .Y(n_1420) );
OAI33xp33_ASAP7_75t_L g1460 ( .A1(n_508), .A2(n_538), .A3(n_1461), .B1(n_1466), .B2(n_1469), .B3(n_1472), .Y(n_1460) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
OR2x6_ASAP7_75t_L g652 ( .A(n_509), .B(n_511), .Y(n_652) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g821 ( .A(n_510), .Y(n_821) );
BUFx3_ASAP7_75t_L g1302 ( .A(n_510), .Y(n_1302) );
INVx2_ASAP7_75t_SL g1560 ( .A(n_510), .Y(n_1560) );
INVx1_ASAP7_75t_L g1950 ( .A(n_510), .Y(n_1950) );
INVx2_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
AND2x4_ASAP7_75t_L g724 ( .A(n_511), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g820 ( .A(n_511), .B(n_821), .Y(n_820) );
AND2x4_ASAP7_75t_L g914 ( .A(n_511), .B(n_725), .Y(n_914) );
BUFx2_ASAP7_75t_L g1134 ( .A(n_511), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_513), .A2(n_517), .B1(n_551), .B2(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_516), .A2(n_657), .B1(n_658), .B2(n_660), .Y(n_656) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_516), .Y(n_1106) );
INVx1_ASAP7_75t_L g1214 ( .A(n_516), .Y(n_1214) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g659 ( .A(n_520), .Y(n_659) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_520), .B(n_684), .Y(n_1313) );
OAI22xp33_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_523), .B1(n_525), .B2(n_526), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_522), .A2(n_525), .B1(n_546), .B2(n_547), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g1328 ( .A1(n_523), .A2(n_1329), .B1(n_1330), .B2(n_1332), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_523), .A2(n_1334), .B1(n_1335), .B2(n_1336), .Y(n_1333) );
OAI22xp33_ASAP7_75t_L g1381 ( .A1(n_523), .A2(n_1330), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_523), .A2(n_1216), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1469 ( .A1(n_523), .A2(n_1424), .B1(n_1470), .B2(n_1471), .Y(n_1469) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1370 ( .A(n_524), .Y(n_1370) );
INVx2_ASAP7_75t_L g1385 ( .A(n_524), .Y(n_1385) );
OAI221xp5_ASAP7_75t_L g1427 ( .A1(n_526), .A2(n_1422), .B1(n_1428), .B2(n_1429), .C(n_1430), .Y(n_1427) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g1217 ( .A(n_527), .Y(n_1217) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g531 ( .A(n_528), .Y(n_531) );
BUFx4f_ASAP7_75t_L g1292 ( .A(n_528), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_528), .Y(n_1331) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x6_ASAP7_75t_L g695 ( .A(n_531), .B(n_683), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_533) );
INVx2_ASAP7_75t_L g687 ( .A(n_535), .Y(n_687) );
INVx1_ASAP7_75t_L g994 ( .A(n_535), .Y(n_994) );
OAI22xp5_ASAP7_75t_SL g1570 ( .A1(n_538), .A2(n_652), .B1(n_1571), .B2(n_1576), .Y(n_1570) );
OAI22xp5_ASAP7_75t_L g1971 ( .A1(n_538), .A2(n_652), .B1(n_1972), .B2(n_1976), .Y(n_1971) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_539), .A2(n_641), .B1(n_651), .B2(n_653), .C(n_661), .Y(n_640) );
AOI33xp33_ASAP7_75t_L g929 ( .A1(n_539), .A2(n_930), .A3(n_931), .B1(n_936), .B2(n_938), .B3(n_940), .Y(n_929) );
AOI33xp33_ASAP7_75t_L g1033 ( .A1(n_539), .A2(n_930), .A3(n_1034), .B1(n_1037), .B2(n_1039), .B3(n_1042), .Y(n_1033) );
BUFx4f_ASAP7_75t_L g1109 ( .A(n_539), .Y(n_1109) );
BUFx4f_ASAP7_75t_L g1162 ( .A(n_539), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_540), .Y(n_1296) );
INVx2_ASAP7_75t_L g1548 ( .A(n_540), .Y(n_1548) );
INVx2_ASAP7_75t_SL g1940 ( .A(n_540), .Y(n_1940) );
AND2x4_ASAP7_75t_L g667 ( .A(n_541), .B(n_668), .Y(n_667) );
OAI33xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .A3(n_550), .B1(n_556), .B2(n_565), .B3(n_572), .Y(n_542) );
INVx1_ASAP7_75t_L g1253 ( .A(n_543), .Y(n_1253) );
OAI33xp33_ASAP7_75t_L g1521 ( .A1(n_543), .A2(n_1273), .A3(n_1522), .B1(n_1527), .B2(n_1535), .B3(n_1538), .Y(n_1521) );
OAI33xp33_ASAP7_75t_L g1915 ( .A1(n_543), .A2(n_1273), .A3(n_1916), .B1(n_1923), .B2(n_1926), .B3(n_1931), .Y(n_1915) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_546), .A2(n_566), .B1(n_567), .B2(n_571), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_546), .A2(n_569), .B1(n_1074), .B2(n_1075), .C(n_1076), .Y(n_1073) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_546), .A2(n_594), .B1(n_1063), .B2(n_1079), .C(n_1080), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_546), .Y(n_1270) );
INVx1_ASAP7_75t_L g1634 ( .A(n_546), .Y(n_1634) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_549), .B(n_612), .Y(n_611) );
OR2x6_ASAP7_75t_L g868 ( .A(n_549), .B(n_618), .Y(n_868) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_549), .B(n_618), .Y(n_1493) );
HB1xp67_ASAP7_75t_L g1922 ( .A(n_549), .Y(n_1922) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_551), .A2(n_1185), .B1(n_1379), .B2(n_1380), .Y(n_1397) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g987 ( .A(n_553), .Y(n_987) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g629 ( .A(n_554), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g866 ( .A(n_555), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_557), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_557), .A2(n_921), .B1(n_1325), .B2(n_1327), .Y(n_1350) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g1438 ( .A(n_558), .Y(n_1438) );
INVx2_ASAP7_75t_L g1446 ( .A(n_558), .Y(n_1446) );
INVx2_ASAP7_75t_L g1496 ( .A(n_558), .Y(n_1496) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g1263 ( .A(n_559), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_560), .A2(n_1260), .B1(n_1261), .B2(n_1264), .Y(n_1259) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g811 ( .A(n_562), .Y(n_811) );
INVx3_ASAP7_75t_L g1085 ( .A(n_562), .Y(n_1085) );
INVx2_ASAP7_75t_L g1929 ( .A(n_562), .Y(n_1929) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g590 ( .A(n_563), .Y(n_590) );
INVx3_ASAP7_75t_L g1186 ( .A(n_563), .Y(n_1186) );
OAI22xp33_ASAP7_75t_L g1931 ( .A1(n_567), .A2(n_1918), .B1(n_1932), .B2(n_1933), .Y(n_1931) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_569), .Y(n_1180) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_569), .A2(n_1076), .B1(n_1329), .B2(n_1332), .C(n_1352), .Y(n_1351) );
BUFx3_ASAP7_75t_L g1399 ( .A(n_569), .Y(n_1399) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI33xp33_ASAP7_75t_L g723 ( .A1(n_573), .A2(n_724), .A3(n_726), .B1(n_729), .B2(n_733), .B3(n_735), .Y(n_723) );
AOI33xp33_ASAP7_75t_L g912 ( .A1(n_573), .A2(n_913), .A3(n_915), .B1(n_918), .B2(n_923), .B3(n_928), .Y(n_912) );
AOI33xp33_ASAP7_75t_L g1028 ( .A1(n_573), .A2(n_724), .A3(n_1029), .B1(n_1030), .B2(n_1031), .B3(n_1032), .Y(n_1028) );
INVx6_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx5_ASAP7_75t_L g813 ( .A(n_574), .Y(n_813) );
OR2x6_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_575), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g683 ( .A(n_576), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g1232 ( .A(n_576), .B(n_624), .Y(n_1232) );
BUFx2_ASAP7_75t_L g607 ( .A(n_577), .Y(n_607) );
INVx2_ASAP7_75t_L g851 ( .A(n_577), .Y(n_851) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_583), .B(n_640), .C(n_678), .D(n_690), .Y(n_582) );
OAI31xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_621), .A3(n_632), .B(n_638), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_592), .B1(n_598), .B2(n_602), .C(n_608), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_589), .B2(n_591), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_586), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g1635 ( .A1(n_586), .A2(n_921), .B1(n_1636), .B2(n_1637), .Y(n_1635) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g1083 ( .A(n_587), .Y(n_1083) );
INVx1_ASAP7_75t_L g1356 ( .A(n_587), .Y(n_1356) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_588), .A2(n_591), .B1(n_648), .B2(n_650), .Y(n_647) );
INVx2_ASAP7_75t_L g734 ( .A(n_589), .Y(n_734) );
INVx2_ASAP7_75t_SL g804 ( .A(n_589), .Y(n_804) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g600 ( .A(n_590), .Y(n_600) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_590), .Y(n_845) );
INVx1_ASAP7_75t_L g1592 ( .A(n_590), .Y(n_1592) );
INVx2_ASAP7_75t_L g1988 ( .A(n_590), .Y(n_1988) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_595), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g1487 ( .A1(n_594), .A2(n_1467), .B1(n_1468), .B2(n_1488), .C(n_1491), .Y(n_1487) );
BUFx2_ASAP7_75t_L g727 ( .A(n_596), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_596), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g606 ( .A(n_597), .Y(n_606) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_597), .Y(n_1122) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_599), .A2(n_609), .B1(n_679), .B2(n_685), .C1(n_686), .C2(n_688), .Y(n_678) );
INVx1_ASAP7_75t_L g732 ( .A(n_600), .Y(n_732) );
INVx2_ASAP7_75t_L g982 ( .A(n_600), .Y(n_982) );
INVx1_ASAP7_75t_L g1486 ( .A(n_600), .Y(n_1486) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_601), .A2(n_603), .B1(n_691), .B2(n_694), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_605), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g1193 ( .A1(n_604), .A2(n_1194), .B(n_1195), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1538 ( .A1(n_604), .A2(n_1352), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
OAI221xp5_ASAP7_75t_L g1594 ( .A1(n_604), .A2(n_1270), .B1(n_1491), .B2(n_1572), .C(n_1573), .Y(n_1594) );
BUFx3_ASAP7_75t_L g916 ( .A(n_606), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .C(n_617), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g1248 ( .A(n_615), .B(n_1245), .Y(n_1248) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x6_ASAP7_75t_L g858 ( .A(n_616), .B(n_618), .Y(n_858) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g840 ( .A(n_618), .Y(n_840) );
INVx1_ASAP7_75t_L g857 ( .A(n_618), .Y(n_857) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_623), .A2(n_629), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx3_ASAP7_75t_L g1092 ( .A(n_623), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_623), .A2(n_629), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_623), .A2(n_629), .B1(n_1174), .B2(n_1175), .Y(n_1173) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_L g631 ( .A(n_624), .Y(n_631) );
INVx1_ASAP7_75t_L g731 ( .A(n_625), .Y(n_731) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_625), .Y(n_844) );
BUFx2_ASAP7_75t_L g919 ( .A(n_625), .Y(n_919) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_625), .Y(n_926) );
BUFx2_ASAP7_75t_L g986 ( .A(n_625), .Y(n_986) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g1093 ( .A(n_629), .Y(n_1093) );
AND2x4_ASAP7_75t_L g636 ( .A(n_630), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
CKINVDCx6p67_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_634), .A2(n_863), .B1(n_864), .B2(n_865), .C(n_867), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g1128 ( .A1(n_634), .A2(n_867), .B1(n_1129), .B2(n_1131), .C(n_1132), .Y(n_1128) );
AOI222xp33_ASAP7_75t_L g1168 ( .A1(n_634), .A2(n_636), .B1(n_1169), .B2(n_1170), .C1(n_1171), .C2(n_1172), .Y(n_1168) );
INVx8_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI221xp5_ASAP7_75t_SL g842 ( .A1(n_636), .A2(n_843), .B1(n_846), .B2(n_852), .C(n_853), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_636), .A2(n_1116), .B1(n_1119), .B2(n_1123), .C(n_1124), .Y(n_1115) );
INVx1_ASAP7_75t_L g849 ( .A(n_637), .Y(n_849) );
INVx1_ASAP7_75t_L g869 ( .A(n_638), .Y(n_869) );
OAI31xp33_ASAP7_75t_L g1628 ( .A1(n_638), .A2(n_1629), .A3(n_1630), .B(n_1638), .Y(n_1628) );
OAI31xp33_ASAP7_75t_L g1981 ( .A1(n_638), .A2(n_1982), .A3(n_1994), .B(n_2000), .Y(n_1981) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp67_ASAP7_75t_L g838 ( .A(n_639), .B(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g875 ( .A(n_643), .Y(n_875) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_646), .Y(n_655) );
INVx2_ASAP7_75t_L g745 ( .A(n_646), .Y(n_745) );
INVx2_ASAP7_75t_L g764 ( .A(n_646), .Y(n_764) );
INVx1_ASAP7_75t_L g824 ( .A(n_646), .Y(n_824) );
INVx2_ASAP7_75t_L g933 ( .A(n_646), .Y(n_933) );
INVx1_ASAP7_75t_L g1158 ( .A(n_646), .Y(n_1158) );
INVx2_ASAP7_75t_SL g1295 ( .A(n_646), .Y(n_1295) );
INVx1_ASAP7_75t_L g1035 ( .A(n_648), .Y(n_1035) );
INVx1_ASAP7_75t_L g1101 ( .A(n_648), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1472 ( .A1(n_648), .A2(n_1340), .B1(n_1473), .B2(n_1474), .Y(n_1472) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g937 ( .A(n_649), .Y(n_937) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_649), .B(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1943 ( .A(n_649), .Y(n_1943) );
INVx1_ASAP7_75t_L g1036 ( .A(n_650), .Y(n_1036) );
INVx1_ASAP7_75t_L g1043 ( .A(n_650), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1377 ( .A1(n_650), .A2(n_1378), .B1(n_1379), .B2(n_1380), .Y(n_1377) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_652), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_652), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_652), .A2(n_1207), .B1(n_1215), .B2(n_1219), .Y(n_1206) );
OAI22xp5_ASAP7_75t_SL g1616 ( .A1(n_652), .A2(n_1219), .B1(n_1617), .B2(n_1621), .Y(n_1616) );
INVx4_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g992 ( .A(n_655), .Y(n_992) );
INVx1_ASAP7_75t_L g1545 ( .A(n_655), .Y(n_1545) );
INVx1_ASAP7_75t_L g979 ( .A(n_658), .Y(n_979) );
INVx1_ASAP7_75t_L g995 ( .A(n_658), .Y(n_995) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g1944 ( .A(n_659), .Y(n_1944) );
INVx2_ASAP7_75t_L g887 ( .A(n_662), .Y(n_887) );
INVx1_ASAP7_75t_L g1058 ( .A(n_662), .Y(n_1058) );
INVx2_ASAP7_75t_L g1148 ( .A(n_662), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1582 ( .A(n_662), .Y(n_1582) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g1287 ( .A(n_664), .Y(n_1287) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
OR2x6_ASAP7_75t_L g671 ( .A(n_666), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_666), .Y(n_677) );
OR2x2_ASAP7_75t_L g1433 ( .A(n_666), .B(n_672), .Y(n_1433) );
AND2x4_ASAP7_75t_L g1286 ( .A(n_667), .B(n_1287), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_667), .B(n_673), .Y(n_1289) );
INVx1_ASAP7_75t_L g1308 ( .A(n_667), .Y(n_1308) );
AND2x4_ASAP7_75t_L g1553 ( .A(n_667), .B(n_1287), .Y(n_1553) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g885 ( .A(n_671), .Y(n_885) );
OR2x2_ASAP7_75t_L g1946 ( .A(n_672), .B(n_1308), .Y(n_1946) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g1146 ( .A(n_674), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_675), .Y(n_1160) );
BUFx2_ASAP7_75t_SL g1949 ( .A(n_675), .Y(n_1949) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g749 ( .A(n_676), .Y(n_749) );
INVx2_ASAP7_75t_SL g1013 ( .A(n_676), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_676), .Y(n_1038) );
BUFx4f_ASAP7_75t_L g1099 ( .A(n_676), .Y(n_1099) );
INVx1_ASAP7_75t_L g1204 ( .A(n_676), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_676), .B(n_1283), .Y(n_1305) );
AND2x2_ASAP7_75t_L g889 ( .A(n_677), .B(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_679), .A2(n_686), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_679), .A2(n_686), .B1(n_1062), .B2(n_1063), .C(n_1064), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_679), .A2(n_686), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g939 ( .A(n_681), .Y(n_939) );
AND2x2_ASAP7_75t_L g686 ( .A(n_682), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x6_ASAP7_75t_L g692 ( .A(n_683), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_683), .B(n_693), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_683), .B(n_1370), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_683), .B(n_1372), .Y(n_1371) );
INVx2_ASAP7_75t_L g1283 ( .A(n_684), .Y(n_1283) );
OR2x6_ASAP7_75t_L g837 ( .A(n_688), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g1278 ( .A(n_688), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_691), .A2(n_694), .B1(n_879), .B2(n_880), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_691), .A2(n_694), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
CKINVDCx6p67_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g873 ( .A(n_693), .Y(n_873) );
CKINVDCx6p67_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
OA22x2_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_770), .B1(n_771), .B2(n_828), .Y(n_696) );
INVx1_ASAP7_75t_L g828 ( .A(n_697), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_722), .C(n_753), .Y(n_699) );
AOI221x1_ASAP7_75t_L g772 ( .A1(n_700), .A2(n_773), .B1(n_786), .B2(n_788), .C(n_801), .Y(n_772) );
CKINVDCx16_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
AOI31xp33_ASAP7_75t_L g996 ( .A1(n_701), .A2(n_997), .A3(n_1001), .B(n_1004), .Y(n_996) );
AO21x1_ASAP7_75t_SL g1020 ( .A1(n_701), .A2(n_1021), .B(n_1025), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_705), .A2(n_707), .B1(n_790), .B2(n_791), .Y(n_789) );
INVx4_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx5_ASAP7_75t_L g954 ( .A(n_712), .Y(n_954) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g917 ( .A(n_716), .Y(n_917) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_717), .Y(n_728) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_738), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_724), .B(n_803), .C(n_805), .Y(n_802) );
BUFx2_ASAP7_75t_SL g1076 ( .A(n_725), .Y(n_1076) );
INVx1_ASAP7_75t_L g1492 ( .A(n_725), .Y(n_1492) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g808 ( .A(n_737), .Y(n_808) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_737), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .A3(n_743), .B1(n_746), .B2(n_750), .B3(n_752), .Y(n_738) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_752), .B(n_823), .C(n_825), .Y(n_822) );
AOI33xp33_ASAP7_75t_L g871 ( .A1(n_752), .A2(n_819), .A3(n_872), .B1(n_874), .B2(n_876), .B3(n_877), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_752), .B(n_991), .C(n_993), .Y(n_990) );
INVx1_ASAP7_75t_L g1343 ( .A(n_752), .Y(n_1343) );
AOI31xp33_ASAP7_75t_SL g753 ( .A1(n_754), .A2(n_761), .A3(n_765), .B(n_769), .Y(n_753) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g782 ( .A(n_758), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_766), .A2(n_775), .B1(n_909), .B2(n_910), .Y(n_908) );
CKINVDCx6p67_ASAP7_75t_R g1018 ( .A(n_766), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_766), .A2(n_775), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g827 ( .A(n_772), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
INVx1_ASAP7_75t_L g935 ( .A(n_785), .Y(n_935) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_785), .Y(n_1041) );
INVx1_ASAP7_75t_L g1300 ( .A(n_785), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1306 ( .A(n_785), .B(n_1307), .Y(n_1306) );
AOI221x1_ASAP7_75t_SL g1166 ( .A1(n_786), .A2(n_1134), .B1(n_1167), .B2(n_1196), .C(n_1206), .Y(n_1166) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AOI211x1_ASAP7_75t_SL g895 ( .A1(n_787), .A2(n_896), .B(n_911), .C(n_943), .Y(n_895) );
AO211x2_ASAP7_75t_L g961 ( .A1(n_787), .A2(n_962), .B(n_974), .C(n_996), .Y(n_961) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g801 ( .A(n_802), .B(n_809), .C(n_814), .D(n_822), .Y(n_801) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_812), .C(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g1440 ( .A(n_811), .Y(n_1440) );
NAND3xp33_ASAP7_75t_L g980 ( .A(n_813), .B(n_981), .C(n_983), .Y(n_980) );
CKINVDCx8_ASAP7_75t_R g1273 ( .A(n_813), .Y(n_1273) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .C(n_819), .Y(n_814) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g1103 ( .A(n_817), .Y(n_1103) );
INVx1_ASAP7_75t_L g1326 ( .A(n_817), .Y(n_1326) );
INVx1_ASAP7_75t_L g1464 ( .A(n_817), .Y(n_1464) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_819), .B(n_976), .C(n_977), .Y(n_975) );
INVx3_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_958), .B2(n_1046), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AOI21x1_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_893), .B(n_957), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g957 ( .A(n_833), .B(n_894), .Y(n_957) );
XOR2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_892), .Y(n_833) );
NOR3xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_841), .C(n_870), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_837), .B(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1143 ( .A(n_837), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_837), .B(n_1346), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_837), .B(n_1393), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_837), .B(n_1418), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_837), .B(n_1480), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_837), .B(n_1584), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_837), .B(n_1614), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g2001 ( .A(n_837), .B(n_2002), .Y(n_2001) );
INVx1_ASAP7_75t_L g1170 ( .A(n_839), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_840), .B(n_1089), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_840), .B(n_1089), .Y(n_1363) );
AOI31xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_859), .A3(n_862), .B(n_869), .Y(n_841) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1080 ( .A(n_850), .Y(n_1080) );
INVx2_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
NAND2x1p5_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .Y(n_854) );
NAND2x1_ASAP7_75t_SL g1244 ( .A(n_855), .B(n_1245), .Y(n_1244) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx11_ASAP7_75t_R g1090 ( .A(n_858), .Y(n_1090) );
INVx1_ASAP7_75t_L g1601 ( .A(n_866), .Y(n_1601) );
NOR3xp33_ASAP7_75t_L g1176 ( .A(n_867), .B(n_1177), .C(n_1191), .Y(n_1176) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_869), .A2(n_1275), .B1(n_1542), .B2(n_1563), .Y(n_1541) );
AOI22xp33_ASAP7_75t_L g1934 ( .A1(n_869), .A2(n_1275), .B1(n_1935), .B2(n_1953), .Y(n_1934) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_878), .C(n_881), .D(n_884), .Y(n_870) );
BUFx2_ASAP7_75t_L g1550 ( .A(n_873), .Y(n_1550) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B1(n_887), .B2(n_888), .C(n_889), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_885), .A2(n_889), .B1(n_1058), .B2(n_1059), .C(n_1060), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1147 ( .A1(n_885), .A2(n_1148), .B1(n_1149), .B2(n_1150), .Y(n_1147) );
INVx2_ASAP7_75t_L g1432 ( .A(n_887), .Y(n_1432) );
NOR3xp33_ASAP7_75t_L g1320 ( .A(n_889), .B(n_1321), .C(n_1344), .Y(n_1320) );
NOR3xp33_ASAP7_75t_L g1375 ( .A(n_889), .B(n_1376), .C(n_1391), .Y(n_1375) );
NOR3xp33_ASAP7_75t_SL g1419 ( .A(n_889), .B(n_1420), .C(n_1431), .Y(n_1419) );
NOR3xp33_ASAP7_75t_SL g1459 ( .A(n_889), .B(n_1460), .C(n_1475), .Y(n_1459) );
BUFx2_ASAP7_75t_L g1569 ( .A(n_889), .Y(n_1569) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g1557 ( .A(n_891), .Y(n_1557) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g956 ( .A(n_895), .Y(n_956) );
NAND4xp25_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .C(n_901), .D(n_908), .Y(n_896) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_897), .Y(n_1205) );
BUFx4f_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g967 ( .A(n_906), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_929), .Y(n_911) );
BUFx3_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_914), .B(n_985), .C(n_988), .Y(n_984) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g1192 ( .A(n_921), .Y(n_1192) );
OAI221xp5_ASAP7_75t_L g1445 ( .A1(n_921), .A2(n_1446), .B1(n_1447), .B2(n_1448), .C(n_1449), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g1495 ( .A1(n_921), .A2(n_1496), .B1(n_1497), .B2(n_1498), .C(n_1499), .Y(n_1495) );
INVx4_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
BUFx3_ASAP7_75t_L g927 ( .A(n_922), .Y(n_927) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_922), .Y(n_1071) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_922), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1358 ( .A(n_922), .Y(n_1358) );
INVx2_ASAP7_75t_SL g1405 ( .A(n_922), .Y(n_1405) );
INVx3_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_SL g925 ( .A(n_926), .Y(n_925) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_926), .B(n_1232), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_926), .B(n_1232), .Y(n_1518) );
INVx1_ASAP7_75t_L g1267 ( .A(n_927), .Y(n_1267) );
AOI33xp33_ASAP7_75t_L g1151 ( .A1(n_930), .A2(n_1152), .A3(n_1155), .B1(n_1159), .B2(n_1161), .B3(n_1162), .Y(n_1151) );
BUFx3_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_933), .Y(n_1040) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
BUFx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
BUFx4f_ASAP7_75t_L g978 ( .A(n_942), .Y(n_978) );
INVx1_ASAP7_75t_L g1372 ( .A(n_942), .Y(n_1372) );
INVx1_ASAP7_75t_L g1046 ( .A(n_958), .Y(n_1046) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
XNOR2x1_ASAP7_75t_L g959 ( .A(n_960), .B(n_1006), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_968), .C(n_971), .Y(n_962) );
NAND4xp25_ASAP7_75t_L g974 ( .A(n_975), .B(n_980), .C(n_984), .D(n_990), .Y(n_974) );
INVx1_ASAP7_75t_L g1641 ( .A(n_987), .Y(n_1641) );
AND4x1_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1020), .C(n_1028), .D(n_1033), .Y(n_1007) );
NAND4xp25_ASAP7_75t_L g1045 ( .A(n_1008), .B(n_1020), .C(n_1028), .D(n_1033), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1043), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1504), .B2(n_1652), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
XNOR2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1316), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1052), .B1(n_1163), .B2(n_1315), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1054), .B1(n_1110), .B2(n_1111), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
NAND4xp75_ASAP7_75t_SL g1055 ( .A(n_1056), .B(n_1065), .C(n_1067), .D(n_1096), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1061), .Y(n_1056) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1058), .Y(n_1627) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_1059), .A2(n_1060), .B1(n_1088), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1062), .A2(n_1082), .B1(n_1084), .B2(n_1086), .Y(n_1081) );
OAI31xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1077), .A3(n_1091), .B(n_1094), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_1088), .A2(n_1090), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_1088), .A2(n_1090), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1604 ( .A1(n_1088), .A2(n_1090), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_1088), .A2(n_1090), .B1(n_1645), .B2(n_1646), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_1090), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_1090), .A2(n_1363), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_1090), .A2(n_1363), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1991 ( .A1(n_1090), .A2(n_1363), .B1(n_1992), .B2(n_1993), .Y(n_1991) );
OAI31xp33_ASAP7_75t_L g1347 ( .A1(n_1094), .A2(n_1348), .A3(n_1349), .B(n_1354), .Y(n_1347) );
OAI31xp33_ASAP7_75t_L g1394 ( .A1(n_1094), .A2(n_1395), .A3(n_1396), .B(n_1402), .Y(n_1394) );
OAI31xp33_ASAP7_75t_L g1434 ( .A1(n_1094), .A2(n_1435), .A3(n_1436), .B(n_1444), .Y(n_1434) );
BUFx8_ASAP7_75t_SL g1094 ( .A(n_1095), .Y(n_1094) );
AOI33xp33_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1098), .A3(n_1100), .B1(n_1104), .B2(n_1105), .B3(n_1109), .Y(n_1096) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_1109), .Y(n_1219) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
XNOR2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
NOR4xp75_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1135), .C(n_1142), .D(n_1144), .Y(n_1113) );
AOI31xp33_ASAP7_75t_SL g1114 ( .A1(n_1115), .A2(n_1125), .A3(n_1128), .B(n_1133), .Y(n_1114) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
OAI22xp5_ASAP7_75t_SL g1996 ( .A1(n_1118), .A2(n_1997), .B1(n_1998), .B2(n_1999), .Y(n_1996) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
BUFx2_ASAP7_75t_L g1130 ( .A(n_1122), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1122), .B(n_1232), .Y(n_1238) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1133), .Y(n_1314) );
CKINVDCx8_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
OAI31xp33_ASAP7_75t_SL g1585 ( .A1(n_1134), .A2(n_1586), .A3(n_1587), .B(n_1595), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1139), .Y(n_1135) );
NAND3xp33_ASAP7_75t_SL g1144 ( .A(n_1145), .B(n_1147), .C(n_1151), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1154), .Y(n_1462) );
BUFx3_ASAP7_75t_L g1556 ( .A(n_1154), .Y(n_1556) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1163), .Y(n_1315) );
AOI22xp5_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1165), .B1(n_1222), .B2(n_1223), .Y(n_1163) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1166), .Y(n_1221) );
NAND3xp33_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1173), .C(n_1176), .Y(n_1167) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_1171), .A2(n_1172), .B1(n_1209), .B2(n_1216), .C(n_1218), .Y(n_1215) );
OAI21xp5_ASAP7_75t_SL g1177 ( .A1(n_1178), .A2(n_1182), .B(n_1188), .Y(n_1177) );
OAI21xp5_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1180), .B(n_1181), .Y(n_1178) );
BUFx3_ASAP7_75t_L g1526 ( .A(n_1180), .Y(n_1526) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .B1(n_1185), .B2(n_1187), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1926 ( .A1(n_1183), .A2(n_1927), .B1(n_1928), .B2(n_1930), .Y(n_1926) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_1186), .B(n_1232), .Y(n_1231) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_1187), .A2(n_1208), .B1(n_1211), .B2(n_1212), .C(n_1213), .Y(n_1207) );
NAND4xp25_ASAP7_75t_SL g1196 ( .A(n_1197), .B(n_1200), .C(n_1202), .D(n_1205), .Y(n_1196) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1571 ( .A1(n_1208), .A2(n_1572), .B1(n_1573), .B2(n_1574), .C(n_1575), .Y(n_1571) );
OAI221xp5_ASAP7_75t_L g1617 ( .A1(n_1208), .A2(n_1574), .B1(n_1618), .B2(n_1619), .C(n_1620), .Y(n_1617) );
OAI221xp5_ASAP7_75t_L g1972 ( .A1(n_1208), .A2(n_1574), .B1(n_1973), .B2(n_1974), .C(n_1975), .Y(n_1972) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_1216), .A2(n_1385), .B1(n_1386), .B2(n_1387), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1576 ( .A1(n_1216), .A2(n_1385), .B1(n_1577), .B2(n_1578), .C(n_1579), .Y(n_1576) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
XNOR2x1_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1225), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1274), .Y(n_1225) );
NOR3xp33_ASAP7_75t_SL g1226 ( .A(n_1227), .B(n_1241), .C(n_1251), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1236), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1230), .B1(n_1233), .B2(n_1234), .Y(n_1228) );
BUFx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
BUFx2_ASAP7_75t_L g1513 ( .A(n_1231), .Y(n_1513) );
BUFx2_ASAP7_75t_L g1908 ( .A(n_1231), .Y(n_1908) );
AND2x6_ASAP7_75t_L g1234 ( .A(n_1232), .B(n_1235), .Y(n_1234) );
OAI211xp5_ASAP7_75t_L g1290 ( .A1(n_1233), .A2(n_1291), .B(n_1293), .C(n_1294), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_1234), .A2(n_1512), .B1(n_1513), .B2(n_1514), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1906 ( .A1(n_1234), .A2(n_1907), .B1(n_1908), .B2(n_1909), .Y(n_1906) );
NAND2x1p5_ASAP7_75t_L g1250 ( .A(n_1235), .B(n_1245), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1238), .B1(n_1239), .B2(n_1240), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_1238), .A2(n_1516), .B1(n_1517), .B2(n_1518), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g1910 ( .A1(n_1238), .A2(n_1518), .B1(n_1911), .B2(n_1912), .Y(n_1910) );
INVx2_ASAP7_75t_SL g1242 ( .A(n_1243), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx3_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
BUFx4f_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
BUFx4f_ASAP7_75t_L g1914 ( .A(n_1248), .Y(n_1914) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1520 ( .A(n_1250), .Y(n_1520) );
OAI33xp33_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1254), .A3(n_1259), .B1(n_1265), .B2(n_1269), .B3(n_1273), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1265 ( .A1(n_1261), .A2(n_1266), .B1(n_1267), .B2(n_1268), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1588 ( .A1(n_1261), .A2(n_1589), .B1(n_1590), .B2(n_1593), .Y(n_1588) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx2_ASAP7_75t_L g1597 ( .A(n_1262), .Y(n_1597) );
INVx1_ASAP7_75t_L g1984 ( .A(n_1262), .Y(n_1984) );
INVx2_ASAP7_75t_L g1998 ( .A(n_1262), .Y(n_1998) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
AOI21xp5_ASAP7_75t_L g1281 ( .A1(n_1266), .A2(n_1282), .B(n_1284), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_1268), .A2(n_1271), .B1(n_1310), .B2(n_1312), .Y(n_1309) );
AOI221xp5_ASAP7_75t_L g1297 ( .A1(n_1272), .A2(n_1298), .B1(n_1303), .B2(n_1304), .C(n_1306), .Y(n_1297) );
AOI21xp33_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1279), .B(n_1280), .Y(n_1274) );
INVx5_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
AOI31xp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1297), .A3(n_1309), .B(n_1314), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_1282), .A2(n_1536), .B1(n_1544), .B2(n_1549), .C(n_1551), .Y(n_1543) );
AOI221xp5_ASAP7_75t_L g1936 ( .A1(n_1282), .A2(n_1927), .B1(n_1937), .B2(n_1941), .C(n_1945), .Y(n_1936) );
INVx1_ASAP7_75t_SL g1285 ( .A(n_1286), .Y(n_1285) );
INVx2_ASAP7_75t_SL g1288 ( .A(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1292), .Y(n_1335) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1292), .Y(n_1424) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_1304), .A2(n_1306), .B1(n_1540), .B2(n_1555), .C(n_1561), .Y(n_1554) );
AOI221xp5_ASAP7_75t_L g1947 ( .A1(n_1304), .A2(n_1306), .B1(n_1933), .B2(n_1948), .C(n_1951), .Y(n_1947) );
BUFx6f_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_SL g1307 ( .A(n_1308), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1562 ( .A1(n_1310), .A2(n_1312), .B1(n_1537), .B2(n_1539), .Y(n_1562) );
AOI22xp33_ASAP7_75t_L g1952 ( .A1(n_1310), .A2(n_1312), .B1(n_1930), .B2(n_1932), .Y(n_1952) );
INVx6_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx4_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
OAI31xp33_ASAP7_75t_L g1481 ( .A1(n_1314), .A2(n_1482), .A3(n_1483), .B(n_1494), .Y(n_1481) );
XNOR2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1414), .Y(n_1316) );
XOR2xp5_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1373), .Y(n_1317) );
AND4x1_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1345), .C(n_1347), .D(n_1365), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1325), .B1(n_1326), .B2(n_1327), .Y(n_1322) );
INVx2_ASAP7_75t_SL g1323 ( .A(n_1324), .Y(n_1323) );
BUFx3_ASAP7_75t_L g1625 ( .A(n_1324), .Y(n_1625) );
OAI22xp5_ASAP7_75t_L g1388 ( .A1(n_1326), .A2(n_1338), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
INVx2_ASAP7_75t_SL g1330 ( .A(n_1331), .Y(n_1330) );
BUFx2_ASAP7_75t_L g1574 ( .A(n_1335), .Y(n_1574) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1339), .B1(n_1340), .B2(n_1342), .Y(n_1337) );
INVx2_ASAP7_75t_SL g1340 ( .A(n_1341), .Y(n_1340) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1353), .Y(n_1524) );
OAI221xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B1(n_1358), .B2(n_1359), .C(n_1360), .Y(n_1355) );
OAI221xp5_ASAP7_75t_L g1403 ( .A1(n_1356), .A2(n_1404), .B1(n_1405), .B2(n_1406), .C(n_1407), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_1358), .A2(n_1529), .B1(n_1536), .B2(n_1537), .Y(n_1535) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1368), .Y(n_1365) );
AND4x1_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1392), .C(n_1394), .D(n_1411), .Y(n_1374) );
OAI21xp33_ASAP7_75t_SL g1398 ( .A1(n_1383), .A2(n_1399), .B(n_1400), .Y(n_1398) );
OAI221xp5_ASAP7_75t_L g1621 ( .A1(n_1385), .A2(n_1424), .B1(n_1622), .B2(n_1623), .C(n_1624), .Y(n_1621) );
OAI221xp5_ASAP7_75t_L g1976 ( .A1(n_1385), .A2(n_1424), .B1(n_1977), .B2(n_1978), .C(n_1979), .Y(n_1976) );
OAI21xp33_ASAP7_75t_L g1442 ( .A1(n_1399), .A2(n_1425), .B(n_1443), .Y(n_1442) );
NOR2xp33_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1413), .Y(n_1411) );
AO22x2_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1456), .B1(n_1457), .B2(n_1503), .Y(n_1414) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1415), .Y(n_1503) );
AND4x1_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .C(n_1434), .D(n_1453), .Y(n_1416) );
OAI221xp5_ASAP7_75t_L g1421 ( .A1(n_1422), .A2(n_1423), .B1(n_1424), .B2(n_1425), .C(n_1426), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1437 ( .A1(n_1438), .A2(n_1439), .B1(n_1440), .B2(n_1441), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g1484 ( .A1(n_1438), .A2(n_1463), .B1(n_1465), .B2(n_1485), .Y(n_1484) );
INVx2_ASAP7_75t_L g1530 ( .A(n_1446), .Y(n_1530) );
NOR2xp33_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1455), .Y(n_1453) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AND4x1_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1476), .C(n_1479), .D(n_1481), .Y(n_1458) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1463), .B1(n_1464), .B2(n_1465), .Y(n_1461) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1462), .Y(n_1580) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx2_ASAP7_75t_SL g1488 ( .A(n_1489), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1489 ( .A(n_1490), .Y(n_1489) );
OAI221xp5_ASAP7_75t_L g1631 ( .A1(n_1491), .A2(n_1618), .B1(n_1619), .B2(n_1632), .C(n_1633), .Y(n_1631) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g1923 ( .A1(n_1496), .A2(n_1590), .B1(n_1924), .B2(n_1925), .Y(n_1923) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1504), .Y(n_1652) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_1505), .A2(n_1564), .B1(n_1650), .B2(n_1651), .Y(n_1504) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1505), .Y(n_1650) );
HB1xp67_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1541), .Y(n_1508) );
NOR3xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1519), .C(n_1521), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1515), .Y(n_1510) );
OAI22xp33_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1524), .B1(n_1525), .B2(n_1526), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1529), .B1(n_1531), .B2(n_1532), .Y(n_1527) );
INVx2_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
NAND3xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1554), .C(n_1562), .Y(n_1542) );
BUFx2_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1564), .Y(n_1651) );
HB1xp67_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
XOR2x2_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1610), .Y(n_1565) );
AND4x1_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1583), .C(n_1585), .D(n_1607), .Y(n_1567) );
NOR3xp33_ASAP7_75t_SL g1568 ( .A(n_1569), .B(n_1570), .C(n_1581), .Y(n_1568) );
NOR3xp33_ASAP7_75t_SL g1615 ( .A(n_1569), .B(n_1616), .C(n_1626), .Y(n_1615) );
NOR3xp33_ASAP7_75t_L g1970 ( .A(n_1569), .B(n_1971), .C(n_1980), .Y(n_1970) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1596 ( .A1(n_1597), .A2(n_1598), .B1(n_1599), .B2(n_1602), .C(n_1603), .Y(n_1596) );
OAI221xp5_ASAP7_75t_L g1639 ( .A1(n_1597), .A2(n_1640), .B1(n_1641), .B2(n_1642), .C(n_1643), .Y(n_1639) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
NOR2xp33_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
XNOR2xp5_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1612), .Y(n_1610) );
AND4x1_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1615), .C(n_1628), .D(n_1647), .Y(n_1612) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
NOR2xp33_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1649), .Y(n_1647) );
OAI221xp5_ASAP7_75t_L g1653 ( .A1(n_1654), .A2(n_1898), .B1(n_1900), .B2(n_1955), .C(n_1960), .Y(n_1653) );
AOI21xp5_ASAP7_75t_L g1654 ( .A1(n_1655), .A2(n_1819), .B(n_1864), .Y(n_1654) );
NAND3xp33_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1737), .C(n_1758), .Y(n_1655) );
O2A1O1Ixp33_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1705), .B(n_1720), .C(n_1722), .Y(n_1656) );
O2A1O1Ixp33_ASAP7_75t_L g1737 ( .A1(n_1657), .A2(n_1738), .B(n_1741), .C(n_1743), .Y(n_1737) );
NOR2xp33_ASAP7_75t_SL g1657 ( .A(n_1658), .B(n_1701), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1679), .Y(n_1658) );
OAI21xp33_ASAP7_75t_L g1738 ( .A1(n_1659), .A2(n_1706), .B(n_1739), .Y(n_1738) );
INVx3_ASAP7_75t_L g1747 ( .A(n_1659), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1843 ( .A(n_1659), .B(n_1740), .Y(n_1843) );
NAND2xp5_ASAP7_75t_L g1877 ( .A(n_1659), .B(n_1775), .Y(n_1877) );
CKINVDCx5p33_ASAP7_75t_R g1659 ( .A(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1660), .Y(n_1721) );
INVx1_ASAP7_75t_SL g1731 ( .A(n_1660), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1660), .B(n_1729), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1660), .B(n_1740), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1660), .B(n_1701), .Y(n_1786) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1660), .Y(n_1832) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1660), .B(n_1681), .Y(n_1849) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1660), .Y(n_1872) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1669), .Y(n_1660) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1662), .Y(n_1812) );
AND2x4_ASAP7_75t_L g1662 ( .A(n_1663), .B(n_1666), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1663), .B(n_1666), .Y(n_1703) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AND2x4_ASAP7_75t_L g1668 ( .A(n_1664), .B(n_1666), .Y(n_1668) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1665), .B(n_1673), .Y(n_1672) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1667), .Y(n_1673) );
INVx2_ASAP7_75t_L g1712 ( .A(n_1668), .Y(n_1712) );
AND2x4_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1674), .Y(n_1670) );
OAI21xp33_ASAP7_75t_SL g2007 ( .A1(n_1671), .A2(n_1959), .B(n_2008), .Y(n_2007) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OR2x2_ASAP7_75t_L g1693 ( .A(n_1672), .B(n_1675), .Y(n_1693) );
AND2x4_ASAP7_75t_L g1676 ( .A(n_1674), .B(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1675), .B(n_1678), .Y(n_1695) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1679), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1688), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1885 ( .A(n_1680), .B(n_1718), .Y(n_1885) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1684), .Y(n_1680) );
INVx4_ASAP7_75t_L g1729 ( .A(n_1681), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1681), .B(n_1688), .Y(n_1742) );
INVx3_ASAP7_75t_L g1756 ( .A(n_1681), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1798 ( .A(n_1681), .B(n_1718), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1807 ( .A(n_1681), .B(n_1751), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1681), .B(n_1730), .Y(n_1828) );
NAND2xp5_ASAP7_75t_L g1860 ( .A(n_1681), .B(n_1762), .Y(n_1860) );
AND2x4_ASAP7_75t_L g1681 ( .A(n_1682), .B(n_1683), .Y(n_1681) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1684), .B(n_1767), .Y(n_1766) );
OR2x2_ASAP7_75t_L g1769 ( .A(n_1684), .B(n_1770), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1790 ( .A(n_1684), .B(n_1696), .Y(n_1790) );
OAI322xp33_ASAP7_75t_L g1826 ( .A1(n_1684), .A2(n_1748), .A3(n_1798), .B1(n_1827), .B2(n_1829), .C1(n_1830), .C2(n_1833), .Y(n_1826) );
NOR2xp33_ASAP7_75t_L g1839 ( .A(n_1684), .B(n_1696), .Y(n_1839) );
OR2x2_ASAP7_75t_L g1867 ( .A(n_1684), .B(n_1742), .Y(n_1867) );
OR2x2_ASAP7_75t_L g1875 ( .A(n_1684), .B(n_1734), .Y(n_1875) );
BUFx3_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1685), .B(n_1718), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1685), .B(n_1688), .Y(n_1724) );
INVx2_ASAP7_75t_L g1735 ( .A(n_1685), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1778 ( .A(n_1685), .B(n_1762), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1685), .B(n_1752), .Y(n_1823) );
AND2x2_ASAP7_75t_L g1834 ( .A(n_1685), .B(n_1734), .Y(n_1834) );
OR2x2_ASAP7_75t_L g1890 ( .A(n_1685), .B(n_1801), .Y(n_1890) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1688), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1688), .B(n_1782), .Y(n_1781) );
NAND2xp5_ASAP7_75t_L g1853 ( .A(n_1688), .B(n_1756), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1696), .Y(n_1688) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1689), .Y(n_1719) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1689), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1689), .B(n_1697), .Y(n_1752) );
OAI22xp33_ASAP7_75t_L g1690 ( .A1(n_1691), .A2(n_1692), .B1(n_1694), .B2(n_1695), .Y(n_1690) );
OAI22xp5_ASAP7_75t_L g1698 ( .A1(n_1692), .A2(n_1695), .B1(n_1699), .B2(n_1700), .Y(n_1698) );
OAI22xp33_ASAP7_75t_L g1713 ( .A1(n_1692), .A2(n_1714), .B1(n_1715), .B2(n_1716), .Y(n_1713) );
BUFx3_ASAP7_75t_L g1815 ( .A(n_1692), .Y(n_1815) );
BUFx6f_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
HB1xp67_ASAP7_75t_L g1716 ( .A(n_1695), .Y(n_1716) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1695), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1762 ( .A(n_1696), .B(n_1719), .Y(n_1762) );
INVx2_ASAP7_75t_L g1767 ( .A(n_1696), .Y(n_1767) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1697), .B(n_1719), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1701), .B(n_1709), .Y(n_1708) );
CKINVDCx5p33_ASAP7_75t_R g1725 ( .A(n_1701), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1701), .B(n_1731), .Y(n_1730) );
CKINVDCx6p67_ASAP7_75t_R g1740 ( .A(n_1701), .Y(n_1740) );
OR2x6_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1704), .Y(n_1701) );
INVxp67_ASAP7_75t_SL g1705 ( .A(n_1706), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1717), .Y(n_1706) );
OAI221xp5_ASAP7_75t_L g1804 ( .A1(n_1707), .A2(n_1747), .B1(n_1805), .B2(n_1806), .C(n_1808), .Y(n_1804) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_1708), .B(n_1832), .Y(n_1831) );
AOI221xp5_ASAP7_75t_L g1835 ( .A1(n_1708), .A2(n_1768), .B1(n_1836), .B2(n_1838), .C(n_1840), .Y(n_1835) );
OR2x2_ASAP7_75t_L g1739 ( .A(n_1709), .B(n_1740), .Y(n_1739) );
AND2x4_ASAP7_75t_SL g1775 ( .A(n_1709), .B(n_1740), .Y(n_1775) );
NAND2xp5_ASAP7_75t_L g1825 ( .A(n_1709), .B(n_1747), .Y(n_1825) );
NOR2xp33_ASAP7_75t_L g1859 ( .A(n_1709), .B(n_1729), .Y(n_1859) );
INVx2_ASAP7_75t_SL g1709 ( .A(n_1710), .Y(n_1709) );
INVx2_ASAP7_75t_L g1736 ( .A(n_1710), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1710), .B(n_1740), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1829 ( .A(n_1710), .B(n_1747), .Y(n_1829) );
INVx2_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1717), .Y(n_1841) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1718), .B(n_1729), .Y(n_1745) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1718), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1821 ( .A(n_1718), .B(n_1782), .Y(n_1821) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
O2A1O1Ixp33_ASAP7_75t_L g1722 ( .A1(n_1723), .A2(n_1725), .B(n_1726), .C(n_1736), .Y(n_1722) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1897 ( .A(n_1724), .B(n_1786), .Y(n_1897) );
AOI21xp33_ASAP7_75t_L g1850 ( .A1(n_1725), .A2(n_1851), .B(n_1854), .Y(n_1850) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1732), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1727), .B(n_1765), .Y(n_1791) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
NOR2xp33_ASAP7_75t_L g1800 ( .A(n_1728), .B(n_1801), .Y(n_1800) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1782 ( .A(n_1729), .B(n_1735), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1729), .B(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_L g1883 ( .A(n_1729), .Y(n_1883) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_1730), .B(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1730), .Y(n_1845) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1731), .B(n_1750), .Y(n_1749) );
NAND3xp33_ASAP7_75t_L g1847 ( .A(n_1732), .B(n_1740), .C(n_1848), .Y(n_1847) );
AOI322xp5_ASAP7_75t_L g1888 ( .A1(n_1732), .A2(n_1750), .A3(n_1836), .B1(n_1848), .B2(n_1889), .C1(n_1891), .C2(n_1893), .Y(n_1888) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
NAND2xp5_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1735), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1735), .B(n_1752), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1735), .B(n_1762), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1735), .B(n_1797), .Y(n_1796) );
OR2x2_ASAP7_75t_L g1852 ( .A(n_1735), .B(n_1853), .Y(n_1852) );
OAI321xp33_ASAP7_75t_L g1854 ( .A1(n_1735), .A2(n_1746), .A3(n_1809), .B1(n_1855), .B2(n_1858), .C(n_1860), .Y(n_1854) );
INVx2_ASAP7_75t_L g1748 ( .A(n_1736), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1736), .B(n_1786), .Y(n_1794) );
NAND3xp33_ASAP7_75t_L g1803 ( .A(n_1736), .B(n_1757), .C(n_1777), .Y(n_1803) );
INVx2_ASAP7_75t_L g1837 ( .A(n_1736), .Y(n_1837) );
AOI221xp5_ASAP7_75t_L g1878 ( .A1(n_1736), .A2(n_1779), .B1(n_1879), .B2(n_1880), .C(n_1886), .Y(n_1878) );
AND2x2_ASAP7_75t_L g1882 ( .A(n_1740), .B(n_1883), .Y(n_1882) );
A2O1A1Ixp33_ASAP7_75t_L g1870 ( .A1(n_1741), .A2(n_1775), .B(n_1821), .C(n_1871), .Y(n_1870) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
OAI221xp5_ASAP7_75t_L g1743 ( .A1(n_1744), .A2(n_1746), .B1(n_1749), .B2(n_1751), .C(n_1753), .Y(n_1743) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1748), .Y(n_1746) );
OR2x2_ASAP7_75t_L g1884 ( .A(n_1747), .B(n_1885), .Y(n_1884) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1748), .B(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1749), .Y(n_1893) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1750), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_1750), .B(n_1756), .Y(n_1771) );
AOI32xp33_ASAP7_75t_L g1861 ( .A1(n_1750), .A2(n_1757), .A3(n_1777), .B1(n_1786), .B2(n_1862), .Y(n_1861) );
NAND2xp5_ASAP7_75t_L g1856 ( .A(n_1751), .B(n_1857), .Y(n_1856) );
OAI21xp33_ASAP7_75t_L g1891 ( .A1(n_1751), .A2(n_1756), .B(n_1892), .Y(n_1891) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVxp67_ASAP7_75t_SL g1868 ( .A(n_1753), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1755), .B(n_1757), .Y(n_1754) );
INVx2_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
OR2x2_ASAP7_75t_L g1760 ( .A(n_1756), .B(n_1761), .Y(n_1760) );
AND2x2_ASAP7_75t_L g1822 ( .A(n_1756), .B(n_1823), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1838 ( .A(n_1756), .B(n_1839), .Y(n_1838) );
O2A1O1Ixp33_ASAP7_75t_SL g1886 ( .A1(n_1756), .A2(n_1793), .B(n_1806), .C(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1757), .Y(n_1789) );
NOR5xp2_ASAP7_75t_L g1758 ( .A(n_1759), .B(n_1783), .C(n_1792), .D(n_1802), .E(n_1804), .Y(n_1758) );
OAI221xp5_ASAP7_75t_L g1759 ( .A1(n_1760), .A2(n_1763), .B1(n_1764), .B2(n_1771), .C(n_1772), .Y(n_1759) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1760), .Y(n_1879) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1762), .Y(n_1857) );
NAND2xp5_ASAP7_75t_L g1863 ( .A(n_1762), .B(n_1782), .Y(n_1863) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1765), .B(n_1768), .Y(n_1764) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
OAI21xp33_ASAP7_75t_L g1880 ( .A1(n_1766), .A2(n_1881), .B(n_1884), .Y(n_1880) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
AOI22xp33_ASAP7_75t_SL g1772 ( .A1(n_1773), .A2(n_1778), .B1(n_1779), .B2(n_1780), .Y(n_1772) );
NAND2xp33_ASAP7_75t_L g1773 ( .A(n_1774), .B(n_1776), .Y(n_1773) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1778), .Y(n_1887) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
OAI211xp5_ASAP7_75t_L g1873 ( .A1(n_1782), .A2(n_1874), .B(n_1875), .C(n_1876), .Y(n_1873) );
OAI21xp5_ASAP7_75t_L g1783 ( .A1(n_1784), .A2(n_1787), .B(n_1791), .Y(n_1783) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
AOI221xp5_ASAP7_75t_L g1865 ( .A1(n_1786), .A2(n_1831), .B1(n_1866), .B2(n_1868), .C(n_1869), .Y(n_1865) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
NAND2xp5_ASAP7_75t_SL g1788 ( .A(n_1789), .B(n_1790), .Y(n_1788) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1790), .Y(n_1895) );
OAI21xp5_ASAP7_75t_L g1792 ( .A1(n_1793), .A2(n_1795), .B(n_1799), .Y(n_1792) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
NOR2xp33_ASAP7_75t_L g1844 ( .A(n_1798), .B(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVxp67_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx2_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
BUFx3_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
OAI22xp33_ASAP7_75t_L g1813 ( .A1(n_1814), .A2(n_1815), .B1(n_1816), .B2(n_1817), .Y(n_1813) );
INVx1_ASAP7_75t_L g1899 ( .A(n_1815), .Y(n_1899) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
NAND5xp2_ASAP7_75t_L g1819 ( .A(n_1820), .B(n_1835), .C(n_1842), .D(n_1850), .E(n_1861), .Y(n_1819) );
O2A1O1Ixp33_ASAP7_75t_L g1820 ( .A1(n_1821), .A2(n_1822), .B(n_1824), .C(n_1826), .Y(n_1820) );
AOI211xp5_ASAP7_75t_L g1842 ( .A1(n_1821), .A2(n_1843), .B(n_1844), .C(n_1846), .Y(n_1842) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1823), .Y(n_1892) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
A2O1A1Ixp33_ASAP7_75t_L g1894 ( .A1(n_1828), .A2(n_1837), .B(n_1895), .C(n_1896), .Y(n_1894) );
NOR2xp33_ASAP7_75t_L g1840 ( .A(n_1829), .B(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1853), .Y(n_1874) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
NAND4xp25_ASAP7_75t_L g1864 ( .A(n_1865), .B(n_1878), .C(n_1888), .D(n_1894), .Y(n_1864) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
NAND2xp5_ASAP7_75t_SL g1869 ( .A(n_1870), .B(n_1873), .Y(n_1869) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
INVxp33_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
INVxp67_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
CKINVDCx16_ASAP7_75t_R g1898 ( .A(n_1899), .Y(n_1898) );
INVx1_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
HB1xp67_ASAP7_75t_L g1902 ( .A(n_1903), .Y(n_1902) );
NAND2xp5_ASAP7_75t_L g1903 ( .A(n_1904), .B(n_1934), .Y(n_1903) );
NOR3xp33_ASAP7_75t_L g1904 ( .A(n_1905), .B(n_1913), .C(n_1915), .Y(n_1904) );
NAND2xp5_ASAP7_75t_L g1905 ( .A(n_1906), .B(n_1910), .Y(n_1905) );
OAI22xp33_ASAP7_75t_L g1916 ( .A1(n_1917), .A2(n_1918), .B1(n_1921), .B2(n_1922), .Y(n_1916) );
BUFx2_ASAP7_75t_L g1918 ( .A(n_1919), .Y(n_1918) );
INVx2_ASAP7_75t_L g1919 ( .A(n_1920), .Y(n_1919) );
INVx1_ASAP7_75t_L g1928 ( .A(n_1929), .Y(n_1928) );
NAND3xp33_ASAP7_75t_L g1935 ( .A(n_1936), .B(n_1947), .C(n_1952), .Y(n_1935) );
INVx1_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
INVx1_ASAP7_75t_L g1939 ( .A(n_1940), .Y(n_1939) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
CKINVDCx14_ASAP7_75t_R g1955 ( .A(n_1956), .Y(n_1955) );
INVx2_ASAP7_75t_L g1956 ( .A(n_1957), .Y(n_1956) );
CKINVDCx5p33_ASAP7_75t_R g1957 ( .A(n_1958), .Y(n_1957) );
INVx1_ASAP7_75t_L g1961 ( .A(n_1962), .Y(n_1961) );
INVx1_ASAP7_75t_L g1962 ( .A(n_1963), .Y(n_1962) );
INVx1_ASAP7_75t_L g1963 ( .A(n_1964), .Y(n_1963) );
INVx1_ASAP7_75t_L g1964 ( .A(n_1965), .Y(n_1964) );
INVx1_ASAP7_75t_L g1966 ( .A(n_1967), .Y(n_1966) );
INVx1_ASAP7_75t_L g1967 ( .A(n_1968), .Y(n_1967) );
AND4x1_ASAP7_75t_L g1969 ( .A(n_1970), .B(n_1981), .C(n_2001), .D(n_2003), .Y(n_1969) );
OAI221xp5_ASAP7_75t_L g1983 ( .A1(n_1984), .A2(n_1985), .B1(n_1986), .B2(n_1989), .C(n_1990), .Y(n_1983) );
INVx1_ASAP7_75t_L g1986 ( .A(n_1987), .Y(n_1986) );
INVx2_ASAP7_75t_L g1987 ( .A(n_1988), .Y(n_1987) );
NOR2xp33_ASAP7_75t_L g2003 ( .A(n_2004), .B(n_2005), .Y(n_2003) );
HB1xp67_ASAP7_75t_L g2006 ( .A(n_2007), .Y(n_2006) );
endmodule