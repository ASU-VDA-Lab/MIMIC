module fake_jpeg_3467_n_231 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_24),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_84),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_2),
.CON(n_84),
.SN(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_59),
.B1(n_70),
.B2(n_66),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_90),
.B1(n_94),
.B2(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_70),
.B1(n_59),
.B2(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_63),
.B1(n_76),
.B2(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_64),
.B1(n_57),
.B2(n_69),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_71),
.B1(n_55),
.B2(n_68),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_71),
.B1(n_55),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_74),
.B1(n_76),
.B2(n_64),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_64),
.B1(n_85),
.B2(n_54),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_86),
.B1(n_85),
.B2(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_116),
.B1(n_92),
.B2(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_35),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_52),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_80),
.B1(n_82),
.B2(n_53),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_108),
.B1(n_114),
.B2(n_118),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_85),
.B1(n_79),
.B2(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_58),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_78),
.C(n_61),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_77),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_61),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_57),
.B1(n_77),
.B2(n_58),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_119),
.Y(n_149)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_134),
.Y(n_159)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_72),
.Y(n_130)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_48),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_60),
.B(n_56),
.C(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_2),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_3),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_50),
.C(n_49),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_120),
.C(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_29),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_152),
.B1(n_154),
.B2(n_120),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_23),
.B(n_25),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_156),
.B1(n_122),
.B2(n_120),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_17),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_30),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_123),
.B(n_137),
.C(n_128),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_163),
.B(n_20),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_18),
.B(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_18),
.B(n_19),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_120),
.B(n_21),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_170),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_174),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_132),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_162),
.B1(n_161),
.B2(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_176),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_20),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_156),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_47),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_22),
.B(n_23),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_153),
.B1(n_163),
.B2(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_197),
.B1(n_183),
.B2(n_178),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_155),
.B1(n_150),
.B2(n_143),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_177),
.B1(n_172),
.B2(n_167),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.C(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_166),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_186),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_144),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_196),
.C(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_203),
.B(n_197),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_194),
.B(n_205),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_220),
.B(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_190),
.B1(n_198),
.B2(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_222),
.B1(n_215),
.B2(n_217),
.Y(n_224)
);

OAI211xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_216),
.C(n_212),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_178),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_168),
.A3(n_142),
.B1(n_27),
.B2(n_28),
.C1(n_25),
.C2(n_26),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_142),
.A3(n_26),
.B1(n_28),
.B2(n_174),
.C(n_39),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_34),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_42),
.Y(n_231)
);


endmodule