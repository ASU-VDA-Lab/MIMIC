module fake_jpeg_14374_n_222 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

XNOR2x1_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_16),
.Y(n_49)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_45),
.B(n_49),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_1),
.B(n_2),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_70),
.Y(n_82)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_0),
.Y(n_86)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_27),
.B1(n_14),
.B2(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_40),
.B1(n_34),
.B2(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_23),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_30),
.B(n_26),
.C(n_25),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_36),
.B(n_17),
.C(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_23),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_41),
.B1(n_33),
.B2(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_53),
.B1(n_64),
.B2(n_47),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_98),
.B1(n_104),
.B2(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_61),
.Y(n_118)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_54),
.B(n_64),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_93),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_102),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_35),
.B1(n_31),
.B2(n_3),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_7),
.B(n_10),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_1),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_97),
.B1(n_99),
.B2(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_116),
.Y(n_133)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_129),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_128),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_80),
.B(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_47),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_58),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_62),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.C(n_95),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_68),
.C(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_7),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_96),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_126),
.B(n_118),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_86),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_103),
.C(n_87),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_102),
.B1(n_92),
.B2(n_81),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_146),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_109),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_92),
.B1(n_85),
.B2(n_83),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_148),
.B(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_87),
.C(n_80),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_89),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_11),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_116),
.B(n_108),
.C(n_105),
.D(n_127),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_161),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_149),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_166),
.C(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_149),
.B(n_146),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_117),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_125),
.A3(n_128),
.B1(n_109),
.B2(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_120),
.B1(n_131),
.B2(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_132),
.B1(n_111),
.B2(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_154),
.A2(n_74),
.B1(n_110),
.B2(n_113),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_164),
.B1(n_137),
.B2(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_178),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_158),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_152),
.B(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_143),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_133),
.C(n_153),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_167),
.A3(n_168),
.B1(n_166),
.B2(n_163),
.C1(n_141),
.C2(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_150),
.C(n_138),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.C(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_137),
.C(n_119),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_178),
.CI(n_179),
.CON(n_186),
.SN(n_186)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.C(n_195),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_182),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_141),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_196),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_185),
.B(n_172),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_197),
.B(n_195),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_174),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_183),
.B(n_175),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_190),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_202),
.B(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_210),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_193),
.B1(n_175),
.B2(n_187),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_201),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_207),
.B1(n_187),
.B2(n_180),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_159),
.B(n_119),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_207),
.B(n_186),
.C(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_159),
.B(n_13),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_219),
.B(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_216),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_12),
.Y(n_222)
);


endmodule