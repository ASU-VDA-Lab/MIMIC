module fake_jpeg_29415_n_311 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_17),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_22),
.B1(n_24),
.B2(n_13),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_29),
.B1(n_13),
.B2(n_15),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_60),
.B1(n_15),
.B2(n_36),
.Y(n_81)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_13),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_28),
.B1(n_22),
.B2(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_41),
.C(n_45),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_71),
.C(n_54),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_45),
.B(n_18),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_31),
.B(n_30),
.C(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_30),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_81),
.B1(n_36),
.B2(n_39),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_39),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_57),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_30),
.Y(n_123)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_52),
.C(n_62),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_83),
.C(n_40),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_49),
.B1(n_47),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_76),
.B1(n_71),
.B2(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_77),
.B1(n_69),
.B2(n_67),
.Y(n_108)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_39),
.B1(n_61),
.B2(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_36),
.B1(n_39),
.B2(n_83),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_55),
.B1(n_46),
.B2(n_56),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_90),
.B(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_89),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_112),
.B1(n_103),
.B2(n_16),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_82),
.B(n_64),
.C(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_82),
.B1(n_64),
.B2(n_80),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_85),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_75),
.B1(n_78),
.B2(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_103),
.B1(n_22),
.B2(n_53),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_72),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.C(n_134),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_30),
.CI(n_40),
.CON(n_122),
.SN(n_122)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_29),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_63),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_130),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_63),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_61),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_40),
.B1(n_48),
.B2(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_44),
.B1(n_34),
.B2(n_21),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_97),
.C(n_96),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_92),
.C(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_103),
.C(n_98),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_166),
.C(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_150),
.B1(n_159),
.B2(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_14),
.A3(n_18),
.B1(n_19),
.B2(n_12),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_30),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_160),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_30),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_22),
.B1(n_24),
.B2(n_36),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_143),
.B1(n_137),
.B2(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_22),
.B1(n_23),
.B2(n_51),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_156)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_22),
.B1(n_23),
.B2(n_51),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_30),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_19),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_23),
.B1(n_12),
.B2(n_16),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_110),
.B(n_33),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_29),
.C(n_26),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_14),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_155),
.B1(n_165),
.B2(n_124),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_130),
.B1(n_107),
.B2(n_110),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_178),
.C(n_182),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_121),
.C(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_129),
.C(n_111),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_176),
.B1(n_188),
.B2(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_146),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_159),
.B1(n_142),
.B2(n_177),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_26),
.C(n_44),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_44),
.C(n_26),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_21),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_160),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_198),
.B(n_12),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_16),
.B(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_139),
.B1(n_176),
.B2(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

NAND2x1_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_139),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_220),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_182),
.B(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_216),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_21),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_145),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_184),
.B1(n_173),
.B2(n_195),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_218),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_150),
.B1(n_152),
.B2(n_149),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_166),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_221),
.B(n_185),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_1),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_192),
.C(n_186),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_238),
.C(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_242),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_190),
.B(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_183),
.C(n_26),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_217),
.B1(n_200),
.B2(n_199),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_33),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_215),
.CI(n_202),
.CON(n_242),
.SN(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_33),
.B(n_2),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_1),
.B(n_2),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_239),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_201),
.B(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_222),
.C(n_218),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_34),
.C(n_33),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_253),
.C(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_34),
.C(n_33),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_1),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_258),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_233),
.A2(n_33),
.B(n_3),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_259),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_34),
.C(n_33),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_232),
.A2(n_33),
.B(n_3),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_231),
.B1(n_234),
.B2(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_236),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_239),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_270),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_242),
.B(n_229),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_276),
.C(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_242),
.B(n_240),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_5),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_257),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_276),
.B(n_4),
.Y(n_290)
);

AOI21x1_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_253),
.B(n_241),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_21),
.C(n_23),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_2),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_262),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_271),
.B1(n_275),
.B2(n_273),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_266),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_290),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_3),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_5),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_5),
.B(n_6),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_6),
.B(n_7),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_6),
.C(n_7),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_302),
.B(n_10),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_7),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_11),
.C(n_8),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_294),
.B(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_301),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.C(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_300),
.C(n_308),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_10),
.B(n_8),
.Y(n_311)
);


endmodule