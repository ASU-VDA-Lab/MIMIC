module fake_aes_2081_n_1081 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1081);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1081;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_1042;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1025;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_818;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_1069;
wire n_1021;
wire n_972;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_100), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_272), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_188), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_13), .Y(n_279) );
BUFx2_ASAP7_75t_SL g280 ( .A(n_166), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_250), .B(n_43), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_178), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_273), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_114), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_84), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_145), .Y(n_288) );
NOR2xp67_ASAP7_75t_L g289 ( .A(n_85), .B(n_82), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_34), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_44), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_53), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_57), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_104), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_8), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_36), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_63), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_123), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_187), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_63), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_243), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_247), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_141), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_189), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_143), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_174), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_21), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_62), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_205), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_5), .Y(n_310) );
INVxp33_ASAP7_75t_SL g311 ( .A(n_254), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_211), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_175), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_101), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_0), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_115), .B(n_12), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_69), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_139), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_218), .Y(n_319) );
INVxp33_ASAP7_75t_SL g320 ( .A(n_164), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_190), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_199), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_17), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_216), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_161), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_86), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_10), .Y(n_327) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_185), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_230), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_28), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_105), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_274), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_186), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_245), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_156), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_87), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_176), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_116), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_253), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_56), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_12), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_195), .Y(n_344) );
INVx4_ASAP7_75t_R g345 ( .A(n_73), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_165), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_130), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_94), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_58), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_0), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_242), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_268), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_237), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_182), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_44), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_57), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_142), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_64), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_266), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_269), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_252), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_16), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_62), .Y(n_363) );
INVxp33_ASAP7_75t_L g364 ( .A(n_263), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_98), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_97), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_198), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_146), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_30), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_118), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_92), .Y(n_371) );
INVxp33_ASAP7_75t_SL g372 ( .A(n_22), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_207), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_23), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_217), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_260), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_83), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_167), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_258), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_179), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_204), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_257), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_72), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_36), .Y(n_384) );
CKINVDCx14_ASAP7_75t_R g385 ( .A(n_18), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_222), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_241), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_265), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_38), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_6), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_240), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_159), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_128), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_89), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_184), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_70), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_39), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_223), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_80), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_231), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_150), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_2), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_206), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_171), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_45), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_214), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_219), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_249), .Y(n_408) );
INVxp33_ASAP7_75t_L g409 ( .A(n_56), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_103), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_102), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_233), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_208), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_96), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_122), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_248), .Y(n_416) );
BUFx2_ASAP7_75t_SL g417 ( .A(n_246), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_284), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_298), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_303), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_284), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_356), .B(n_1), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_356), .B(n_1), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_303), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_319), .B(n_2), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_296), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_385), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_299), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_297), .B(n_3), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_305), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_319), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_299), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_305), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_298), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_335), .B(n_4), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_351), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_297), .B(n_6), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_304), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_310), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_310), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_304), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_323), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_409), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_341), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_409), .B(n_7), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_323), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_341), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_389), .B(n_9), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_296), .B(n_10), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_452), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_431), .B(n_359), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_438), .B(n_359), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_420), .B(n_348), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_439), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_420), .A2(n_278), .B(n_277), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_424), .B(n_364), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_452), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_427), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_452), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_419), .Y(n_466) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_429), .B(n_276), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_434), .B(n_348), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_433), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_434), .B(n_364), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_425), .B(n_365), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_423), .Y(n_478) );
AND2x6_ASAP7_75t_L g479 ( .A(n_423), .B(n_395), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_437), .B(n_384), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_436), .B(n_374), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_437), .Y(n_482) );
NOR2xp33_ASAP7_75t_SL g483 ( .A(n_446), .B(n_276), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_418), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_418), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_442), .B(n_346), .Y(n_487) );
INVx4_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_421), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_440), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_442), .B(n_443), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_459), .B(n_448), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_474), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_478), .Y(n_495) );
OR2x6_ASAP7_75t_L g496 ( .A(n_471), .B(n_451), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_465), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_467), .Y(n_498) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_471), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_477), .B(n_422), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_473), .B(n_384), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_453), .A2(n_421), .B1(n_432), .B2(n_428), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_455), .B(n_294), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_471), .B(n_311), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_454), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_465), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_467), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_483), .A2(n_372), .B1(n_338), .B2(n_370), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_480), .B(n_301), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_492), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_457), .Y(n_512) );
OR2x2_ASAP7_75t_SL g513 ( .A(n_461), .B(n_342), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_479), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_479), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_475), .B(n_337), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_484), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_478), .B(n_292), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_488), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_472), .B(n_282), .Y(n_521) );
NAND2xp33_ASAP7_75t_L g522 ( .A(n_479), .B(n_301), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_484), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_465), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_476), .B(n_337), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_476), .B(n_311), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_481), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_463), .B(n_306), .Y(n_530) );
BUFx12f_ASAP7_75t_L g531 ( .A(n_481), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_460), .A2(n_428), .B(n_444), .C(n_432), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_479), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_487), .B(n_338), .Y(n_534) );
INVx5_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
XNOR2xp5_ASAP7_75t_L g536 ( .A(n_461), .B(n_342), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_466), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_462), .B(n_283), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_491), .B(n_320), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_464), .B(n_469), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_487), .B(n_377), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_458), .B(n_306), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_456), .A2(n_355), .B(n_441), .C(n_432), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_466), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_470), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_458), .B(n_317), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_466), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_470), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_466), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_468), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_468), .B(n_317), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_490), .B(n_324), .Y(n_555) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_490), .B(n_349), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_459), .B(n_324), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_465), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_500), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_515), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_515), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_500), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_494), .B(n_426), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_494), .B(n_320), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_529), .B(n_308), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_495), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_541), .A2(n_328), .B(n_302), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_506), .B(n_428), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_506), .B(n_349), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_493), .B(n_444), .Y(n_571) );
CKINVDCx6p67_ASAP7_75t_R g572 ( .A(n_531), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_556), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_535), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_501), .A2(n_450), .B1(n_447), .B2(n_444), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_501), .B(n_326), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_535), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_557), .B(n_326), .Y(n_580) );
BUFx8_ASAP7_75t_SL g581 ( .A(n_512), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_551), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_556), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_541), .A2(n_378), .B(n_376), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_539), .A2(n_286), .B(n_285), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_537), .Y(n_587) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_516), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_511), .A2(n_450), .B1(n_447), .B2(n_290), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_537), .Y(n_590) );
INVx6_ASAP7_75t_L g591 ( .A(n_518), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_539), .A2(n_288), .B(n_287), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_532), .A2(n_291), .B(n_293), .C(n_279), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g594 ( .A1(n_513), .A2(n_397), .B1(n_330), .B2(n_295), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_526), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_532), .A2(n_300), .B(n_315), .C(n_307), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_536), .B(n_443), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_540), .B(n_327), .Y(n_598) );
CKINVDCx14_ASAP7_75t_R g599 ( .A(n_509), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_535), .B(n_333), .Y(n_600) );
OR2x6_ASAP7_75t_SL g601 ( .A(n_534), .B(n_333), .Y(n_601) );
INVx3_ASAP7_75t_SL g602 ( .A(n_498), .Y(n_602) );
AOI21x1_ASAP7_75t_L g603 ( .A1(n_543), .A2(n_450), .B(n_447), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_505), .B(n_336), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_503), .A2(n_350), .B1(n_358), .B2(n_343), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_496), .B(n_362), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_534), .B(n_445), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_520), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_508), .A2(n_374), .B1(n_390), .B2(n_363), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_502), .B(n_445), .Y(n_611) );
AO32x2_ASAP7_75t_L g612 ( .A1(n_503), .A2(n_435), .A3(n_419), .B1(n_280), .B2(n_417), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_505), .B(n_402), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_516), .B(n_449), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_540), .B(n_405), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_517), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_496), .B(n_449), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_525), .B(n_280), .Y(n_618) );
INVx3_ASAP7_75t_SL g619 ( .A(n_542), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_514), .B(n_336), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_354), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_527), .A2(n_309), .B1(n_313), .B2(n_312), .Y(n_622) );
BUFx12f_ASAP7_75t_L g623 ( .A(n_525), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_521), .B(n_281), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_554), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_544), .Y(n_626) );
AND2x2_ASAP7_75t_SL g627 ( .A(n_522), .B(n_316), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_547), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_527), .A2(n_314), .B1(n_321), .B2(n_318), .Y(n_629) );
INVx4_ASAP7_75t_L g630 ( .A(n_496), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_530), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_514), .B(n_396), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_550), .Y(n_633) );
NAND2x1_ASAP7_75t_SL g634 ( .A(n_523), .B(n_289), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_504), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_545), .A2(n_325), .B(n_329), .C(n_322), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_533), .B(n_399), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_521), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_510), .A2(n_332), .B(n_331), .Y(n_639) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_548), .A2(n_339), .B(n_334), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_553), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_533), .B(n_400), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_555), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_SL g644 ( .A1(n_552), .A2(n_344), .B(n_347), .C(n_340), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_524), .B(n_412), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_538), .B(n_360), .Y(n_646) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_546), .A2(n_353), .B(n_352), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_497), .B(n_360), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_625), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_568), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_639), .A2(n_549), .B(n_499), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_572), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_613), .A2(n_499), .B(n_497), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_625), .Y(n_654) );
OAI21x1_ASAP7_75t_L g655 ( .A1(n_603), .A2(n_379), .B(n_365), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_566), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_630), .B(n_357), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_584), .A2(n_371), .B1(n_367), .B2(n_361), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_625), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_569), .B(n_367), .Y(n_660) );
INVx4_ASAP7_75t_L g661 ( .A(n_584), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_573), .Y(n_662) );
AND2x4_ASAP7_75t_SL g663 ( .A(n_630), .B(n_497), .Y(n_663) );
INVx5_ASAP7_75t_L g664 ( .A(n_618), .Y(n_664) );
OAI21x1_ASAP7_75t_L g665 ( .A1(n_641), .A2(n_382), .B(n_379), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_643), .A2(n_392), .B(n_382), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_581), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_568), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_563), .A2(n_368), .B(n_366), .Y(n_669) );
OA21x2_ASAP7_75t_L g670 ( .A1(n_647), .A2(n_416), .B(n_394), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_593), .A2(n_375), .B(n_380), .C(n_373), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_571), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_563), .A2(n_383), .B(n_381), .Y(n_673) );
OAI21x1_ASAP7_75t_L g674 ( .A1(n_616), .A2(n_387), .B(n_386), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_571), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_582), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_576), .A2(n_391), .B1(n_393), .B2(n_388), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_560), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_613), .A2(n_398), .B(n_403), .C(n_401), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_594), .A2(n_371), .B1(n_417), .B2(n_404), .Y(n_680) );
OR2x6_ASAP7_75t_L g681 ( .A(n_618), .B(n_406), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_619), .B(n_407), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_601), .A2(n_414), .B1(n_408), .B2(n_410), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_604), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_623), .B(n_411), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_598), .A2(n_413), .B1(n_415), .B2(n_435), .C(n_497), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_596), .A2(n_435), .B(n_507), .C(n_499), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_611), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_560), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_617), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_617), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_564), .B(n_507), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_561), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_640), .A2(n_558), .B(n_507), .Y(n_695) );
AO21x2_ASAP7_75t_L g696 ( .A1(n_640), .A2(n_435), .B(n_558), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_626), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_589), .A2(n_345), .B(n_13), .C(n_14), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_570), .A2(n_558), .B(n_435), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_628), .A2(n_68), .B(n_67), .Y(n_700) );
CKINVDCx6p67_ASAP7_75t_R g701 ( .A(n_602), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_633), .Y(n_702) );
OAI21x1_ASAP7_75t_L g703 ( .A1(n_590), .A2(n_74), .B(n_71), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_648), .A2(n_76), .B(n_75), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_594), .A2(n_11), .B1(n_14), .B2(n_15), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_574), .Y(n_706) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_579), .A2(n_78), .B(n_77), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_615), .A2(n_15), .B(n_16), .C(n_17), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_614), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_576), .Y(n_710) );
INVx6_ASAP7_75t_L g711 ( .A(n_591), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_627), .A2(n_18), .B(n_19), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_618), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_713) );
OA21x2_ASAP7_75t_L g714 ( .A1(n_647), .A2(n_81), .B(n_79), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_609), .Y(n_715) );
OAI21x1_ASAP7_75t_L g716 ( .A1(n_579), .A2(n_90), .B(n_88), .Y(n_716) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_587), .A2(n_93), .B(n_91), .Y(n_717) );
AO32x2_ASAP7_75t_L g718 ( .A1(n_606), .A2(n_612), .A3(n_644), .B1(n_634), .B2(n_624), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_631), .B(n_20), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_599), .B(n_22), .C(n_23), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_636), .A2(n_24), .B(n_25), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_564), .B(n_635), .Y(n_722) );
INVx4_ASAP7_75t_L g723 ( .A(n_587), .Y(n_723) );
BUFx8_ASAP7_75t_L g724 ( .A(n_565), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_565), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_597), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_607), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_622), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_728) );
AO21x2_ASAP7_75t_L g729 ( .A1(n_612), .A2(n_99), .B(n_95), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_588), .B(n_26), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_607), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_621), .B(n_27), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_577), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_586), .A2(n_107), .B(n_106), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_608), .Y(n_736) );
OAI21x1_ASAP7_75t_L g737 ( .A1(n_592), .A2(n_109), .B(n_108), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_595), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_595), .B(n_29), .Y(n_739) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_606), .B(n_610), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_638), .Y(n_741) );
NOR2xp67_ASAP7_75t_SL g742 ( .A(n_561), .B(n_31), .Y(n_742) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_600), .A2(n_153), .B(n_270), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_622), .B(n_32), .Y(n_744) );
CKINVDCx11_ASAP7_75t_R g745 ( .A(n_575), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_605), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_746) );
BUFx3_ASAP7_75t_L g747 ( .A(n_562), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_580), .B(n_33), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_567), .A2(n_154), .B(n_267), .Y(n_749) );
OAI21x1_ASAP7_75t_L g750 ( .A1(n_585), .A2(n_152), .B(n_264), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_701), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_719), .A2(n_642), .B1(n_637), .B2(n_632), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_683), .A2(n_629), .B1(n_642), .B2(n_637), .C(n_632), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_695), .A2(n_629), .B(n_645), .Y(n_754) );
BUFx8_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
BUFx2_ASAP7_75t_L g756 ( .A(n_724), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_688), .A2(n_620), .B1(n_646), .B2(n_583), .C(n_578), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_672), .A2(n_561), .B(n_583), .C(n_578), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g759 ( .A1(n_679), .A2(n_583), .B(n_578), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_740), .A2(n_575), .B1(n_612), .B2(n_38), .Y(n_760) );
OAI221xp5_ASAP7_75t_SL g761 ( .A1(n_705), .A2(n_35), .B1(n_37), .B2(n_39), .C(n_40), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_675), .B(n_575), .Y(n_762) );
AO21x1_ASAP7_75t_L g763 ( .A1(n_713), .A2(n_37), .B(n_40), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_681), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_764) );
OAI221xp5_ASAP7_75t_SL g765 ( .A1(n_705), .A2(n_41), .B1(n_42), .B2(n_45), .C(n_46), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_722), .B(n_46), .Y(n_766) );
OAI211xp5_ASAP7_75t_SL g767 ( .A1(n_680), .A2(n_47), .B(n_48), .C(n_49), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_722), .B(n_47), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_650), .A2(n_48), .B(n_49), .C(n_50), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_681), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_770) );
NOR2xp67_ASAP7_75t_L g771 ( .A(n_656), .B(n_51), .Y(n_771) );
BUFx8_ASAP7_75t_SL g772 ( .A(n_667), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_709), .A2(n_54), .B1(n_55), .B2(n_58), .C(n_59), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g774 ( .A1(n_668), .A2(n_55), .B(n_59), .C(n_60), .Y(n_774) );
OAI211xp5_ASAP7_75t_SL g775 ( .A1(n_680), .A2(n_60), .B(n_61), .C(n_64), .Y(n_775) );
AOI322xp5_ASAP7_75t_L g776 ( .A1(n_720), .A2(n_61), .A3(n_65), .B1(n_66), .B2(n_110), .C1(n_111), .C2(n_112), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_744), .B(n_113), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_653), .A2(n_695), .B(n_651), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_684), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_726), .A2(n_117), .B1(n_119), .B2(n_120), .Y(n_780) );
AND2x4_ASAP7_75t_L g781 ( .A(n_661), .B(n_121), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_710), .B(n_124), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_697), .B(n_125), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_702), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_669), .B(n_126), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_719), .A2(n_127), .B1(n_129), .B2(n_131), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_730), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_664), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_788) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_745), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_730), .A2(n_138), .B1(n_140), .B2(n_144), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_662), .B(n_147), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_677), .A2(n_148), .B1(n_149), .B2(n_151), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_732), .A2(n_155), .B1(n_157), .B2(n_158), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_724), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_748), .A2(n_160), .B(n_162), .C(n_163), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_736), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_685), .A2(n_168), .B1(n_169), .B2(n_170), .C(n_172), .Y(n_797) );
OAI211xp5_ASAP7_75t_L g798 ( .A1(n_712), .A2(n_173), .B(n_177), .C(n_180), .Y(n_798) );
INVx4_ASAP7_75t_L g799 ( .A(n_664), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_660), .A2(n_181), .B1(n_183), .B2(n_191), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_664), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_661), .B(n_196), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_698), .A2(n_197), .B1(n_200), .B2(n_201), .C(n_202), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_679), .A2(n_203), .B1(n_209), .B2(n_210), .C(n_212), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_677), .A2(n_213), .B1(n_215), .B2(n_220), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_713), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_739), .Y(n_807) );
CKINVDCx6p67_ASAP7_75t_R g808 ( .A(n_676), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g809 ( .A(n_706), .Y(n_809) );
BUFx12f_ASAP7_75t_L g810 ( .A(n_711), .Y(n_810) );
INVx11_ASAP7_75t_L g811 ( .A(n_711), .Y(n_811) );
AO221x2_ASAP7_75t_L g812 ( .A1(n_728), .A2(n_224), .B1(n_225), .B2(n_226), .C(n_227), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_728), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_712), .A2(n_228), .B1(n_229), .B2(n_232), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_727), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_669), .B(n_238), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_727), .B(n_244), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_741), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_698), .A2(n_255), .B1(n_256), .B2(n_259), .C(n_261), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_699), .A2(n_262), .B(n_271), .Y(n_820) );
AO21x2_ASAP7_75t_L g821 ( .A1(n_729), .A2(n_655), .B(n_687), .Y(n_821) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_739), .A2(n_721), .B1(n_725), .B2(n_657), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_682), .A2(n_658), .B1(n_731), .B2(n_690), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_686), .A2(n_673), .B1(n_721), .B2(n_671), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_715), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_673), .A2(n_708), .B(n_674), .C(n_692), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_657), .A2(n_691), .B1(n_746), .B2(n_734), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_686), .A2(n_738), .B1(n_747), .B2(n_692), .Y(n_828) );
BUFx12f_ASAP7_75t_L g829 ( .A(n_649), .Y(n_829) );
BUFx4f_ASAP7_75t_SL g830 ( .A(n_689), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_733), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_714), .A2(n_723), .B1(n_670), .B2(n_663), .Y(n_832) );
AND2x4_ASAP7_75t_L g833 ( .A(n_723), .B(n_694), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_689), .B(n_693), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_693), .B(n_696), .Y(n_835) );
OA21x2_ASAP7_75t_L g836 ( .A1(n_665), .A2(n_666), .B(n_703), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_742), .A2(n_678), .B1(n_694), .B2(n_659), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_718), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_718), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_718), .Y(n_840) );
INVx1_ASAP7_75t_SL g841 ( .A(n_678), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_749), .A2(n_750), .B(n_704), .C(n_743), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_654), .A2(n_707), .B1(n_716), .B2(n_717), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_735), .B(n_737), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_700), .A2(n_594), .B1(n_719), .B2(n_467), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_719), .A2(n_594), .B1(n_467), .B2(n_584), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_818), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_829), .Y(n_848) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_833), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_813), .B(n_796), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_784), .Y(n_851) );
INVx2_ASAP7_75t_SL g852 ( .A(n_755), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_806), .B(n_846), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_779), .Y(n_854) );
AND2x4_ASAP7_75t_SL g855 ( .A(n_789), .B(n_808), .Y(n_855) );
CKINVDCx11_ASAP7_75t_R g856 ( .A(n_789), .Y(n_856) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_771), .B(n_799), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_835), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_766), .B(n_768), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_799), .B(n_841), .Y(n_860) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_807), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_836), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_825), .B(n_831), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_836), .Y(n_864) );
INVx4_ASAP7_75t_L g865 ( .A(n_830), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_835), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_820), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_809), .B(n_756), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_777), .B(n_812), .Y(n_869) );
OAI222xp33_ASAP7_75t_L g870 ( .A1(n_822), .A2(n_845), .B1(n_761), .B2(n_765), .C1(n_752), .C2(n_819), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_838), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_839), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_841), .B(n_781), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_812), .B(n_763), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_753), .B(n_823), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_840), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_794), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_781), .Y(n_878) );
INVx3_ASAP7_75t_L g879 ( .A(n_802), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_802), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_782), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_827), .B(n_791), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_754), .B(n_783), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_844), .Y(n_884) );
OR2x6_ASAP7_75t_L g885 ( .A(n_792), .B(n_805), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_821), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_783), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_834), .B(n_824), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_834), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_754), .B(n_828), .Y(n_890) );
BUFx3_ASAP7_75t_L g891 ( .A(n_810), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_821), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_824), .B(n_776), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_778), .Y(n_894) );
NOR2x1_ASAP7_75t_L g895 ( .A(n_792), .B(n_805), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_755), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_843), .Y(n_897) );
AND2x4_ASAP7_75t_L g898 ( .A(n_758), .B(n_762), .Y(n_898) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_785), .Y(n_899) );
INVx2_ASAP7_75t_SL g900 ( .A(n_789), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_816), .B(n_826), .Y(n_901) );
BUFx3_ASAP7_75t_L g902 ( .A(n_751), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_759), .B(n_760), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_817), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_769), .B(n_774), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_842), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_764), .B(n_770), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_795), .B(n_800), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_832), .Y(n_909) );
AND2x4_ASAP7_75t_L g910 ( .A(n_787), .B(n_790), .Y(n_910) );
NOR2x1_ASAP7_75t_L g911 ( .A(n_767), .B(n_775), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_803), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_773), .B(n_786), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_797), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_798), .Y(n_915) );
INVx2_ASAP7_75t_SL g916 ( .A(n_811), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_814), .B(n_757), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_788), .Y(n_918) );
INVx2_ASAP7_75t_SL g919 ( .A(n_837), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_815), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_804), .B(n_780), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_801), .B(n_793), .Y(n_922) );
OR2x6_ASAP7_75t_L g923 ( .A(n_772), .B(n_681), .Y(n_923) );
OAI31xp33_ASAP7_75t_L g924 ( .A1(n_870), .A2(n_893), .A3(n_869), .B(n_875), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_923), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_858), .B(n_866), .Y(n_926) );
INVx4_ASAP7_75t_L g927 ( .A(n_878), .Y(n_927) );
INVxp67_ASAP7_75t_SL g928 ( .A(n_880), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_890), .B(n_858), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_890), .B(n_866), .Y(n_930) );
NAND2x1_ASAP7_75t_L g931 ( .A(n_878), .B(n_879), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_871), .Y(n_932) );
BUFx3_ASAP7_75t_L g933 ( .A(n_848), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_883), .B(n_884), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_862), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_888), .B(n_853), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_871), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_888), .B(n_850), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_884), .B(n_889), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_862), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_889), .B(n_859), .Y(n_941) );
OAI21x1_ASAP7_75t_SL g942 ( .A1(n_895), .A2(n_857), .B(n_918), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_883), .B(n_847), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_864), .Y(n_944) );
INVx5_ASAP7_75t_L g945 ( .A(n_878), .Y(n_945) );
BUFx6f_ASAP7_75t_SL g946 ( .A(n_923), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_872), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_864), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_859), .B(n_854), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g950 ( .A1(n_893), .A2(n_869), .B1(n_874), .B2(n_907), .C1(n_882), .C2(n_913), .Y(n_950) );
CKINVDCx16_ASAP7_75t_R g951 ( .A(n_923), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_851), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_894), .Y(n_953) );
OAI31xp33_ASAP7_75t_L g954 ( .A1(n_913), .A2(n_874), .A3(n_907), .B(n_918), .Y(n_954) );
BUFx3_ASAP7_75t_L g955 ( .A(n_848), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g956 ( .A(n_911), .B(n_894), .C(n_895), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_851), .B(n_863), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_876), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_877), .B(n_896), .Y(n_959) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_879), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_906), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g962 ( .A(n_905), .B(n_909), .C(n_904), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_861), .A2(n_852), .B(n_868), .C(n_909), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_852), .B(n_916), .Y(n_964) );
INVx3_ASAP7_75t_L g965 ( .A(n_873), .Y(n_965) );
BUFx3_ASAP7_75t_L g966 ( .A(n_848), .Y(n_966) );
OAI21xp5_ASAP7_75t_L g967 ( .A1(n_914), .A2(n_921), .B(n_917), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_849), .B(n_860), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_914), .A2(n_885), .B1(n_915), .B2(n_920), .C(n_900), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_910), .A2(n_912), .B1(n_908), .B2(n_922), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_860), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_881), .B(n_887), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_881), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_887), .B(n_901), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_897), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_901), .B(n_849), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_936), .B(n_903), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_958), .Y(n_978) );
NOR2xp67_ASAP7_75t_L g979 ( .A(n_963), .B(n_900), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_964), .B(n_891), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_934), .B(n_886), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_936), .B(n_903), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_935), .Y(n_983) );
AND2x2_ASAP7_75t_SL g984 ( .A(n_951), .B(n_855), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_934), .B(n_892), .Y(n_985) );
INVx1_ASAP7_75t_SL g986 ( .A(n_933), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_938), .B(n_892), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_957), .B(n_919), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_929), .B(n_886), .Y(n_989) );
BUFx2_ASAP7_75t_L g990 ( .A(n_971), .Y(n_990) );
NOR2xp67_ASAP7_75t_L g991 ( .A(n_925), .B(n_865), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_924), .A2(n_902), .B1(n_865), .B2(n_915), .C(n_891), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_940), .Y(n_993) );
INVxp67_ASAP7_75t_L g994 ( .A(n_959), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_940), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_930), .B(n_899), .Y(n_996) );
INVx1_ASAP7_75t_SL g997 ( .A(n_933), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_930), .B(n_899), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_944), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_944), .Y(n_1000) );
NOR2x1_ASAP7_75t_L g1001 ( .A(n_955), .B(n_898), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_943), .B(n_899), .Y(n_1002) );
NAND2x1p5_ASAP7_75t_L g1003 ( .A(n_945), .B(n_898), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_932), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_932), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_968), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_948), .Y(n_1007) );
INVx3_ASAP7_75t_L g1008 ( .A(n_927), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_974), .B(n_867), .Y(n_1009) );
NOR3xp33_ASAP7_75t_L g1010 ( .A(n_956), .B(n_856), .C(n_922), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_948), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_937), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_947), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_947), .Y(n_1014) );
INVx1_ASAP7_75t_SL g1015 ( .A(n_955), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g1016 ( .A(n_962), .B(n_954), .C(n_967), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_949), .B(n_941), .Y(n_1017) );
NAND2xp33_ASAP7_75t_L g1018 ( .A(n_1010), .B(n_925), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_990), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_1017), .B(n_926), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1004), .Y(n_1021) );
NAND4xp25_ASAP7_75t_L g1022 ( .A(n_1016), .B(n_950), .C(n_970), .D(n_969), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1004), .Y(n_1023) );
NOR2x1_ASAP7_75t_L g1024 ( .A(n_991), .B(n_966), .Y(n_1024) );
NAND2x1_ASAP7_75t_L g1025 ( .A(n_1008), .B(n_942), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1005), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_988), .B(n_952), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1012), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_992), .B(n_928), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_977), .B(n_982), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_990), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_983), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_983), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1013), .Y(n_1034) );
INVx3_ASAP7_75t_L g1035 ( .A(n_1008), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1002), .B(n_953), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_994), .B(n_946), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_987), .B(n_939), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1014), .Y(n_1039) );
NOR2xp67_ASAP7_75t_SL g1040 ( .A(n_1035), .B(n_1008), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1030), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1020), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1019), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_1022), .A2(n_979), .B(n_984), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1021), .Y(n_1045) );
AOI21xp33_ASAP7_75t_L g1046 ( .A1(n_1029), .A2(n_980), .B(n_942), .Y(n_1046) );
AOI21xp33_ASAP7_75t_L g1047 ( .A1(n_1029), .A2(n_1001), .B(n_997), .Y(n_1047) );
OAI21xp5_ASAP7_75t_L g1048 ( .A1(n_1018), .A2(n_1003), .B(n_960), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1023), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1025), .A2(n_986), .B1(n_1015), .B2(n_1006), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_1038), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1026), .Y(n_1052) );
AOI32xp33_ASAP7_75t_L g1053 ( .A1(n_1037), .A2(n_1002), .A3(n_996), .B1(n_998), .B2(n_989), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1045), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1049), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1056 ( .A(n_1046), .B(n_1041), .Y(n_1056) );
AOI21xp5_ASAP7_75t_L g1057 ( .A1(n_1048), .A2(n_1024), .B(n_1035), .Y(n_1057) );
OA22x2_ASAP7_75t_L g1058 ( .A1(n_1044), .A2(n_1035), .B1(n_1031), .B2(n_1027), .Y(n_1058) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_1043), .Y(n_1059) );
NAND2xp5_ASAP7_75t_SL g1060 ( .A(n_1050), .B(n_1032), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1052), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1051), .B(n_1036), .Y(n_1062) );
OAI211xp5_ASAP7_75t_L g1063 ( .A1(n_1048), .A2(n_1039), .B(n_1028), .C(n_1034), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1042), .Y(n_1064) );
NAND5xp2_ASAP7_75t_L g1065 ( .A(n_1057), .B(n_1056), .C(n_1063), .D(n_1047), .E(n_1053), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1054), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1067 ( .A1(n_1058), .A2(n_945), .B1(n_931), .B2(n_1040), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1055), .Y(n_1068) );
OAI211xp5_ASAP7_75t_SL g1069 ( .A1(n_1060), .A2(n_965), .B(n_976), .C(n_961), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_1065), .A2(n_1064), .B1(n_1061), .B2(n_1059), .C(n_1062), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_1069), .A2(n_1067), .B1(n_1068), .B2(n_1066), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_1071), .B(n_1033), .Y(n_1072) );
NAND5xp2_ASAP7_75t_L g1073 ( .A(n_1070), .B(n_972), .C(n_973), .D(n_1009), .E(n_985), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_1072), .Y(n_1074) );
NOR2x1_ASAP7_75t_L g1075 ( .A(n_1073), .B(n_978), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1076 ( .A(n_1074), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_1076), .A2(n_1075), .B(n_953), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1077), .Y(n_1078) );
AOI222xp33_ASAP7_75t_SL g1079 ( .A1(n_1078), .A2(n_1007), .B1(n_1000), .B2(n_999), .C1(n_995), .C2(n_993), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_1079), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g1081 ( .A1(n_1080), .A2(n_975), .B1(n_981), .B2(n_999), .C1(n_995), .C2(n_1011), .Y(n_1081) );
endmodule