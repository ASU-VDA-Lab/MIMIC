module fake_jpeg_17367_n_58 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_3),
.B1(n_0),
.B2(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_1),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_37),
.B(n_4),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.C(n_41),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_10),
.C(n_14),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_4),
.B(n_5),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_32),
.B(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.C(n_36),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_32),
.Y(n_47)
);

XOR2x1_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_33),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_46),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_46),
.C(n_47),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.B(n_7),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_6),
.B(n_7),
.Y(n_58)
);


endmodule