module real_jpeg_5942_n_17 (n_8, n_116, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_117, n_3, n_5, n_4, n_109, n_115, n_1, n_118, n_16, n_15, n_13, n_113, n_17);

input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_117;
input n_3;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_0),
.B(n_81),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_2),
.B(n_46),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_4),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_6),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_6),
.B(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_8),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_31),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_16),
.B(n_35),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_27),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_74),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_50),
.B(n_100),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR4xp25_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_40),
.D(n_45),
.Y(n_29)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_39),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_96),
.B(n_99),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_88),
.B(n_95),
.Y(n_52)
);

AO221x1_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_65),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_84),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_69),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_83),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_79),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_94),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_105),
.C(n_106),
.D(n_107),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_109),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_110),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_111),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_112),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_113),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_114),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_115),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_116),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_117),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_118),
.Y(n_98)
);


endmodule