module real_aes_6498_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_729;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g550 ( .A1(n_0), .A2(n_155), .B(n_551), .C(n_554), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_1), .B(n_495), .Y(n_555) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g189 ( .A(n_3), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_4), .B(n_147), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_5), .A2(n_464), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_6), .A2(n_132), .B(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_7), .A2(n_36), .B1(n_141), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_8), .B(n_132), .Y(n_158) );
AND2x6_ASAP7_75t_L g156 ( .A(n_9), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_10), .A2(n_156), .B(n_454), .C(n_456), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_11), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_11), .B(n_37), .Y(n_440) );
INVx1_ASAP7_75t_L g137 ( .A(n_12), .Y(n_137) );
INVx1_ASAP7_75t_L g182 ( .A(n_13), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_14), .B(n_145), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_15), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_16), .B(n_147), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_17), .B(n_133), .Y(n_194) );
AO32x2_ASAP7_75t_L g216 ( .A1(n_18), .A2(n_132), .A3(n_162), .B1(n_173), .B2(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_19), .B(n_141), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_20), .B(n_133), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_21), .A2(n_54), .B1(n_141), .B2(n_219), .Y(n_220) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_22), .A2(n_81), .B1(n_141), .B2(n_145), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_23), .B(n_141), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_24), .A2(n_173), .B(n_454), .C(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_25), .A2(n_173), .B(n_454), .C(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_26), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_27), .B(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_28), .A2(n_464), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_29), .B(n_175), .Y(n_213) );
INVx2_ASAP7_75t_L g143 ( .A(n_30), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_31), .A2(n_466), .B(n_474), .C(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_32), .A2(n_103), .B1(n_115), .B2(n_759), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_33), .B(n_141), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_34), .B(n_175), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_35), .B(n_227), .Y(n_484) );
INVx1_ASAP7_75t_L g114 ( .A(n_37), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_38), .B(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_39), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_40), .A2(n_78), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_40), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_41), .B(n_147), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_42), .B(n_464), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_43), .A2(n_79), .B1(n_435), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_43), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_44), .A2(n_466), .B(n_468), .C(n_474), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_45), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g552 ( .A(n_46), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_47), .A2(n_90), .B1(n_219), .B2(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g469 ( .A(n_48), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_49), .B(n_141), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_50), .B(n_141), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_51), .B(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_51), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_52), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_53), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_SL g198 ( .A1(n_55), .A2(n_59), .B1(n_141), .B2(n_145), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_56), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_57), .B(n_141), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_58), .B(n_141), .Y(n_224) );
INVx1_ASAP7_75t_L g157 ( .A(n_60), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_61), .B(n_464), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_62), .B(n_495), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_63), .A2(n_153), .B(n_185), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_64), .B(n_141), .Y(n_190) );
INVx1_ASAP7_75t_L g136 ( .A(n_65), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_66), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_67), .B(n_147), .Y(n_505) );
AO32x2_ASAP7_75t_L g237 ( .A1(n_68), .A2(n_132), .A3(n_173), .B1(n_238), .B2(n_242), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_69), .B(n_148), .Y(n_457) );
INVx1_ASAP7_75t_L g168 ( .A(n_70), .Y(n_168) );
INVx1_ASAP7_75t_L g208 ( .A(n_71), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_72), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_73), .B(n_471), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_74), .A2(n_454), .B(n_474), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_75), .B(n_145), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_76), .Y(n_490) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_78), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_79), .A2(n_124), .B1(n_434), .B2(n_435), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_79), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_80), .B(n_470), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_82), .B(n_219), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_83), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_84), .B(n_145), .Y(n_212) );
INVx2_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_86), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_87), .B(n_172), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_88), .B(n_145), .Y(n_144) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_89), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g438 ( .A(n_89), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g728 ( .A(n_89), .Y(n_728) );
OR2x2_ASAP7_75t_L g752 ( .A(n_89), .B(n_738), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_91), .A2(n_101), .B1(n_145), .B2(n_146), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_92), .B(n_464), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_93), .Y(n_735) );
INVx1_ASAP7_75t_L g504 ( .A(n_94), .Y(n_504) );
INVxp67_ASAP7_75t_L g493 ( .A(n_95), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_96), .B(n_145), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g450 ( .A(n_98), .Y(n_450) );
INVx1_ASAP7_75t_L g528 ( .A(n_99), .Y(n_528) );
AND2x2_ASAP7_75t_L g476 ( .A(n_100), .B(n_175), .Y(n_476) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g439 ( .A(n_108), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_739), .B1(n_742), .B2(n_753), .C(n_755), .Y(n_115) );
OAI222xp33_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_120), .B1(n_729), .B2(n_730), .C1(n_735), .C2(n_736), .Y(n_116) );
INVx1_ASAP7_75t_L g729 ( .A(n_117), .Y(n_729) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_436), .B1(n_441), .B2(n_725), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_123), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g434 ( .A(n_124), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_124), .A2(n_434), .B1(n_745), .B2(n_746), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_125), .B(n_358), .Y(n_124) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_316), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_256), .C(n_292), .D(n_306), .Y(n_126) );
OAI221xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_200), .B1(n_232), .B2(n_243), .C(n_247), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_128), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_176), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_159), .Y(n_130) );
AND2x2_ASAP7_75t_L g253 ( .A(n_131), .B(n_160), .Y(n_253) );
INVx3_ASAP7_75t_L g261 ( .A(n_131), .Y(n_261) );
AND2x2_ASAP7_75t_L g315 ( .A(n_131), .B(n_179), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_131), .B(n_178), .Y(n_351) );
AND2x2_ASAP7_75t_L g409 ( .A(n_131), .B(n_271), .Y(n_409) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_138), .B(n_158), .Y(n_131) );
INVx4_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_132), .A2(n_481), .B(n_482), .Y(n_480) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_132), .Y(n_487) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_134), .B(n_135), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_150), .B(n_156), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_144), .B(n_147), .Y(n_139) );
INVx3_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_141), .Y(n_530) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
BUFx3_ASAP7_75t_L g240 ( .A(n_142), .Y(n_240) );
AND2x6_ASAP7_75t_L g454 ( .A(n_142), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
INVx2_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_147), .A2(n_165), .B(n_166), .Y(n_164) );
O2A1O1Ixp5_ASAP7_75t_SL g206 ( .A1(n_147), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_147), .B(n_493), .Y(n_492) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_148), .A2(n_172), .B1(n_239), .B2(n_241), .Y(n_238) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
AND2x2_ASAP7_75t_L g452 ( .A(n_149), .B(n_154), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_149), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .Y(n_150) );
INVx2_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_169), .B(n_189), .C(n_190), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_155), .A2(n_172), .B1(n_197), .B2(n_198), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_155), .A2(n_172), .B1(n_218), .B2(n_220), .Y(n_217) );
BUFx3_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_156), .A2(n_181), .B(n_188), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_156), .A2(n_206), .B(n_210), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_156), .A2(n_223), .B(n_228), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_156), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g464 ( .A(n_156), .B(n_452), .Y(n_464) );
INVx4_ASAP7_75t_SL g475 ( .A(n_156), .Y(n_475) );
AND2x2_ASAP7_75t_L g244 ( .A(n_159), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g258 ( .A(n_159), .B(n_179), .Y(n_258) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_160), .B(n_179), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_160), .B(n_261), .Y(n_285) );
OR2x2_ASAP7_75t_L g287 ( .A(n_160), .B(n_245), .Y(n_287) );
AND2x2_ASAP7_75t_L g322 ( .A(n_160), .B(n_245), .Y(n_322) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_160), .Y(n_367) );
INVx1_ASAP7_75t_L g375 ( .A(n_160), .Y(n_375) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_174), .Y(n_160) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_161), .A2(n_180), .B(n_191), .Y(n_179) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_162), .B(n_460), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_173), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_171), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_169), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g553 ( .A(n_172), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_173), .B(n_196), .C(n_199), .Y(n_195) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_175), .A2(n_205), .B(n_213), .Y(n_204) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_222), .B(n_231), .Y(n_221) );
INVx2_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_175), .A2(n_463), .B(n_465), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_175), .A2(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g521 ( .A(n_175), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_176), .A2(n_293), .B1(n_297), .B2(n_301), .C(n_302), .Y(n_292) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g252 ( .A(n_177), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_192), .Y(n_177) );
INVx2_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
AND2x2_ASAP7_75t_L g304 ( .A(n_178), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g323 ( .A(n_178), .B(n_261), .Y(n_323) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g386 ( .A(n_179), .B(n_261), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_185), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_183), .A2(n_457), .B(n_458), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_183), .A2(n_484), .B(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_185), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_186), .A2(n_211), .B(n_212), .Y(n_210) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g471 ( .A(n_187), .Y(n_471) );
AND2x2_ASAP7_75t_L g308 ( .A(n_192), .B(n_253), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g376 ( .A1(n_192), .A2(n_332), .A3(n_377), .B1(n_379), .B2(n_382), .C1(n_384), .C2(n_388), .Y(n_376) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_193), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g272 ( .A(n_193), .Y(n_272) );
AND2x2_ASAP7_75t_L g381 ( .A(n_193), .B(n_261), .Y(n_381) );
AND2x2_ASAP7_75t_L g413 ( .A(n_193), .B(n_285), .Y(n_413) );
OR2x2_ASAP7_75t_L g416 ( .A(n_193), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g246 ( .A(n_194), .Y(n_246) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_196), .A2(n_199), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_199), .A2(n_449), .B(n_459), .Y(n_448) );
INVx3_ASAP7_75t_L g495 ( .A(n_199), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_199), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_199), .A2(n_525), .B(n_532), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_199), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_214), .Y(n_201) );
INVx1_ASAP7_75t_L g429 ( .A(n_202), .Y(n_429) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g234 ( .A(n_203), .B(n_221), .Y(n_234) );
INVx2_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g291 ( .A(n_204), .Y(n_291) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_204), .Y(n_299) );
OR2x2_ASAP7_75t_L g423 ( .A(n_204), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g248 ( .A(n_214), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g288 ( .A(n_214), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g340 ( .A(n_214), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
AND2x2_ASAP7_75t_L g235 ( .A(n_215), .B(n_236), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_215), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g349 ( .A(n_215), .B(n_237), .Y(n_349) );
OR2x2_ASAP7_75t_L g357 ( .A(n_215), .B(n_291), .Y(n_357) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g266 ( .A(n_216), .Y(n_266) );
AND2x2_ASAP7_75t_L g276 ( .A(n_216), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g300 ( .A(n_216), .B(n_221), .Y(n_300) );
AND2x2_ASAP7_75t_L g364 ( .A(n_216), .B(n_237), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_221), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_221), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
INVx1_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
AND2x2_ASAP7_75t_L g294 ( .A(n_221), .B(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_221), .Y(n_372) );
INVx1_ASAP7_75t_L g424 ( .A(n_221), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g401 ( .A(n_233), .B(n_310), .Y(n_401) );
INVx2_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g328 ( .A(n_235), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g427 ( .A(n_235), .B(n_362), .Y(n_427) );
INVx1_ASAP7_75t_L g249 ( .A(n_236), .Y(n_249) );
AND2x2_ASAP7_75t_L g275 ( .A(n_236), .B(n_269), .Y(n_275) );
BUFx2_ASAP7_75t_L g334 ( .A(n_236), .Y(n_334) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_237), .Y(n_255) );
INVx1_ASAP7_75t_L g265 ( .A(n_237), .Y(n_265) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_240), .Y(n_473) );
INVx2_ASAP7_75t_L g554 ( .A(n_240), .Y(n_554) );
INVx1_ASAP7_75t_L g518 ( .A(n_242), .Y(n_518) );
NOR2xp67_ASAP7_75t_L g403 ( .A(n_243), .B(n_250), .Y(n_403) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI32xp33_ASAP7_75t_L g247 ( .A1(n_244), .A2(n_248), .A3(n_250), .B1(n_252), .B2(n_254), .Y(n_247) );
AND2x2_ASAP7_75t_L g387 ( .A(n_244), .B(n_260), .Y(n_387) );
AND2x2_ASAP7_75t_L g425 ( .A(n_244), .B(n_323), .Y(n_425) );
INVx1_ASAP7_75t_L g305 ( .A(n_245), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_249), .B(n_311), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_250), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_250), .B(n_253), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_250), .B(n_322), .Y(n_404) );
OR2x2_ASAP7_75t_L g418 ( .A(n_250), .B(n_287), .Y(n_418) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g345 ( .A(n_251), .B(n_253), .Y(n_345) );
OR2x2_ASAP7_75t_L g354 ( .A(n_251), .B(n_341), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_253), .B(n_304), .Y(n_326) );
INVx2_ASAP7_75t_L g341 ( .A(n_255), .Y(n_341) );
OR2x2_ASAP7_75t_L g356 ( .A(n_255), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g371 ( .A(n_255), .B(n_372), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g428 ( .A1(n_255), .A2(n_348), .B(n_429), .C(n_430), .Y(n_428) );
OAI321xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .A3(n_267), .B1(n_270), .B2(n_274), .C(n_278), .Y(n_256) );
INVx1_ASAP7_75t_L g369 ( .A(n_257), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g380 ( .A(n_258), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g332 ( .A(n_260), .Y(n_332) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_261), .B(n_375), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_262), .A2(n_400), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x2_ASAP7_75t_L g337 ( .A(n_264), .B(n_311), .Y(n_337) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_265), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_267), .A2(n_308), .B(n_353), .C(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g319 ( .A(n_269), .B(n_276), .Y(n_319) );
BUFx2_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
INVx1_ASAP7_75t_L g344 ( .A(n_269), .Y(n_344) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OR2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g433 ( .A(n_272), .Y(n_433) );
INVx1_ASAP7_75t_L g426 ( .A(n_273), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g383 ( .A(n_275), .B(n_300), .Y(n_383) );
INVx1_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_283), .B1(n_286), .B2(n_288), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_280), .B(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g348 ( .A(n_281), .B(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_282), .B(n_291), .Y(n_311) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g303 ( .A(n_285), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g313 ( .A(n_287), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_290), .A2(n_408), .B1(n_410), .B2(n_411), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g296 ( .A(n_291), .Y(n_296) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_291), .Y(n_362) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_294), .B(n_413), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_295), .A2(n_300), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_298), .B(n_308), .Y(n_405) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g374 ( .A(n_299), .Y(n_374) );
AND2x2_ASAP7_75t_L g333 ( .A(n_300), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g422 ( .A(n_300), .Y(n_422) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g393 ( .A(n_304), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_312), .B2(n_313), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_310), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g378 ( .A(n_311), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_311), .B(n_349), .Y(n_415) );
OR2x2_ASAP7_75t_L g388 ( .A(n_312), .B(n_341), .Y(n_388) );
INVx1_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_315), .B(n_366), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_335), .C(n_346), .Y(n_316) );
OAI211xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B(n_324), .C(n_330), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_319), .A2(n_390), .B1(n_394), .B2(n_397), .C(n_399), .Y(n_389) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g385 ( .A(n_322), .B(n_386), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_323), .A2(n_371), .B(n_373), .C(n_375), .Y(n_370) );
INVx2_ASAP7_75t_L g417 ( .A(n_323), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_327), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g396 ( .A(n_329), .B(n_349), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
OAI21xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_338), .B(n_339), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI21xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_342), .B(n_345), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_340), .B(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_345), .B(n_432), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B(n_352), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g373 ( .A(n_349), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND4x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_389), .C(n_406), .D(n_428), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_376), .Y(n_359) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_365), .B(n_368), .C(n_370), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_364), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_375), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g410 ( .A(n_385), .Y(n_410) );
INVx2_ASAP7_75t_SL g398 ( .A(n_386), .Y(n_398) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g411 ( .A(n_396), .Y(n_411) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_414), .Y(n_406) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B1(n_418), .B2(n_419), .C(n_420), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g732 ( .A(n_437), .Y(n_732) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g727 ( .A(n_439), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g738 ( .A(n_439), .Y(n_738) );
INVx2_ASAP7_75t_L g733 ( .A(n_441), .Y(n_733) );
OR3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_623), .C(n_688), .Y(n_441) );
NAND4xp25_ASAP7_75t_SL g442 ( .A(n_443), .B(n_564), .C(n_590), .D(n_613), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_496), .B1(n_534), .B2(n_541), .C(n_556), .Y(n_443) );
CKINVDCx14_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_445), .A2(n_557), .B1(n_581), .B2(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_477), .Y(n_445) );
INVx1_ASAP7_75t_SL g617 ( .A(n_446), .Y(n_617) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_461), .Y(n_446) );
OR2x2_ASAP7_75t_L g539 ( .A(n_447), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g559 ( .A(n_447), .B(n_478), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_447), .B(n_486), .Y(n_572) );
AND2x2_ASAP7_75t_L g589 ( .A(n_447), .B(n_461), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_447), .B(n_537), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_447), .B(n_588), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_447), .B(n_477), .Y(n_710) );
AOI211xp5_ASAP7_75t_SL g721 ( .A1(n_447), .A2(n_627), .B(n_722), .C(n_723), .Y(n_721) );
INVx5_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_448), .B(n_478), .Y(n_593) );
AND2x2_ASAP7_75t_L g596 ( .A(n_448), .B(n_479), .Y(n_596) );
OR2x2_ASAP7_75t_L g641 ( .A(n_448), .B(n_478), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_448), .B(n_486), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_453), .Y(n_449) );
INVx5_ASAP7_75t_L g467 ( .A(n_454), .Y(n_467) );
INVx5_ASAP7_75t_SL g540 ( .A(n_461), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_461), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_461), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g644 ( .A(n_461), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g676 ( .A(n_461), .B(n_486), .Y(n_676) );
OR2x2_ASAP7_75t_L g682 ( .A(n_461), .B(n_572), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_461), .B(n_632), .Y(n_691) );
OR2x6_ASAP7_75t_L g461 ( .A(n_462), .B(n_476), .Y(n_461) );
BUFx2_ASAP7_75t_L g513 ( .A(n_464), .Y(n_513) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_467), .A2(n_475), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g548 ( .A1(n_467), .A2(n_475), .B(n_549), .C(n_550), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_472), .C(n_473), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_470), .A2(n_473), .B(n_504), .C(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
AND2x2_ASAP7_75t_L g573 ( .A(n_478), .B(n_540), .Y(n_573) );
INVx1_ASAP7_75t_SL g586 ( .A(n_478), .Y(n_586) );
OR2x2_ASAP7_75t_L g621 ( .A(n_478), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g627 ( .A(n_478), .B(n_486), .Y(n_627) );
AND2x2_ASAP7_75t_L g685 ( .A(n_478), .B(n_537), .Y(n_685) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_479), .B(n_540), .Y(n_612) );
INVx3_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
OR2x2_ASAP7_75t_L g578 ( .A(n_486), .B(n_540), .Y(n_578) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_586), .Y(n_588) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_486), .Y(n_636) );
AND2x2_ASAP7_75t_L g645 ( .A(n_486), .B(n_559), .Y(n_645) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_494), .Y(n_486) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_495), .A2(n_547), .B(n_555), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_496), .A2(n_662), .B1(n_664), .B2(n_666), .C(n_669), .Y(n_661) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
AND2x2_ASAP7_75t_L g635 ( .A(n_498), .B(n_616), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_498), .B(n_694), .Y(n_698) );
OR2x2_ASAP7_75t_L g719 ( .A(n_498), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_498), .B(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
AND2x2_ASAP7_75t_L g643 ( .A(n_499), .B(n_510), .Y(n_643) );
AND2x2_ASAP7_75t_L g704 ( .A(n_499), .B(n_583), .Y(n_704) );
AND2x2_ASAP7_75t_L g717 ( .A(n_499), .B(n_537), .Y(n_717) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_522), .Y(n_508) );
AND2x4_ASAP7_75t_L g544 ( .A(n_509), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g562 ( .A(n_509), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g569 ( .A(n_509), .Y(n_569) );
AND2x2_ASAP7_75t_L g638 ( .A(n_509), .B(n_616), .Y(n_638) );
AND2x2_ASAP7_75t_L g648 ( .A(n_509), .B(n_566), .Y(n_648) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_509), .Y(n_656) );
AND2x2_ASAP7_75t_L g668 ( .A(n_509), .B(n_546), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_509), .B(n_600), .Y(n_672) );
AND2x2_ASAP7_75t_L g709 ( .A(n_509), .B(n_704), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_509), .B(n_583), .Y(n_720) );
OR2x2_ASAP7_75t_L g722 ( .A(n_509), .B(n_658), .Y(n_722) );
INVx5_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g608 ( .A(n_510), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g618 ( .A(n_510), .B(n_563), .Y(n_618) );
AND2x2_ASAP7_75t_L g630 ( .A(n_510), .B(n_546), .Y(n_630) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_510), .Y(n_660) );
AND2x4_ASAP7_75t_L g694 ( .A(n_510), .B(n_545), .Y(n_694) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
AOI21xp5_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_514), .B(n_518), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
BUFx2_ASAP7_75t_L g543 ( .A(n_522), .Y(n_543) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_523), .B(n_546), .Y(n_616) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g563 ( .A(n_524), .B(n_546), .Y(n_563) );
BUFx2_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .Y(n_525) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_536), .B(n_617), .Y(n_696) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_537), .B(n_559), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_537), .B(n_540), .Y(n_598) );
AND2x2_ASAP7_75t_L g653 ( .A(n_537), .B(n_589), .Y(n_653) );
AOI221xp5_ASAP7_75t_SL g590 ( .A1(n_538), .A2(n_591), .B1(n_599), .B2(n_601), .C(n_605), .Y(n_590) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g585 ( .A(n_539), .B(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g626 ( .A(n_539), .B(n_627), .Y(n_626) );
OAI321xp33_ASAP7_75t_L g633 ( .A1(n_539), .A2(n_592), .A3(n_634), .B1(n_636), .B2(n_637), .C(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_540), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_543), .B(n_694), .Y(n_712) );
AND2x2_ASAP7_75t_L g599 ( .A(n_544), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_544), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_545), .Y(n_575) );
AND2x2_ASAP7_75t_L g582 ( .A(n_545), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_545), .B(n_657), .Y(n_687) );
INVx1_ASAP7_75t_L g724 ( .A(n_545), .Y(n_724) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_561), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_558), .A2(n_668), .B(n_717), .C(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_559), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_559), .B(n_597), .Y(n_663) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_563), .B(n_566), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_563), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_563), .B(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B1(n_579), .B2(n_584), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g580 ( .A(n_566), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g603 ( .A(n_566), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g615 ( .A(n_566), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_566), .B(n_609), .Y(n_651) );
OR2x2_ASAP7_75t_L g658 ( .A(n_566), .B(n_583), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_566), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g708 ( .A(n_566), .B(n_694), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B1(n_574), .B2(n_576), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g614 ( .A(n_569), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_572), .A2(n_587), .B1(n_655), .B2(n_659), .Y(n_654) );
INVx1_ASAP7_75t_L g702 ( .A(n_573), .Y(n_702) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_614), .B1(n_617), .B2(n_618), .C(n_619), .Y(n_613) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g592 ( .A(n_578), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_582), .B(n_648), .Y(n_680) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_583), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_583), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g622 ( .A(n_589), .Y(n_622) );
AND2x2_ASAP7_75t_L g631 ( .A(n_589), .B(n_632), .Y(n_631) );
NAND2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g675 ( .A(n_596), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_599), .A2(n_625), .B1(n_628), .B2(n_631), .C(n_633), .Y(n_624) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_603), .B(n_660), .Y(n_659) );
AOI21xp33_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_607), .B(n_610), .Y(n_605) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
CKINVDCx16_ASAP7_75t_R g707 ( .A(n_610), .Y(n_707) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
OR2x2_ASAP7_75t_L g649 ( .A(n_612), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g670 ( .A(n_615), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_615), .B(n_675), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_618), .B(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_642), .C(n_661), .D(n_674), .Y(n_623) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g632 ( .A(n_627), .Y(n_632) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g665 ( .A(n_636), .B(n_641), .Y(n_665) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_646), .C(n_654), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_644), .A2(n_686), .B(n_714), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_SL g673 ( .A(n_645), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_651), .B2(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g677 ( .A(n_651), .Y(n_677) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_657), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_657), .B(n_668), .Y(n_701) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g678 ( .A(n_668), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B(n_673), .Y(n_669) );
INVxp33_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .A3(n_678), .B1(n_679), .B2(n_681), .C1(n_683), .C2(n_686), .Y(n_674) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g688 ( .A(n_689), .B(n_706), .C(n_713), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B1(n_695), .B2(n_697), .C(n_699), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g705 ( .A(n_694), .Y(n_705) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_709), .B2(n_710), .C(n_711), .Y(n_706) );
NAND2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g734 ( .A(n_726), .Y(n_734) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_728), .B(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g754 ( .A(n_740), .Y(n_754) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_748), .C(n_751), .Y(n_742) );
INVx1_ASAP7_75t_L g750 ( .A(n_744), .Y(n_750) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g758 ( .A(n_752), .Y(n_758) );
BUFx3_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule