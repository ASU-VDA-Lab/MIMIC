module fake_aes_9115_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
OR2x2_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_3), .Y(n_7) );
AOI222xp33_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_0), .B1(n_1), .B2(n_2), .C1(n_4), .C2(n_3), .Y(n_8) );
OAI22xp33_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_9) );
AOI221xp5_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_7), .B1(n_8), .B2(n_1), .C(n_2), .Y(n_10) );
NAND2x1p5_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .Y(n_11) );
AOI222xp33_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_1), .B1(n_2), .B2(n_10), .C1(n_9), .C2(n_7), .Y(n_12) );
endmodule