module fake_jpeg_30700_n_456 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_456);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_456;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_8),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_74),
.Y(n_120)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_9),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_9),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_32),
.Y(n_127)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_38),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_88),
.Y(n_104)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_44),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_32),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_107),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_50),
.A2(n_44),
.B1(n_28),
.B2(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_35),
.B1(n_26),
.B2(n_29),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_44),
.B1(n_28),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_31),
.B1(n_22),
.B2(n_33),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_59),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_46),
.A2(n_30),
.B1(n_28),
.B2(n_32),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_113),
.A2(n_33),
.B1(n_25),
.B2(n_123),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_53),
.B(n_36),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_35),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_36),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_54),
.B(n_36),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_22),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_35),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_185),
.B1(n_137),
.B2(n_131),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_163),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_63),
.B1(n_48),
.B2(n_57),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_161),
.B1(n_173),
.B2(n_174),
.Y(n_195)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_106),
.A2(n_104),
.B(n_101),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_51),
.B1(n_68),
.B2(n_60),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_184),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_55),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_129),
.C(n_124),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_106),
.A2(n_77),
.B1(n_29),
.B2(n_26),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_80),
.B1(n_66),
.B2(n_73),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_179),
.B1(n_131),
.B2(n_94),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_172),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_78),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_110),
.A2(n_84),
.B1(n_49),
.B2(n_62),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_96),
.A2(n_65),
.B1(n_69),
.B2(n_87),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_22),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_98),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_100),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_25),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_13),
.B(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_108),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_100),
.B(n_25),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_121),
.A2(n_72),
.B1(n_33),
.B2(n_31),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_157),
.B1(n_165),
.B2(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_134),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_122),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_166),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_211),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_167),
.A2(n_126),
.B1(n_136),
.B2(n_132),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_158),
.B1(n_180),
.B2(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_155),
.Y(n_212)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_234),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_163),
.B(n_178),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_201),
.B(n_205),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_217),
.A2(n_218),
.B1(n_231),
.B2(n_232),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_181),
.B1(n_154),
.B2(n_161),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_181),
.C(n_177),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_160),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_185),
.B1(n_155),
.B2(n_167),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_223),
.B1(n_229),
.B2(n_212),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_155),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_179),
.B1(n_168),
.B2(n_170),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_170),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_172),
.B1(n_156),
.B2(n_117),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_176),
.C(n_156),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_200),
.C(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_173),
.B1(n_172),
.B2(n_121),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_99),
.B1(n_132),
.B2(n_128),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_204),
.B1(n_207),
.B2(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_244),
.C(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_262),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_197),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_203),
.B1(n_187),
.B2(n_208),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_233),
.B1(n_215),
.B2(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_255),
.B1(n_258),
.B2(n_261),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_251),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_240),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_207),
.C(n_191),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_254),
.A2(n_238),
.B(n_196),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_214),
.B1(n_201),
.B2(n_196),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_228),
.B(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_257),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_149),
.B1(n_139),
.B2(n_118),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_205),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_264),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_214),
.B1(n_149),
.B2(n_118),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_199),
.C(n_153),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_217),
.C(n_235),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_199),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_188),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_250),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_279),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_235),
.B1(n_216),
.B2(n_227),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_270),
.A2(n_271),
.B1(n_294),
.B2(n_287),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_281),
.C(n_288),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_276),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_235),
.C(n_218),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_283),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_286),
.B1(n_255),
.B2(n_258),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_226),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_291),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_287),
.B(n_294),
.Y(n_302)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_246),
.A2(n_237),
.B1(n_236),
.B2(n_234),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_226),
.B(n_190),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_188),
.C(n_182),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_248),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_193),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_242),
.A2(n_193),
.B(n_162),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_245),
.B(n_145),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_265),
.C(n_252),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_306),
.B1(n_308),
.B2(n_312),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_289),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_260),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_300),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_275),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_243),
.B1(n_250),
.B2(n_256),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_274),
.B(n_262),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_318),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_278),
.A2(n_250),
.B1(n_247),
.B2(n_261),
.Y(n_308)
);

OAI21x1_ASAP7_75t_SL g310 ( 
.A1(n_269),
.A2(n_250),
.B(n_264),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_277),
.B(n_270),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_269),
.A2(n_276),
.B1(n_285),
.B2(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_257),
.B1(n_251),
.B2(n_264),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_323),
.B1(n_324),
.B2(n_268),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_150),
.C(n_159),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_283),
.C(n_284),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_319),
.A2(n_295),
.B1(n_268),
.B2(n_291),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_152),
.B1(n_151),
.B2(n_147),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_277),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_128),
.B1(n_112),
.B2(n_94),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_273),
.A2(n_97),
.B1(n_112),
.B2(n_151),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_281),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_349),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_341),
.B1(n_342),
.B2(n_298),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_331),
.B(n_302),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_267),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_336),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_345),
.C(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_339),
.A2(n_344),
.B1(n_323),
.B2(n_322),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_309),
.B1(n_306),
.B2(n_296),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_97),
.B1(n_152),
.B2(n_126),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_343),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_319),
.A2(n_136),
.B1(n_189),
.B2(n_108),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_189),
.C(n_89),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_313),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_189),
.B(n_11),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_348),
.A2(n_10),
.B(n_13),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_108),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_340),
.A2(n_309),
.B1(n_308),
.B2(n_312),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_365),
.B1(n_330),
.B2(n_369),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_363),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_327),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_317),
.C(n_316),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_362),
.C(n_366),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_313),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_359),
.B(n_360),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_311),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_307),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_361),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_326),
.C(n_329),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_301),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_371),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_311),
.B1(n_298),
.B2(n_324),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_301),
.C(n_310),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_369),
.A2(n_346),
.B1(n_325),
.B2(n_342),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_344),
.B1(n_335),
.B2(n_325),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_380),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_364),
.B(n_331),
.CI(n_333),
.CON(n_375),
.SN(n_375)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_363),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_377),
.A2(n_352),
.B1(n_357),
.B2(n_11),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_353),
.A2(n_346),
.B1(n_341),
.B2(n_343),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_379),
.A2(n_382),
.B1(n_7),
.B2(n_17),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_333),
.B(n_347),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_381),
.A2(n_384),
.B(n_371),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_361),
.A2(n_348),
.B(n_11),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_383),
.A2(n_351),
.B(n_372),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_88),
.B(n_10),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_386),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_10),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_27),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_27),
.C(n_1),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_0),
.C(n_1),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_367),
.A2(n_7),
.B(n_17),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_368),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_402),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g410 ( 
.A1(n_397),
.A2(n_398),
.B(n_375),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_366),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_376),
.A2(n_372),
.B1(n_351),
.B2(n_370),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_400),
.A2(n_406),
.B1(n_383),
.B2(n_382),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_404),
.Y(n_413)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_354),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_405),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_391),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_403),
.B(n_389),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_409),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_378),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_417),
.B(n_387),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_394),
.B(n_385),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_393),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_397),
.A2(n_388),
.B(n_384),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_418),
.B(n_420),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_404),
.A2(n_401),
.B1(n_388),
.B2(n_398),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_390),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_422),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_416),
.B(n_399),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_11),
.B(n_17),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_399),
.B1(n_380),
.B2(n_407),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_427),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_413),
.B(n_419),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_27),
.C(n_1),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_432),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_27),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_5),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_27),
.Y(n_434)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_435),
.B(n_437),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_429),
.A2(n_5),
.B(n_14),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_429),
.A2(n_5),
.B(n_14),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_431),
.A2(n_5),
.B(n_13),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_441),
.B(n_12),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_4),
.B(n_12),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_428),
.C(n_423),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_443),
.B(n_444),
.C(n_446),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_445),
.A2(n_6),
.B(n_12),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_436),
.A2(n_430),
.B(n_6),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_6),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_447),
.A2(n_0),
.B(n_1),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_439),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_448),
.A2(n_450),
.B(n_451),
.Y(n_453)
);

AOI321xp33_ASAP7_75t_L g452 ( 
.A1(n_449),
.A2(n_12),
.A3(n_15),
.B1(n_3),
.B2(n_1),
.C(n_2),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_452),
.A2(n_453),
.B(n_15),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_2),
.B(n_3),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_2),
.Y(n_456)
);


endmodule