module real_aes_10281_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_102;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_85;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g123 ( .A(n_0), .B(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_1), .Y(n_530) );
INVx1_ASAP7_75t_L g610 ( .A(n_1), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_2), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_3), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g537 ( .A(n_4), .Y(n_537) );
INVx1_ASAP7_75t_L g533 ( .A(n_5), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_5), .A2(n_60), .B1(n_605), .B2(n_606), .Y(n_604) );
BUFx2_ASAP7_75t_L g527 ( .A(n_6), .Y(n_527) );
BUFx2_ASAP7_75t_L g581 ( .A(n_6), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_7), .B(n_133), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_9), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_10), .B(n_113), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_11), .B(n_119), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_12), .B(n_156), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_13), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_14), .B(n_119), .Y(n_199) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_16), .B(n_133), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_17), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_18), .B(n_156), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_19), .A2(n_76), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_19), .A2(n_76), .B1(n_617), .B2(n_618), .Y(n_616) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_20), .Y(n_677) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_21), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_22), .B(n_113), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_23), .B(n_181), .Y(n_206) );
INVx1_ASAP7_75t_L g579 ( .A(n_24), .Y(n_579) );
INVx1_ASAP7_75t_L g703 ( .A(n_24), .Y(n_703) );
NAND2xp33_ASAP7_75t_SL g170 ( .A(n_25), .B(n_90), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_26), .B(n_159), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_27), .B(n_115), .Y(n_183) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_28), .A2(n_48), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g475 ( .A(n_29), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_29), .A2(n_64), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_30), .A2(n_470), .B1(n_471), .B2(n_636), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_30), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_31), .A2(n_56), .B1(n_589), .B2(n_593), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_31), .A2(n_56), .B1(n_613), .B2(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_32), .B(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g83 ( .A(n_33), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_33), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_33), .B(n_663), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_34), .B(n_147), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_35), .B(n_147), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_36), .B(n_152), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_37), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_38), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_39), .Y(n_519) );
INVx1_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_40), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_41), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_42), .B(n_238), .Y(n_237) );
NAND2xp33_ASAP7_75t_L g168 ( .A(n_43), .B(n_90), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_44), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_45), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_46), .B(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g485 ( .A(n_47), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_49), .B(n_113), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_50), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g568 ( .A(n_51), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_51), .A2(n_67), .B1(n_600), .B2(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_52), .B(n_159), .Y(n_186) );
BUFx10_ASAP7_75t_L g697 ( .A(n_53), .Y(n_697) );
INVx2_ASAP7_75t_L g479 ( .A(n_54), .Y(n_479) );
INVx1_ASAP7_75t_L g503 ( .A(n_54), .Y(n_503) );
INVx1_ASAP7_75t_L g493 ( .A(n_55), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_55), .A2(n_74), .B1(n_626), .B2(n_628), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_55), .A2(n_522), .B(n_640), .C(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_57), .B(n_113), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_58), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_59), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g556 ( .A(n_60), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_60), .A2(n_653), .B(n_658), .C(n_659), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_61), .B(n_119), .Y(n_150) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_61), .Y(n_705) );
INVx2_ASAP7_75t_L g108 ( .A(n_62), .Y(n_108) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_63), .Y(n_682) );
INVx1_ASAP7_75t_L g486 ( .A(n_64), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_65), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_66), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g545 ( .A(n_67), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_68), .B(n_133), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_69), .Y(n_505) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_70), .Y(n_671) );
INVx2_ASAP7_75t_L g482 ( .A(n_71), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_72), .Y(n_197) );
BUFx3_ASAP7_75t_L g542 ( .A(n_73), .Y(n_542) );
INVx1_ASAP7_75t_L g572 ( .A(n_73), .Y(n_572) );
INVx1_ASAP7_75t_L g514 ( .A(n_74), .Y(n_514) );
BUFx3_ASAP7_75t_L g544 ( .A(n_75), .Y(n_544) );
INVx1_ASAP7_75t_L g550 ( .A(n_75), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_95), .B(n_468), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_SL g172 ( .A(n_82), .Y(n_172) );
INVx8_ASAP7_75t_L g185 ( .A(n_82), .Y(n_185) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
A2O1A1Ixp33_ASAP7_75t_L g109 ( .A1(n_83), .A2(n_110), .B(n_112), .C(n_117), .Y(n_109) );
OAI21x1_ASAP7_75t_SL g130 ( .A1(n_83), .A2(n_131), .B(n_138), .Y(n_130) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_83), .A2(n_149), .B(n_153), .Y(n_148) );
INVxp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g713 ( .A1(n_86), .A2(n_714), .B(n_715), .Y(n_713) );
NAND2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
INVx2_ASAP7_75t_L g115 ( .A(n_91), .Y(n_115) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_91), .Y(n_122) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
BUFx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_93), .A2(n_118), .B(n_120), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_93), .A2(n_139), .B(n_141), .Y(n_138) );
BUFx12f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx5_ASAP7_75t_L g111 ( .A(n_94), .Y(n_111) );
INVx5_ASAP7_75t_L g137 ( .A(n_94), .Y(n_137) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx3_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND3x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_345), .C(n_425), .Y(n_98) );
NOR2xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_283), .Y(n_99) );
NAND4xp25_ASAP7_75t_L g100 ( .A(n_101), .B(n_242), .C(n_264), .D(n_275), .Y(n_100) );
AOI322xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_161), .A3(n_187), .B1(n_214), .B2(n_217), .C1(n_223), .C2(n_227), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_126), .Y(n_102) );
INVx4_ASAP7_75t_L g287 ( .A(n_103), .Y(n_287) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g241 ( .A(n_104), .Y(n_241) );
AND2x2_ASAP7_75t_L g249 ( .A(n_104), .B(n_129), .Y(n_249) );
AND2x2_ASAP7_75t_L g280 ( .A(n_104), .B(n_272), .Y(n_280) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_109), .B(n_123), .Y(n_104) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_105), .A2(n_177), .B(n_186), .Y(n_176) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_105), .A2(n_191), .B(n_200), .Y(n_190) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_105), .A2(n_204), .B(n_212), .Y(n_203) );
BUFx5_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_106), .Y(n_213) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_110), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_110), .A2(n_209), .B(n_211), .Y(n_208) );
AOI21x1_ASAP7_75t_L g235 ( .A1(n_110), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g157 ( .A(n_111), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_111), .A2(n_166), .B(n_167), .C(n_168), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_111), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_111), .A2(n_233), .B(n_234), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
INVx2_ASAP7_75t_L g210 ( .A(n_115), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_116), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_116), .Y(n_680) );
INVx5_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
INVx1_ASAP7_75t_L g198 ( .A(n_121), .Y(n_198) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx2_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
INVx2_ASAP7_75t_L g194 ( .A(n_122), .Y(n_194) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_124), .A2(n_130), .B(n_142), .Y(n_129) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_124), .Y(n_230) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
INVx1_ASAP7_75t_L g266 ( .A(n_126), .Y(n_266) );
AND2x2_ASAP7_75t_L g408 ( .A(n_126), .B(n_280), .Y(n_408) );
AND2x2_ASAP7_75t_L g428 ( .A(n_126), .B(n_372), .Y(n_428) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_145), .Y(n_126) );
AND2x2_ASAP7_75t_L g240 ( .A(n_127), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g216 ( .A(n_128), .Y(n_216) );
AND2x2_ASAP7_75t_L g301 ( .A(n_128), .B(n_145), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_128), .B(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_128), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_128), .B(n_241), .Y(n_411) );
INVx1_ASAP7_75t_L g432 ( .A(n_128), .Y(n_432) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_128), .Y(n_451) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_135), .C(n_137), .Y(n_131) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g136 ( .A(n_134), .Y(n_136) );
INVx2_ASAP7_75t_L g238 ( .A(n_136), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_137), .A2(n_150), .B(n_151), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_137), .A2(n_183), .B(n_184), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_L g196 ( .A1(n_137), .A2(n_197), .B(n_198), .C(n_199), .Y(n_196) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_SL g147 ( .A(n_144), .Y(n_147) );
NOR2xp67_ASAP7_75t_L g215 ( .A(n_145), .B(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_145), .Y(n_279) );
INVx1_ASAP7_75t_L g289 ( .A(n_145), .Y(n_289) );
INVx1_ASAP7_75t_L g331 ( .A(n_145), .Y(n_331) );
AND2x2_ASAP7_75t_L g354 ( .A(n_145), .B(n_247), .Y(n_354) );
INVx1_ASAP7_75t_L g445 ( .A(n_145), .Y(n_445) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g344 ( .A(n_146), .B(n_247), .Y(n_344) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_158), .Y(n_146) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_147), .A2(n_164), .B(n_173), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_157), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_157), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_157), .A2(n_193), .B(n_195), .Y(n_192) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_161), .A2(n_389), .B1(n_402), .B2(n_405), .C(n_407), .Y(n_388) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g223 ( .A(n_162), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g446 ( .A(n_162), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_174), .Y(n_162) );
INVx2_ASAP7_75t_L g220 ( .A(n_163), .Y(n_220) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_163), .Y(n_385) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B(n_172), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B(n_196), .Y(n_191) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g258 ( .A(n_174), .Y(n_258) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g221 ( .A(n_175), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g263 ( .A(n_175), .Y(n_263) );
AND2x2_ASAP7_75t_L g295 ( .A(n_175), .B(n_262), .Y(n_295) );
INVx1_ASAP7_75t_L g384 ( .A(n_175), .Y(n_384) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI21x1_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_182), .B(n_185), .Y(n_177) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_185), .A2(n_205), .B(n_208), .Y(n_204) );
INVxp67_ASAP7_75t_L g282 ( .A(n_187), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_187), .A2(n_430), .B1(n_433), .B2(n_435), .Y(n_429) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_201), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_188), .B(n_297), .Y(n_339) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_188), .B(n_376), .Y(n_436) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_189), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
AND2x4_ASAP7_75t_L g224 ( .A(n_201), .B(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g338 ( .A(n_201), .Y(n_338) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_201), .Y(n_447) );
BUFx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g293 ( .A(n_202), .Y(n_293) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g400 ( .A(n_215), .B(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_216), .Y(n_350) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_221), .Y(n_217) );
OR2x2_ASAP7_75t_L g259 ( .A(n_218), .B(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g274 ( .A(n_218), .B(n_253), .Y(n_274) );
AND2x4_ASAP7_75t_L g322 ( .A(n_218), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g415 ( .A(n_218), .B(n_324), .Y(n_415) );
INVx1_ASAP7_75t_L g462 ( .A(n_218), .Y(n_462) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g257 ( .A(n_219), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_219), .B(n_254), .Y(n_269) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g298 ( .A(n_220), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_220), .B(n_255), .Y(n_335) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_220), .Y(n_360) );
AND2x2_ASAP7_75t_L g267 ( .A(n_221), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g307 ( .A(n_221), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g341 ( .A(n_221), .Y(n_341) );
AOI322xp5_ASAP7_75t_L g367 ( .A1(n_221), .A2(n_368), .A3(n_370), .B1(n_373), .B2(n_375), .C1(n_377), .C2(n_380), .Y(n_367) );
AND2x2_ASAP7_75t_L g404 ( .A(n_221), .B(n_292), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_221), .A2(n_355), .B1(n_423), .B2(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g226 ( .A(n_222), .Y(n_226) );
INVx2_ASAP7_75t_L g262 ( .A(n_222), .Y(n_262) );
INVx1_ASAP7_75t_L g310 ( .A(n_224), .Y(n_310) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_226), .B(n_293), .Y(n_324) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_240), .Y(n_227) );
AND2x2_ASAP7_75t_L g398 ( .A(n_228), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g455 ( .A(n_228), .B(n_301), .Y(n_455) );
INVxp67_ASAP7_75t_R g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_247) );
INVx2_ASAP7_75t_L g364 ( .A(n_240), .Y(n_364) );
AND2x2_ASAP7_75t_L g423 ( .A(n_240), .B(n_344), .Y(n_423) );
INVx1_ASAP7_75t_L g321 ( .A(n_241), .Y(n_321) );
AND2x2_ASAP7_75t_L g394 ( .A(n_241), .B(n_293), .Y(n_394) );
AND2x2_ASAP7_75t_L g401 ( .A(n_241), .B(n_272), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_250), .Y(n_242) );
OAI31xp33_ASAP7_75t_L g427 ( .A1(n_243), .A2(n_359), .A3(n_362), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
AND2x2_ASAP7_75t_L g362 ( .A(n_245), .B(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g372 ( .A(n_246), .Y(n_372) );
BUFx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g265 ( .A(n_248), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g314 ( .A(n_249), .B(n_293), .Y(n_314) );
AND2x2_ASAP7_75t_L g353 ( .A(n_249), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_249), .B(n_330), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_256), .Y(n_251) );
INVx1_ASAP7_75t_L g467 ( .A(n_252), .Y(n_467) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g357 ( .A(n_253), .Y(n_357) );
INVx2_ASAP7_75t_L g382 ( .A(n_254), .Y(n_382) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g376 ( .A(n_255), .B(n_298), .Y(n_376) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_256), .B(n_338), .Y(n_439) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g366 ( .A(n_257), .B(n_338), .Y(n_366) );
AND2x2_ASAP7_75t_L g317 ( .A(n_258), .B(n_298), .Y(n_317) );
INVx1_ASAP7_75t_L g412 ( .A(n_259), .Y(n_412) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g375 ( .A(n_261), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_261), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g458 ( .A(n_261), .B(n_292), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_261), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
BUFx2_ASAP7_75t_L g356 ( .A(n_263), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B1(n_270), .B2(n_273), .Y(n_264) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_270), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
AND2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
AND2x4_ASAP7_75t_L g361 ( .A(n_271), .B(n_301), .Y(n_361) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g288 ( .A(n_272), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_281), .C(n_282), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g349 ( .A(n_278), .B(n_350), .Y(n_349) );
NAND2x1_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_311), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .B1(n_299), .B2(n_302), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_287), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g329 ( .A(n_287), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_287), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g434 ( .A(n_287), .B(n_392), .Y(n_434) );
INVx2_ASAP7_75t_L g379 ( .A(n_288), .Y(n_379) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_292), .B(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g305 ( .A(n_295), .Y(n_305) );
AND2x2_ASAP7_75t_L g359 ( .A(n_295), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_297), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g374 ( .A(n_301), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .C(n_309), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_309), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_325), .B(n_327), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B(n_318), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_315), .A2(n_453), .B(n_456), .Y(n_452) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g466 ( .A(n_320), .B(n_344), .Y(n_466) );
AND2x2_ASAP7_75t_L g444 ( .A(n_321), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g457 ( .A(n_326), .B(n_410), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_332), .B(n_336), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_331), .B(n_399), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_334), .A2(n_443), .B1(n_446), .B2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_340), .B(n_342), .Y(n_336) );
NOR2x1_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_338), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g460 ( .A(n_338), .Y(n_460) );
INVx1_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
INVx1_ASAP7_75t_L g441 ( .A(n_340), .Y(n_441) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_344), .B(n_410), .Y(n_421) );
AND2x2_ASAP7_75t_L g424 ( .A(n_344), .B(n_410), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_344), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g464 ( .A(n_344), .B(n_451), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_388), .C(n_413), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_358), .C(n_367), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_351), .B(n_355), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g378 ( .A(n_350), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
INVx2_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_354), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_362), .B2(n_365), .Y(n_358) );
INVx2_ASAP7_75t_L g440 ( .A(n_361), .Y(n_440) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x6_ASAP7_75t_L g405 ( .A(n_364), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_381), .B(n_386), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI221xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_393), .B1(n_395), .B2(n_398), .C(n_400), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g454 ( .A(n_393), .B(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_395), .A2(n_408), .B1(n_409), .B2(n_412), .Y(n_407) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g443 ( .A(n_398), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_416), .C(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_421), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_418), .A2(n_438), .B1(n_440), .B2(n_441), .C(n_442), .Y(n_437) );
OR2x6_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_437), .C(n_452), .D(n_461), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_465), .C(n_467), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_661), .B2(n_666), .C(n_709), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_471), .A2(n_705), .B1(n_710), .B2(n_712), .Y(n_709) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI221x1_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_525), .B1(n_531), .B2(n_576), .C(n_582), .Y(n_472) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_492), .C(n_513), .D(n_522), .Y(n_473) );
INVx1_ASAP7_75t_L g649 ( .A(n_474), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_486), .B2(n_487), .Y(n_474) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .Y(n_476) );
AND2x4_ASAP7_75t_L g487 ( .A(n_477), .B(n_488), .Y(n_487) );
OR2x6_ASAP7_75t_L g521 ( .A(n_477), .B(n_517), .Y(n_521) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g512 ( .A(n_479), .Y(n_512) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_480), .Y(n_586) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_480), .Y(n_600) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g490 ( .A(n_482), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_482), .Y(n_497) );
INVx1_ASAP7_75t_L g509 ( .A(n_482), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_482), .B(n_485), .Y(n_518) );
AND2x2_ASAP7_75t_L g592 ( .A(n_482), .B(n_485), .Y(n_592) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g491 ( .A(n_485), .Y(n_491) );
INVx1_ASAP7_75t_L g504 ( .A(n_485), .Y(n_504) );
INVx1_ASAP7_75t_L g644 ( .A(n_485), .Y(n_644) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
INVx3_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
AND2x4_ASAP7_75t_L g496 ( .A(n_491), .B(n_497), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_498), .B2(n_499), .C1(n_505), .C2(n_506), .Y(n_492) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g523 ( .A(n_496), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g594 ( .A(n_496), .Y(n_594) );
BUFx3_ASAP7_75t_L g606 ( .A(n_496), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g551 ( .A1(n_498), .A2(n_505), .B1(n_552), .B2(n_556), .C1(n_557), .C2(n_564), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_498), .A2(n_505), .B1(n_646), .B2(n_648), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_498), .A2(n_505), .B1(n_558), .B2(n_564), .Y(n_659) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g647 ( .A(n_501), .Y(n_647) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
OR2x6_ASAP7_75t_L g516 ( .A(n_502), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_529), .Y(n_597) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_510), .Y(n_506) );
AND2x4_ASAP7_75t_L g648 ( .A(n_507), .B(n_510), .Y(n_648) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g643 ( .A(n_509), .B(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g524 ( .A(n_511), .Y(n_524) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_512), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g638 ( .A(n_513), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_519), .B2(n_520), .Y(n_513) );
INVx8_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_519), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx11_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
OAI31xp33_ASAP7_75t_L g637 ( .A1(n_525), .A2(n_638), .A3(n_639), .B(n_649), .Y(n_637) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x4_ASAP7_75t_L g633 ( .A(n_527), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_532), .B(n_551), .C(n_566), .D(n_573), .Y(n_531) );
INVxp67_ASAP7_75t_L g651 ( .A(n_532), .Y(n_651) );
AOI22xp5_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_534), .B1(n_545), .B2(n_546), .Y(n_532) );
AND2x4_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
AND2x6_ASAP7_75t_L g569 ( .A(n_535), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_537), .Y(n_560) );
AND2x2_ASAP7_75t_L g623 ( .A(n_537), .B(n_579), .Y(n_623) );
INVx2_ASAP7_75t_L g635 ( .A(n_537), .Y(n_635) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_539), .Y(n_627) );
INVx6_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g567 ( .A(n_540), .B(n_559), .Y(n_567) );
BUFx2_ASAP7_75t_L g613 ( .A(n_540), .Y(n_613) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g565 ( .A(n_541), .Y(n_565) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g549 ( .A(n_542), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g555 ( .A(n_542), .B(n_544), .Y(n_555) );
INVx1_ASAP7_75t_L g563 ( .A(n_543), .Y(n_563) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g571 ( .A(n_544), .B(n_572), .Y(n_571) );
AND2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g575 ( .A(n_547), .Y(n_575) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x6_ASAP7_75t_L g564 ( .A(n_548), .B(n_565), .Y(n_564) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_549), .Y(n_617) );
BUFx3_ASAP7_75t_L g631 ( .A(n_549), .Y(n_631) );
INVx1_ASAP7_75t_L g657 ( .A(n_550), .Y(n_657) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g574 ( .A(n_554), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g629 ( .A(n_554), .Y(n_629) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_555), .Y(n_615) );
BUFx4f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g695 ( .A(n_563), .Y(n_695) );
INVxp67_ASAP7_75t_L g660 ( .A(n_566), .Y(n_660) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_570), .Y(n_632) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g619 ( .A(n_571), .Y(n_619) );
INVx1_ASAP7_75t_L g656 ( .A(n_572), .Y(n_656) );
INVx5_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx8_ASAP7_75t_R g658 ( .A(n_574), .Y(n_658) );
OAI31xp33_ASAP7_75t_L g650 ( .A1(n_576), .A2(n_651), .A3(n_652), .B(n_660), .Y(n_650) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g634 ( .A(n_579), .B(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g596 ( .A(n_581), .Y(n_596) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_583), .B(n_637), .C(n_650), .Y(n_636) );
AND4x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_598), .C(n_611), .D(n_624), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .C(n_595), .Y(n_584) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g605 ( .A(n_591), .Y(n_605) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g607 ( .A(n_596), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g621 ( .A(n_596), .B(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_604), .C(n_607), .Y(n_598) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .C(n_620), .Y(n_611) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g691 ( .A(n_623), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_630), .C(n_633), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g701 ( .A(n_635), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_663), .B(n_665), .Y(n_687) );
INVx1_ASAP7_75t_SL g714 ( .A(n_663), .Y(n_714) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_683), .B1(n_705), .B2(n_706), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_667), .A2(n_705), .B1(n_708), .B2(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_678), .B2(n_679), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx8_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx8_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
CKINVDCx20_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_686), .Y(n_711) );
OR2x6_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OR2x4_ASAP7_75t_L g708 ( .A(n_687), .B(n_689), .Y(n_708) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI31xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .A3(n_696), .B(n_698), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g704 ( .A(n_695), .Y(n_704) );
INVx6_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx8_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
BUFx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
endmodule