module real_jpeg_6680_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_0),
.A2(n_150),
.B1(n_153),
.B2(n_156),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_0),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_173),
.C(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_0),
.B(n_78),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_0),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_0),
.B(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_0),
.B(n_266),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_1),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_1),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_2),
.A2(n_57),
.B1(n_92),
.B2(n_132),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_2),
.A2(n_92),
.B1(n_386),
.B2(n_388),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_2),
.A2(n_92),
.B1(n_251),
.B2(n_419),
.Y(n_418)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_3),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_3),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_3),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_3),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_4),
.A2(n_122),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_4),
.A2(n_181),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_4),
.A2(n_181),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_4),
.A2(n_60),
.B1(n_181),
.B2(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_5),
.Y(n_335)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_7),
.A2(n_61),
.B1(n_226),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_7),
.A2(n_61),
.B1(n_166),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_7),
.A2(n_61),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_8),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_12),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_162),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_162),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_12),
.A2(n_162),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_159),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_14),
.A2(n_208),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_14),
.A2(n_45),
.B1(n_208),
.B2(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_14),
.A2(n_36),
.B1(n_52),
.B2(n_208),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_15),
.A2(n_53),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_15),
.A2(n_53),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_15),
.A2(n_53),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_16),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_16),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_16),
.A2(n_98),
.B1(n_104),
.B2(n_126),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_16),
.A2(n_36),
.B1(n_98),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_16),
.A2(n_98),
.B1(n_182),
.B2(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_17),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_17),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_17),
.A2(n_279),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_17),
.A2(n_279),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_L g458 ( 
.A1(n_17),
.A2(n_279),
.B1(n_332),
.B2(n_459),
.Y(n_458)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_534),
.B(n_537),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_139),
.B(n_533),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_136),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_27),
.B(n_136),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_130),
.C(n_133),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_28),
.A2(n_29),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_62),
.C(n_99),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_30),
.B(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_31),
.A2(n_54),
.B1(n_56),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_31),
.A2(n_54),
.B1(n_131),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_31),
.A2(n_359),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_31),
.A2(n_54),
.B1(n_413),
.B2(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_31),
.A2(n_50),
.B1(n_54),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_32),
.A2(n_339),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_32),
.B(n_360),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_32),
.A2(n_55),
.B(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_40),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_36),
.Y(n_361)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_44),
.Y(n_411)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_49),
.Y(n_337)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_51),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_54),
.B(n_156),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_54),
.A2(n_433),
.B(n_460),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_55),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_55),
.B(n_458),
.Y(n_457)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_62),
.A2(n_99),
.B1(n_100),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_62),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_62)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_63),
.A2(n_93),
.B1(n_303),
.B2(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_63),
.A2(n_93),
.B1(n_402),
.B2(n_407),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_63),
.A2(n_88),
.B1(n_93),
.B2(n_510),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_69),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_72),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_72),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_72),
.Y(n_331)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_72),
.Y(n_338)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_77),
.Y(n_305)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_77),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_78),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_78),
.A2(n_134),
.B1(n_307),
.B2(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_78),
.A2(n_134),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_81),
.Y(n_374)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_81),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_82),
.Y(n_256)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_83),
.Y(n_399)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_86),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_90),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_91),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_93),
.B(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_93),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_99),
.A2(n_100),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_99),
.B(n_505),
.C(n_508),
.Y(n_516)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_114),
.B(n_125),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_149),
.B(n_157),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_101),
.A2(n_114),
.B1(n_206),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_101),
.A2(n_157),
.B(n_250),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_101),
.A2(n_114),
.B1(n_372),
.B2(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_102),
.B(n_158),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_102),
.A2(n_167),
.B1(n_393),
.B2(n_396),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_102),
.A2(n_167),
.B1(n_396),
.B2(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_102),
.A2(n_167),
.B1(n_418),
.B2(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_106),
.Y(n_253)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_106),
.Y(n_376)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_114),
.A2(n_206),
.B(n_209),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_114),
.A2(n_209),
.B(n_372),
.Y(n_371)
);

AOI22x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_120),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_122),
.B(n_216),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_123),
.Y(n_316)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_123),
.Y(n_387)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_125),
.Y(n_449)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_130),
.B(n_133),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_134),
.A2(n_259),
.B(n_267),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_134),
.B(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_134),
.A2(n_267),
.B(n_473),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_136),
.B(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_136),
.B(n_535),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_137),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_527),
.B(n_532),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_499),
.B(n_524),
.Y(n_140)
);

OAI311xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_379),
.A3(n_475),
.B1(n_493),
.C1(n_498),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_322),
.B(n_378),
.Y(n_142)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_294),
.B(n_321),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_244),
.B(n_293),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_212),
.B(n_243),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_178),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_147),
.B(n_178),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_168),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_148),
.A2(n_168),
.B1(n_169),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_156),
.A2(n_187),
.B(n_190),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_156),
.A2(n_260),
.B(n_264),
.Y(n_259)
);

HAxp5_ASAP7_75t_SL g339 ( 
.A(n_156),
.B(n_340),
.CON(n_339),
.SN(n_339)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_167),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_SL g420 ( 
.A(n_171),
.Y(n_420)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_203),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_204),
.C(n_211),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_187),
.B(n_190),
.Y(n_179)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_187),
.A2(n_345),
.B1(n_346),
.B2(n_349),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_187),
.A2(n_282),
.B1(n_385),
.B2(n_389),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_187),
.A2(n_230),
.B(n_389),
.Y(n_421)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_188),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_188),
.A2(n_277),
.B1(n_311),
.B2(n_317),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_188),
.A2(n_350),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_199),
.Y(n_312)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_201),
.Y(n_391)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_210),
.B2(n_211),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_234),
.B(n_242),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B(n_233),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_232),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_230),
.B(n_231),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_276),
.B(n_282),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_240),
.Y(n_242)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_246),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_274),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_257),
.B2(n_258),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_257),
.C(n_274),
.Y(n_295)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_252),
.B(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_253),
.Y(n_395)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_263),
.Y(n_408)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_263),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_285),
.A3(n_286),
.B1(n_289),
.B2(n_291),
.Y(n_284)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_281),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_295),
.B(n_296),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_320),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_300),
.C(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_309),
.C(n_310),
.Y(n_352)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_323),
.B(n_324),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_355),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_325)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_343),
.B2(n_344),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_328),
.B(n_343),
.Y(n_471)
);

OAI32xp33_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_332),
.A3(n_334),
.B1(n_336),
.B2(n_339),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_352),
.B(n_354),
.C(n_355),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_364),
.B2(n_377),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_356),
.B(n_365),
.C(n_371),
.Y(n_484)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_371),
.Y(n_364)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_461),
.Y(n_379)
);

A2O1A1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_380),
.A2(n_461),
.B(n_494),
.C(n_497),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_436),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_381),
.B(n_436),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_415),
.C(n_423),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_382),
.B(n_415),
.CI(n_423),
.CON(n_474),
.SN(n_474)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_400),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_401),
.C(n_412),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_392),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_392),
.Y(n_467)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_412),
.Y(n_400)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_421),
.B2(n_422),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_421),
.Y(n_453)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_421),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_422),
.B1(n_455),
.B2(n_456),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_421),
.A2(n_453),
.B(n_456),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_431),
.C(n_434),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_427),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_427),
.Y(n_483)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_434),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_440),
.C(n_451),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_451),
.B2(n_452),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_447),
.B(n_450),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_448),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_450),
.B(n_502),
.CI(n_503),
.CON(n_501),
.SN(n_501)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_450),
.B(n_502),
.C(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_474),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.C(n_468),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.C(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_472),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_474),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_485),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.C(n_484),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_491),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_490),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_513),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_512),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_512),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_501),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_507),
.B2(n_511),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_505),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_515),
.C(n_519),
.Y(n_531)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_523),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_523),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_531),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_530),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_538),
.Y(n_537)
);


endmodule