module fake_jpeg_14236_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_56),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_21),
.B(n_46),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_0),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_70),
.B1(n_52),
.B2(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_25),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_73),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_61),
.B(n_68),
.C(n_59),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_112),
.B(n_8),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_117),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_67),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_110),
.C(n_114),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_60),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_109),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_69),
.B(n_65),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_22),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_87),
.B1(n_97),
.B2(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_52),
.C(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_13),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_56),
.B1(n_55),
.B2(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_55),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_123),
.B1(n_131),
.B2(n_20),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_128),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_7),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_107),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_27),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_136),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_16),
.CI(n_19),
.CON(n_136),
.SN(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_122),
.B1(n_132),
.B2(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_144),
.B1(n_147),
.B2(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_26),
.B(n_29),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_125),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_31),
.B(n_32),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_39),
.B1(n_42),
.B2(n_48),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_125),
.C(n_121),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_141),
.C(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_154),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_146),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_155),
.A3(n_145),
.B1(n_163),
.B2(n_147),
.C1(n_152),
.C2(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_142),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_160),
.Y(n_168)
);


endmodule