module real_jpeg_14087_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_248, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_248;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_58),
.B1(n_61),
.B2(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_108),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_7),
.B(n_61),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_7),
.A2(n_63),
.B(n_165),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_98),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_44),
.B(n_48),
.C(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_7),
.B(n_104),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_32),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_84),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_61),
.B(n_156),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_52),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_10),
.A2(n_52),
.B1(n_58),
.B2(n_61),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_58),
.B1(n_61),
.B2(n_67),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_67),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_58),
.B1(n_61),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_12),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_77),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_77),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_58),
.B1(n_61),
.B2(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_69),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_15),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_16),
.A2(n_42),
.B1(n_58),
.B2(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_146)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_21),
.B(n_112),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_79),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_22),
.A2(n_23),
.B1(n_79),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_55),
.C(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_26),
.B(n_39),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_27),
.A2(n_31),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_28),
.A2(n_32),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_28),
.A2(n_32),
.B(n_87),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_28),
.A2(n_32),
.B1(n_94),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_28),
.A2(n_32),
.B1(n_146),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_28),
.A2(n_32),
.B1(n_159),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_28),
.A2(n_32),
.B1(n_98),
.B2(n_205),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_28),
.A2(n_32),
.B1(n_198),
.B2(n_205),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_36),
.A2(n_49),
.B(n_98),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_41),
.A2(n_46),
.B1(n_84),
.B2(n_150),
.Y(n_168)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_44),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_43),
.A2(n_61),
.A3(n_73),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_44),
.B(n_74),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_45),
.A2(n_50),
.B1(n_149),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_46),
.A2(n_83),
.B1(n_84),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_46),
.A2(n_84),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_46),
.A2(n_84),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_46),
.A2(n_84),
.B1(n_184),
.B2(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_70),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_56),
.A2(n_57),
.B1(n_68),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_56),
.A2(n_57),
.B1(n_107),
.B2(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_61),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_60),
.A3(n_63),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_61),
.Y(n_96)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_71),
.A2(n_75),
.B1(n_101),
.B2(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_71),
.A2(n_75),
.B1(n_140),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_79),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_89),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_90),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_105),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_91),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_97),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_99),
.B(n_105),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_104),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_118),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI221xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_232),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_176),
.B(n_231),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_160),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_136),
.B(n_160),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.C(n_151),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_137),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_144),
.C(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_147),
.A2(n_151),
.B1(n_152),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_153),
.A2(n_154),
.B1(n_158),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_175),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_172),
.C(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_225),
.B(n_230),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_224),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_194),
.B(n_213),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_202),
.B(n_212),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_200),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);


endmodule