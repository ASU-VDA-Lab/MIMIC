module fake_jpeg_28645_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_28),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_12),
.B1(n_18),
.B2(n_13),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_49),
.B1(n_36),
.B2(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_14),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_31),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_70),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_22),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_17),
.B1(n_44),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_30),
.B1(n_50),
.B2(n_52),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_74),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_54),
.B(n_46),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_80),
.B(n_70),
.C(n_69),
.D(n_54),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_17),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_86),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_58),
.B(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_80),
.C(n_77),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_72),
.A3(n_75),
.B1(n_54),
.B2(n_46),
.C1(n_59),
.C2(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_77),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_90),
.C(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_83),
.B1(n_72),
.B2(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_89),
.B1(n_67),
.B2(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_62),
.B1(n_63),
.B2(n_2),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_94),
.B(n_81),
.C(n_10),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_2),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_98),
.C(n_10),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_9),
.C(n_46),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_27),
.Y(n_102)
);


endmodule