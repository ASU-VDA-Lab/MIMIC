module fake_netlist_5_424_n_15103 (n_924, n_1263, n_3304, n_977, n_1378, n_2253, n_2417, n_611, n_2756, n_1126, n_1423, n_1729, n_2739, n_1166, n_2380, n_1751, n_469, n_1508, n_82, n_2771, n_785, n_3241, n_549, n_2617, n_2200, n_3261, n_3006, n_532, n_1161, n_3027, n_1859, n_2746, n_1677, n_1150, n_2327, n_3179, n_3127, n_226, n_1780, n_3256, n_1488, n_667, n_2899, n_2955, n_790, n_3619, n_1055, n_3541, n_3622, n_2386, n_3596, n_1501, n_111, n_2395, n_880, n_3086, n_3297, n_544, n_1007, n_2369, n_155, n_2927, n_552, n_1528, n_2683, n_1370, n_1292, n_2347, n_2520, n_2821, n_1198, n_1360, n_2388, n_1099, n_2568, n_956, n_564, n_423, n_1738, n_2021, n_21, n_2134, n_3064, n_2391, n_105, n_3088, n_1021, n_1960, n_2843, n_2185, n_4, n_3270, n_551, n_2143, n_2853, n_3615, n_2059, n_1323, n_1466, n_688, n_1695, n_2487, n_1353, n_800, n_3595, n_3246, n_3202, n_1347, n_2495, n_2880, n_1535, n_1789, n_1666, n_3350, n_2389, n_671, n_819, n_1451, n_1022, n_2302, n_915, n_1545, n_2374, n_864, n_173, n_859, n_951, n_3341, n_1947, n_1264, n_3587, n_2114, n_3445, n_447, n_247, n_2001, n_1494, n_3407, n_3571, n_3599, n_292, n_625, n_854, n_1462, n_1799, n_2069, n_2396, n_3621, n_1580, n_674, n_417, n_1939, n_2486, n_3434, n_1806, n_516, n_933, n_2244, n_2257, n_1152, n_3501, n_3448, n_497, n_1869, n_1607, n_1563, n_606, n_3019, n_275, n_3039, n_2011, n_2096, n_26, n_877, n_2105, n_2538, n_2024, n_2, n_2530, n_1696, n_2483, n_3163, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_307, n_1860, n_2543, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_2031, n_2076, n_2482, n_3036, n_2677, n_1230, n_668, n_375, n_301, n_1896, n_2165, n_2147, n_929, n_3010, n_3180, n_3379, n_3532, n_2770, n_1124, n_1818, n_2127, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_2584, n_1257, n_2639, n_171, n_1182, n_3188, n_3325, n_3107, n_3531, n_3403, n_579, n_1698, n_1261, n_2329, n_938, n_1098, n_2963, n_3624, n_2142, n_3186, n_3461, n_3082, n_320, n_1154, n_2189, n_3332, n_1242, n_3283, n_1135, n_3048, n_3258, n_24, n_406, n_519, n_2323, n_2203, n_2597, n_1016, n_1243, n_546, n_2959, n_101, n_3340, n_2047, n_1280, n_3277, n_1845, n_281, n_240, n_2052, n_2193, n_2978, n_2058, n_2458, n_2478, n_291, n_231, n_257, n_2761, n_731, n_371, n_1483, n_2888, n_1314, n_1512, n_3157, n_709, n_1490, n_317, n_1236, n_1633, n_2537, n_2983, n_569, n_2669, n_2144, n_1778, n_3214, n_227, n_2306, n_920, n_2515, n_3022, n_1289, n_1517, n_2091, n_2466, n_2635, n_2652, n_94, n_335, n_3631, n_2715, n_3087, n_2085, n_3489, n_1669, n_2566, n_370, n_976, n_1949, n_343, n_1449, n_308, n_1946, n_2936, n_1566, n_2032, n_297, n_2587, n_156, n_2149, n_1078, n_2782, n_1670, n_2672, n_775, n_219, n_3060, n_157, n_2651, n_3490, n_600, n_1484, n_2071, n_2561, n_1374, n_1328, n_2643, n_223, n_2141, n_1948, n_3013, n_3183, n_1984, n_3437, n_2099, n_2408, n_3446, n_3353, n_264, n_1877, n_1831, n_1598, n_3049, n_1723, n_955, n_1850, n_163, n_3028, n_339, n_1146, n_882, n_183, n_243, n_2384, n_1036, n_1097, n_1749, n_347, n_3156, n_59, n_550, n_696, n_3101, n_897, n_215, n_350, n_196, n_798, n_3376, n_646, n_1428, n_2663, n_436, n_1394, n_2659, n_1414, n_1216, n_290, n_580, n_2693, n_1040, n_2202, n_2648, n_1872, n_3389, n_1852, n_2159, n_578, n_2976, n_926, n_2180, n_2249, n_344, n_2353, n_1218, n_1931, n_2439, n_2632, n_2276, n_3089, n_422, n_475, n_777, n_1070, n_1547, n_2089, n_3420, n_1030, n_72, n_2470, n_1755, n_3222, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1801, n_1391, n_958, n_1034, n_670, n_1513, n_2908, n_2970, n_3361, n_1600, n_48, n_521, n_663, n_845, n_2235, n_1862, n_673, n_837, n_1239, n_2915, n_528, n_2300, n_2791, n_1796, n_2551, n_3291, n_680, n_1473, n_1587, n_2682, n_395, n_164, n_553, n_901, n_2432, n_813, n_1521, n_1284, n_1590, n_3440, n_3405, n_214, n_2174, n_2714, n_1748, n_3563, n_2934, n_1672, n_2506, n_675, n_2699, n_888, n_1880, n_2769, n_3542, n_2337, n_3436, n_1167, n_1626, n_3550, n_637, n_2615, n_1384, n_1556, n_184, n_446, n_1863, n_1064, n_144, n_858, n_2079, n_2238, n_114, n_96, n_923, n_2118, n_691, n_1151, n_2985, n_2944, n_881, n_1405, n_2407, n_1706, n_468, n_3418, n_213, n_129, n_342, n_2932, n_2753, n_464, n_2980, n_363, n_1582, n_197, n_1069, n_3306, n_1784, n_2859, n_2842, n_1075, n_3262, n_3136, n_1836, n_2868, n_3395, n_1450, n_3141, n_1322, n_2101, n_1471, n_1986, n_2863, n_2072, n_3164, n_2738, n_1750, n_3570, n_1459, n_460, n_889, n_2358, n_973, n_2968, n_1700, n_2833, n_477, n_3191, n_571, n_1585, n_461, n_2684, n_2712, n_3593, n_3193, n_1971, n_1599, n_3252, n_2275, n_2855, n_3507, n_3273, n_2713, n_3544, n_2644, n_2700, n_1211, n_1197, n_3367, n_2951, n_1523, n_2730, n_1950, n_3008, n_907, n_1447, n_2251, n_3096, n_1377, n_2370, n_190, n_3496, n_989, n_2544, n_1039, n_2214, n_3339, n_34, n_2055, n_3427, n_228, n_283, n_3025, n_3349, n_1403, n_2248, n_2356, n_488, n_736, n_892, n_3320, n_3007, n_2688, n_1000, n_1202, n_2750, n_2620, n_1278, n_2622, n_2062, n_2668, n_1002, n_1463, n_1581, n_2100, n_49, n_3071, n_310, n_3310, n_54, n_593, n_3487, n_2258, n_12, n_748, n_586, n_1058, n_1667, n_3359, n_838, n_2784, n_2919, n_332, n_3092, n_1053, n_3470, n_1224, n_2865, n_349, n_2557, n_1926, n_2706, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_2150, n_3146, n_2241, n_2757, n_2152, n_3598, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_2590, n_2776, n_2140, n_2385, n_3580, n_1819, n_2330, n_2139, n_2942, n_476, n_2987, n_1527, n_2042, n_534, n_3106, n_1882, n_884, n_3328, n_345, n_944, n_1754, n_3611, n_1623, n_2862, n_2175, n_2921, n_2720, n_2324, n_1854, n_91, n_2606, n_2674, n_3187, n_1565, n_3508, n_2828, n_3371, n_1809, n_1856, n_182, n_143, n_647, n_3433, n_237, n_407, n_1072, n_2218, n_2267, n_832, n_857, n_2305, n_3392, n_3430, n_2636, n_2450, n_3208, n_207, n_561, n_1319, n_2379, n_3331, n_3447, n_2616, n_2911, n_3305, n_2154, n_1825, n_1951, n_1883, n_1906, n_2759, n_1712, n_1387, n_3528, n_2262, n_2462, n_2514, n_1532, n_2322, n_2271, n_2625, n_18, n_3257, n_3625, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_2798, n_2331, n_2945, n_2293, n_686, n_2837, n_847, n_1393, n_2319, n_596, n_1775, n_2979, n_3296, n_2028, n_1368, n_3481, n_2762, n_558, n_2808, n_702, n_1276, n_3009, n_2548, n_822, n_1412, n_2676, n_1709, n_2679, n_2108, n_728, n_266, n_1162, n_272, n_1538, n_2930, n_1838, n_1199, n_1847, n_1779, n_2767, n_2777, n_2603, n_3514, n_3116, n_352, n_1884, n_2434, n_2660, n_53, n_3602, n_1038, n_2967, n_520, n_1369, n_409, n_2611, n_1841, n_1660, n_887, n_1905, n_2553, n_154, n_3207, n_2581, n_71, n_2195, n_2529, n_3224, n_300, n_2698, n_809, n_870, n_931, n_599, n_1711, n_1662, n_1891, n_1481, n_2626, n_3441, n_3042, n_1942, n_434, n_1978, n_1544, n_2510, n_3047, n_3526, n_868, n_2454, n_639, n_2804, n_914, n_2120, n_411, n_414, n_2546, n_1629, n_1293, n_2801, n_3120, n_965, n_1876, n_1743, n_3491, n_935, n_121, n_1175, n_817, n_2763, n_360, n_36, n_1479, n_1810, n_2350, n_2813, n_64, n_2825, n_1888, n_2009, n_759, n_2222, n_1892, n_3510, n_28, n_806, n_2990, n_1997, n_2667, n_1766, n_3218, n_1477, n_3142, n_324, n_1635, n_1963, n_2226, n_1571, n_2891, n_3119, n_187, n_1189, n_2690, n_103, n_97, n_3370, n_11, n_2215, n_3479, n_7, n_1259, n_1690, n_706, n_746, n_1649, n_3150, n_747, n_2064, n_52, n_784, n_110, n_2449, n_1733, n_1244, n_3500, n_2413, n_431, n_1194, n_1925, n_2297, n_1815, n_3279, n_2621, n_615, n_851, n_1759, n_843, n_1788, n_2177, n_2491, n_523, n_913, n_1537, n_705, n_865, n_61, n_2227, n_678, n_2671, n_697, n_127, n_1222, n_75, n_1679, n_2190, n_3346, n_776, n_1798, n_2022, n_1790, n_2518, n_2876, n_1415, n_367, n_2629, n_2592, n_3416, n_452, n_525, n_3484, n_3620, n_1260, n_1746, n_1647, n_2181, n_2479, n_2838, n_1829, n_1464, n_3133, n_3513, n_649, n_547, n_2563, n_43, n_1444, n_1191, n_2387, n_2992, n_1674, n_1833, n_116, n_3138, n_1830, n_2517, n_2073, n_1710, n_284, n_1128, n_2928, n_3128, n_139, n_1734, n_3038, n_744, n_590, n_629, n_2631, n_1308, n_2871, n_2178, n_3068, n_1767, n_3144, n_2943, n_2913, n_2336, n_3143, n_3168, n_254, n_1680, n_1233, n_3469, n_2607, n_23, n_1615, n_1529, n_2005, n_526, n_1916, n_3317, n_293, n_372, n_677, n_244, n_47, n_1333, n_2469, n_1121, n_2723, n_3355, n_314, n_368, n_433, n_604, n_2007, n_8, n_3220, n_949, n_2539, n_3263, n_100, n_2582, n_1443, n_1008, n_946, n_1539, n_2736, n_1001, n_1503, n_2054, n_498, n_1468, n_1559, n_1765, n_3455, n_1866, n_689, n_3158, n_738, n_1624, n_3000, n_640, n_3452, n_1510, n_252, n_624, n_1380, n_1744, n_2623, n_1617, n_295, n_133, n_1010, n_1994, n_1231, n_739, n_1279, n_1406, n_3108, n_3113, n_3111, n_2718, n_1195, n_1837, n_1839, n_610, n_2577, n_1760, n_2875, n_936, n_568, n_1500, n_2960, n_39, n_1090, n_2796, n_757, n_3280, n_2342, n_633, n_2856, n_439, n_3471, n_106, n_1832, n_259, n_448, n_1851, n_758, n_999, n_3205, n_2046, n_2848, n_2741, n_2937, n_3003, n_3610, n_1933, n_2290, n_93, n_1656, n_3564, n_3288, n_1158, n_3095, n_2045, n_3369, n_1509, n_1874, n_2040, n_563, n_2060, n_3199, n_2613, n_1987, n_2805, n_1145, n_878, n_524, n_3457, n_204, n_394, n_1678, n_1049, n_1153, n_2145, n_741, n_1639, n_1306, n_1068, n_3030, n_3558, n_1871, n_2580, n_3630, n_2545, n_2787, n_2914, n_1964, n_2869, n_122, n_331, n_10, n_906, n_1163, n_3271, n_2039, n_1207, n_919, n_908, n_2412, n_2406, n_3623, n_90, n_2846, n_724, n_1781, n_2084, n_2925, n_2035, n_658, n_2061, n_3555, n_3579, n_3075, n_3173, n_2378, n_2509, n_1740, n_3236, n_2398, n_1362, n_2857, n_1586, n_456, n_959, n_2459, n_3031, n_535, n_152, n_3396, n_940, n_1445, n_9, n_3516, n_1492, n_2155, n_2516, n_1923, n_1773, n_592, n_3243, n_1169, n_45, n_1596, n_1692, n_2666, n_2982, n_3385, n_1017, n_2481, n_2947, n_3545, n_2171, n_123, n_978, n_2768, n_2116, n_2314, n_1434, n_1054, n_2507, n_1474, n_1665, n_1269, n_2420, n_2900, n_1095, n_3343, n_3515, n_1828, n_1614, n_2886, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_2093, n_2038, n_2320, n_2339, n_2473, n_3287, n_2137, n_3378, n_603, n_1431, n_2583, n_484, n_1593, n_1033, n_442, n_3426, n_3454, n_2299, n_131, n_2540, n_2873, n_636, n_660, n_3410, n_2087, n_1640, n_2162, n_1732, n_1009, n_2847, n_1148, n_2051, n_109, n_742, n_750, n_2029, n_995, n_454, n_3221, n_2168, n_2790, n_1609, n_374, n_3629, n_3021, n_1989, n_185, n_2359, n_2941, n_396, n_1887, n_3502, n_2523, n_1383, n_3098, n_1073, n_255, n_2346, n_2457, n_662, n_459, n_2312, n_218, n_962, n_3475, n_1215, n_3015, n_1171, n_1578, n_723, n_1920, n_1065, n_1592, n_2536, n_1336, n_2882, n_1721, n_1959, n_1758, n_2338, n_2952, n_2737, n_1574, n_2399, n_3058, n_2812, n_473, n_2048, n_3197, n_3109, n_3607, n_2355, n_2133, n_1921, n_2721, n_1309, n_1878, n_1426, n_1043, n_2585, n_355, n_3505, n_486, n_3002, n_1800, n_1548, n_2725, n_614, n_337, n_1421, n_88, n_2571, n_1286, n_1177, n_3276, n_1355, n_168, n_974, n_2565, n_727, n_1159, n_957, n_773, n_208, n_142, n_2124, n_743, n_3001, n_2081, n_299, n_303, n_3149, n_296, n_613, n_1119, n_2156, n_1240, n_2261, n_1820, n_2729, n_3268, n_3597, n_2418, n_65, n_829, n_2519, n_3354, n_2724, n_1612, n_2179, n_1416, n_2077, n_2897, n_3614, n_2909, n_1724, n_2111, n_2521, n_3301, n_361, n_3466, n_3458, n_700, n_1237, n_573, n_69, n_1420, n_3185, n_1132, n_3330, n_388, n_1366, n_1300, n_2595, n_1127, n_3248, n_2277, n_761, n_2477, n_3523, n_1785, n_1568, n_2829, n_1006, n_3411, n_2110, n_329, n_274, n_1270, n_1664, n_3200, n_1486, n_582, n_3586, n_1332, n_3519, n_2231, n_1390, n_2017, n_73, n_2474, n_2879, n_2604, n_19, n_2090, n_3374, n_3153, n_3045, n_1870, n_309, n_30, n_512, n_2367, n_1591, n_2033, n_84, n_3453, n_130, n_322, n_1682, n_1980, n_2390, n_2628, n_1249, n_3399, n_2896, n_652, n_1111, n_3213, n_1365, n_1927, n_25, n_3065, n_2132, n_1349, n_1093, n_288, n_2400, n_1031, n_263, n_609, n_1041, n_1265, n_3223, n_1909, n_44, n_224, n_3077, n_2681, n_1562, n_383, n_3103, n_834, n_3474, n_112, n_765, n_2255, n_2424, n_2272, n_893, n_1015, n_1140, n_891, n_1651, n_1965, n_239, n_3387, n_630, n_1902, n_2151, n_1941, n_55, n_2106, n_2775, n_2716, n_1913, n_2878, n_504, n_1823, n_511, n_874, n_2464, n_358, n_3422, n_1101, n_2831, n_77, n_102, n_1106, n_1456, n_3557, n_2230, n_3498, n_2015, n_2365, n_1875, n_1982, n_1304, n_2803, n_1324, n_2851, n_987, n_3189, n_1846, n_3037, n_261, n_174, n_2066, n_1885, n_1455, n_3429, n_767, n_993, n_1903, n_2490, n_1407, n_2452, n_1551, n_3154, n_545, n_441, n_860, n_3229, n_450, n_2849, n_1805, n_2176, n_2204, n_2905, n_1816, n_429, n_948, n_3566, n_1217, n_2220, n_2455, n_628, n_365, n_1849, n_2410, n_729, n_1131, n_1084, n_1961, n_970, n_1935, n_911, n_2922, n_1430, n_83, n_3275, n_3499, n_2645, n_2467, n_513, n_3366, n_2727, n_1094, n_1354, n_560, n_1534, n_340, n_2288, n_3421, n_1351, n_2240, n_2696, n_1044, n_1205, n_2436, n_346, n_1209, n_3029, n_1552, n_2508, n_3242, n_3592, n_3618, n_495, n_602, n_3525, n_574, n_2593, n_3486, n_1435, n_879, n_3394, n_16, n_2416, n_58, n_2405, n_623, n_3286, n_2088, n_405, n_2953, n_824, n_359, n_1645, n_2461, n_490, n_1327, n_2858, n_2243, n_996, n_921, n_1684, n_233, n_2658, n_3590, n_1717, n_572, n_366, n_2895, n_815, n_1795, n_2128, n_2578, n_3097, n_3483, n_128, n_1821, n_120, n_2929, n_3424, n_327, n_3478, n_135, n_1381, n_2555, n_2662, n_2740, n_1611, n_1037, n_2368, n_3388, n_2656, n_1080, n_2301, n_1274, n_3583, n_2890, n_3560, n_3059, n_3524, n_2554, n_3465, n_1316, n_1708, n_2419, n_3215, n_426, n_1438, n_1082, n_1840, n_589, n_716, n_1630, n_2122, n_2512, n_3589, n_562, n_1436, n_62, n_3549, n_1691, n_952, n_2786, n_2534, n_2092, n_3171, n_1229, n_391, n_701, n_1437, n_1023, n_2075, n_645, n_539, n_3449, n_803, n_1092, n_2694, n_238, n_1776, n_3559, n_2198, n_2610, n_2661, n_2572, n_2989, n_2281, n_2131, n_2789, n_3026, n_2216, n_531, n_3020, n_1757, n_890, n_1897, n_764, n_1919, n_1056, n_1424, n_162, n_960, n_3462, n_3588, n_2933, n_2308, n_3468, n_1893, n_2910, n_222, n_3419, n_1290, n_1123, n_1467, n_1047, n_2053, n_2163, n_634, n_2328, n_199, n_1958, n_32, n_2254, n_1252, n_348, n_1382, n_1029, n_925, n_3546, n_1206, n_424, n_2647, n_3160, n_1311, n_2191, n_2864, n_2969, n_3195, n_1519, n_256, n_950, n_3190, n_2428, n_1553, n_2664, n_1811, n_2443, n_2624, n_3012, n_3456, n_380, n_419, n_1346, n_3053, n_444, n_1299, n_3244, n_2158, n_1808, n_3290, n_1060, n_1141, n_316, n_2266, n_389, n_3130, n_2465, n_2824, n_3033, n_2650, n_3298, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_3548, n_451, n_619, n_408, n_2440, n_1386, n_1699, n_376, n_3334, n_967, n_1442, n_2923, n_3494, n_2541, n_74, n_1139, n_2731, n_3264, n_515, n_2333, n_57, n_351, n_885, n_2916, n_3166, n_397, n_1432, n_1357, n_483, n_2125, n_683, n_1632, n_3110, n_2998, n_1057, n_1051, n_1085, n_1066, n_721, n_2402, n_1157, n_3073, n_2403, n_841, n_1050, n_22, n_802, n_1954, n_2265, n_46, n_3162, n_1608, n_983, n_1844, n_2760, n_2792, n_3554, n_38, n_3377, n_2870, n_280, n_1305, n_3178, n_873, n_1826, n_378, n_1112, n_3134, n_2304, n_2999, n_762, n_1283, n_1644, n_17, n_2334, n_2637, n_690, n_33, n_1974, n_2463, n_583, n_2086, n_3537, n_2289, n_3080, n_3051, n_302, n_1343, n_2701, n_2783, n_2263, n_3362, n_2881, n_1203, n_1631, n_3282, n_2472, n_821, n_1763, n_2341, n_3105, n_3231, n_1966, n_1768, n_321, n_2294, n_1179, n_621, n_753, n_2475, n_2733, n_455, n_1048, n_1719, n_2993, n_1288, n_212, n_385, n_2785, n_2556, n_507, n_2269, n_2732, n_3569, n_2309, n_2415, n_2948, n_3274, n_3041, n_3299, n_2646, n_1560, n_1605, n_2236, n_330, n_1228, n_2816, n_2123, n_3209, n_972, n_3504, n_692, n_2037, n_2685, n_3040, n_1953, n_1938, n_820, n_1200, n_2499, n_1911, n_3616, n_2460, n_3568, n_2589, n_3203, n_1301, n_1363, n_1668, n_1185, n_991, n_2903, n_3417, n_3482, n_828, n_1967, n_779, n_576, n_1143, n_1579, n_2233, n_1329, n_2743, n_2675, n_3255, n_1312, n_1439, n_804, n_537, n_2827, n_1688, n_3052, n_945, n_2997, n_492, n_3327, n_153, n_1504, n_943, n_3326, n_341, n_3572, n_250, n_992, n_3067, n_1932, n_3375, n_2755, n_543, n_260, n_842, n_650, n_984, n_694, n_3237, n_2082, n_286, n_1992, n_2429, n_1643, n_883, n_1983, n_3167, n_3400, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_3423, n_900, n_2362, n_856, n_2609, n_1793, n_3382, n_1976, n_2223, n_3044, n_3574, n_918, n_3529, n_942, n_2169, n_1804, n_189, n_1147, n_1557, n_1977, n_2153, n_2468, n_1610, n_13, n_1077, n_1422, n_3196, n_3078, n_2364, n_2533, n_540, n_3492, n_618, n_3094, n_896, n_2310, n_2780, n_323, n_2287, n_2860, n_3316, n_195, n_356, n_2291, n_3099, n_2596, n_894, n_1636, n_2056, n_3253, n_1730, n_3601, n_3603, n_831, n_2280, n_2192, n_964, n_3363, n_1373, n_1350, n_1511, n_1865, n_2973, n_1470, n_1096, n_2094, n_2670, n_234, n_1575, n_1697, n_1735, n_833, n_2318, n_2393, n_2020, n_5, n_1646, n_2502, n_225, n_2504, n_1307, n_1881, n_2974, n_988, n_2749, n_2043, n_2901, n_1940, n_814, n_2707, n_2751, n_2793, n_3372, n_3451, n_192, n_2971, n_3442, n_1549, n_1934, n_2311, n_1201, n_1114, n_655, n_3240, n_2025, n_1616, n_1446, n_2285, n_3147, n_2758, n_669, n_472, n_1458, n_1176, n_1472, n_2298, n_2471, n_1807, n_387, n_1149, n_2618, n_398, n_1671, n_635, n_2559, n_763, n_3230, n_1020, n_1062, n_3342, n_211, n_2303, n_1824, n_1917, n_2295, n_1219, n_3386, n_3, n_1204, n_2840, n_2810, n_2325, n_178, n_2747, n_2446, n_3488, n_1814, n_1035, n_2822, n_287, n_555, n_783, n_1848, n_1928, n_2126, n_2893, n_1188, n_2588, n_2962, n_1722, n_661, n_2441, n_41, n_1802, n_3083, n_2600, n_849, n_2795, n_15, n_336, n_584, n_681, n_1638, n_1786, n_2981, n_50, n_430, n_2002, n_2282, n_3608, n_510, n_2800, n_216, n_2371, n_2935, n_311, n_3233, n_3380, n_3177, n_830, n_2098, n_1296, n_2627, n_3409, n_3460, n_2352, n_3538, n_1413, n_801, n_2207, n_2080, n_2377, n_2619, n_2340, n_3085, n_2444, n_2068, n_241, n_3552, n_875, n_357, n_1110, n_1655, n_445, n_2641, n_3198, n_749, n_1895, n_3123, n_3137, n_2574, n_1134, n_1358, n_717, n_165, n_939, n_482, n_2361, n_1088, n_588, n_1173, n_789, n_3393, n_1232, n_1603, n_734, n_638, n_2638, n_866, n_107, n_969, n_1401, n_3520, n_2492, n_1019, n_1105, n_249, n_1998, n_304, n_1338, n_577, n_2016, n_1522, n_2949, n_1687, n_1637, n_2034, n_1419, n_2711, n_338, n_149, n_1653, n_693, n_2270, n_1506, n_3206, n_2653, n_3578, n_14, n_836, n_990, n_2867, n_2496, n_1886, n_1389, n_1894, n_975, n_1908, n_1256, n_1702, n_2259, n_2794, n_567, n_1465, n_3145, n_3124, n_778, n_1122, n_151, n_3192, n_2608, n_306, n_2657, n_458, n_770, n_2995, n_1375, n_2494, n_3547, n_2649, n_1102, n_2852, n_2392, n_3459, n_3093, n_1843, n_711, n_1499, n_3061, n_3155, n_85, n_1187, n_3517, n_2633, n_1441, n_3100, n_2522, n_2435, n_1392, n_1597, n_1929, n_2807, n_1164, n_1659, n_1834, n_2097, n_2313, n_2542, n_489, n_1174, n_2431, n_3324, n_3356, n_2835, n_2558, n_1371, n_617, n_1303, n_2206, n_2063, n_3182, n_1572, n_1968, n_3269, n_2564, n_2252, n_876, n_1516, n_1190, n_3506, n_1736, n_3605, n_1685, n_118, n_2409, n_601, n_917, n_3450, n_1714, n_966, n_253, n_1116, n_2000, n_1661, n_3402, n_1212, n_2074, n_1541, n_2576, n_3565, n_172, n_206, n_217, n_726, n_3174, n_982, n_2575, n_2988, n_3390, n_1573, n_1453, n_1731, n_2217, n_818, n_2373, n_1970, n_861, n_1713, n_1183, n_3398, n_2307, n_2766, n_1658, n_899, n_1253, n_210, n_1737, n_2201, n_2722, n_2117, n_2745, n_3408, n_1904, n_2640, n_1993, n_774, n_1628, n_2493, n_2205, n_3432, n_1335, n_1514, n_1777, n_1957, n_1059, n_1345, n_176, n_1133, n_1771, n_1912, n_3401, n_1899, n_3226, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_3090, n_2067, n_527, n_1168, n_707, n_2219, n_2437, n_2885, n_3533, n_2877, n_3318, n_2148, n_937, n_2445, n_1427, n_2779, n_3485, n_393, n_108, n_487, n_1584, n_665, n_1726, n_1835, n_3035, n_66, n_1440, n_177, n_2164, n_421, n_1988, n_3333, n_2115, n_1853, n_1356, n_2845, n_1787, n_2634, n_910, n_2232, n_3034, n_2212, n_2602, n_1657, n_768, n_1475, n_1302, n_1774, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_2811, n_1496, n_3348, n_179, n_1125, n_125, n_410, n_2547, n_3014, n_708, n_529, n_1812, n_735, n_2501, n_3079, n_232, n_1915, n_1109, n_126, n_895, n_2532, n_1310, n_2605, n_3358, n_2121, n_1803, n_202, n_3308, n_2665, n_427, n_1399, n_1543, n_1991, n_1979, n_791, n_732, n_1533, n_2224, n_193, n_3368, n_2924, n_3467, n_808, n_2484, n_797, n_3530, n_1025, n_1930, n_1955, n_2765, n_3329, n_500, n_2994, n_1067, n_2946, n_1720, n_148, n_2830, n_2401, n_3135, n_435, n_2003, n_159, n_766, n_1457, n_541, n_2692, n_3573, n_3148, n_538, n_2354, n_2246, n_2008, n_1117, n_799, n_2264, n_2754, n_687, n_3534, n_715, n_1742, n_1480, n_1482, n_1213, n_2489, n_1266, n_536, n_3438, n_872, n_2012, n_594, n_200, n_1291, n_3381, n_3503, n_1297, n_1753, n_2283, n_2866, n_3278, n_1782, n_2245, n_3561, n_1155, n_1418, n_89, n_1972, n_1524, n_1689, n_1485, n_2806, n_115, n_1011, n_1184, n_2184, n_985, n_1855, n_2425, n_2917, n_869, n_810, n_2965, n_3536, n_416, n_827, n_3217, n_3404, n_3425, n_401, n_1703, n_3312, n_1352, n_2926, n_626, n_2197, n_2199, n_3540, n_1650, n_1144, n_1137, n_1570, n_2814, n_3046, n_1170, n_305, n_2023, n_2213, n_3249, n_3211, n_3285, n_2351, n_2211, n_2095, n_3121, n_137, n_676, n_294, n_318, n_2103, n_653, n_2160, n_642, n_3337, n_2228, n_2527, n_1602, n_2498, n_194, n_855, n_1178, n_1461, n_2697, n_850, n_684, n_3074, n_124, n_3204, n_268, n_2421, n_2286, n_2902, n_664, n_1999, n_503, n_2372, n_2065, n_2136, n_2480, n_235, n_1372, n_2861, n_605, n_2630, n_1273, n_1822, n_3397, n_353, n_620, n_643, n_2363, n_2430, n_916, n_1081, n_2549, n_493, n_2705, n_3005, n_2332, n_1235, n_703, n_698, n_980, n_1115, n_2433, n_3293, n_3129, n_1282, n_1318, n_1783, n_780, n_2977, n_3606, n_2601, n_3043, n_998, n_2375, n_2550, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_1907, n_3600, n_501, n_823, n_245, n_2686, n_2528, n_725, n_2344, n_1388, n_1417, n_1295, n_2836, n_2316, n_672, n_1985, n_3055, n_1898, n_2107, n_3294, n_3219, n_3315, n_581, n_2906, n_382, n_554, n_1625, n_2130, n_3415, n_2187, n_2284, n_898, n_2817, n_3172, n_3139, n_2773, n_3239, n_3292, n_2598, n_1762, n_1013, n_3365, n_3476, n_1452, n_718, n_2687, n_265, n_3023, n_3553, n_1120, n_719, n_443, n_1791, n_198, n_1890, n_1747, n_714, n_2850, n_1683, n_1817, n_909, n_1944, n_1497, n_1530, n_2654, n_997, n_3431, n_3104, n_932, n_3169, n_3151, n_612, n_3131, n_2078, n_1409, n_788, n_1326, n_3070, n_3284, n_119, n_3176, n_2884, n_1268, n_2996, n_559, n_825, n_2819, n_3126, n_1981, n_508, n_2186, n_506, n_1320, n_1663, n_737, n_1718, n_3609, n_986, n_2315, n_509, n_3228, n_1317, n_147, n_1518, n_1715, n_2102, n_3581, n_2562, n_1281, n_67, n_1952, n_1192, n_2221, n_1024, n_3576, n_1063, n_1889, n_209, n_1792, n_1564, n_1868, n_1613, n_733, n_1489, n_1922, n_2966, n_1376, n_941, n_2326, n_981, n_2560, n_1569, n_2188, n_68, n_3495, n_867, n_186, n_2348, n_2422, n_134, n_2239, n_587, n_2950, n_63, n_792, n_756, n_1429, n_399, n_1238, n_2448, n_3140, n_548, n_3170, n_812, n_298, n_2104, n_2748, n_3311, n_518, n_505, n_2057, n_3272, n_3011, n_1772, n_282, n_752, n_905, n_1476, n_1108, n_2898, n_782, n_2717, n_2818, n_1100, n_1861, n_2129, n_1395, n_3345, n_862, n_3584, n_1425, n_760, n_1901, n_3069, n_1900, n_1620, n_3032, n_381, n_3628, n_2889, n_220, n_390, n_1330, n_1867, n_31, n_1945, n_2772, n_481, n_3018, n_1675, n_3072, n_1924, n_2573, n_3084, n_3081, n_3313, n_1727, n_2710, n_1554, n_2939, n_1745, n_2735, n_769, n_2497, n_2006, n_3412, n_42, n_2844, n_1995, n_2411, n_2138, n_1046, n_271, n_934, n_1618, n_2260, n_826, n_2343, n_1813, n_2447, n_886, n_3439, n_2014, n_3056, n_1221, n_2345, n_2986, n_654, n_1172, n_167, n_2535, n_379, n_428, n_1341, n_2726, n_570, n_2774, n_3295, n_1641, n_1361, n_3184, n_2382, n_1707, n_853, n_3062, n_3161, n_377, n_2317, n_751, n_3289, n_2799, n_2172, n_1973, n_786, n_1083, n_1142, n_2376, n_2488, n_1129, n_392, n_2579, n_3477, n_3017, n_158, n_3626, n_2476, n_704, n_787, n_1770, n_138, n_2781, n_2456, n_961, n_2250, n_2678, n_1756, n_771, n_2778, n_276, n_95, n_1716, n_2788, n_2872, n_1225, n_2984, n_1520, n_2451, n_169, n_2887, n_522, n_3364, n_1287, n_1262, n_2691, n_400, n_930, n_181, n_1873, n_1411, n_3201, n_3054, n_221, n_622, n_1962, n_1577, n_2423, n_1087, n_3472, n_2526, n_2854, n_386, n_994, n_1701, n_3344, n_2194, n_848, n_1550, n_2874, n_2764, n_2703, n_1498, n_2167, n_3302, n_3235, n_1223, n_1272, n_2680, n_3391, n_104, n_682, n_1567, n_56, n_141, n_2567, n_3543, n_1247, n_2709, n_3102, n_922, n_3122, n_816, n_1648, n_591, n_145, n_1536, n_3050, n_3265, n_1857, n_1344, n_2041, n_313, n_631, n_3627, n_479, n_1246, n_1339, n_1478, n_1797, n_432, n_1769, n_2957, n_839, n_3551, n_1210, n_3518, n_2964, n_1364, n_2956, n_2357, n_2183, n_2673, n_2742, n_3314, n_2360, n_3254, n_328, n_140, n_2292, n_1250, n_2173, n_369, n_1842, n_871, n_2442, n_3309, n_598, n_685, n_928, n_608, n_1367, n_78, n_1943, n_1460, n_772, n_2018, n_3464, n_3260, n_1555, n_3117, n_2834, n_3245, n_3357, n_499, n_2531, n_1589, n_517, n_3428, n_98, n_2961, n_402, n_413, n_1086, n_2570, n_2702, n_796, n_1858, n_3351, n_1619, n_3527, n_2815, n_236, n_2119, n_1502, n_2157, n_2552, n_1469, n_1012, n_1, n_1396, n_2744, n_1348, n_2030, n_903, n_2453, n_1525, n_1752, n_2397, n_740, n_2883, n_3115, n_203, n_3509, n_3352, n_384, n_2208, n_3076, n_1404, n_80, n_3063, n_3617, n_2912, n_1794, n_3535, n_2182, n_35, n_1315, n_2234, n_277, n_1061, n_3251, n_92, n_1910, n_333, n_1298, n_2931, n_1652, n_2209, n_462, n_2050, n_2809, n_1193, n_2797, n_1676, n_1255, n_258, n_1113, n_3118, n_29, n_79, n_3227, n_3300, n_2321, n_3511, n_1226, n_722, n_1277, n_2591, n_3443, n_188, n_2146, n_844, n_201, n_3384, n_471, n_852, n_3497, n_1487, n_40, n_1864, n_1028, n_1601, n_3336, n_781, n_474, n_2940, n_542, n_3435, n_3521, n_463, n_3575, n_1546, n_595, n_502, n_3562, n_466, n_2612, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_2841, n_3165, n_1627, n_2918, n_3232, n_3322, n_1245, n_846, n_2427, n_2438, n_2505, n_1673, n_465, n_2832, n_76, n_362, n_1321, n_170, n_1975, n_27, n_2296, n_2070, n_161, n_273, n_1937, n_585, n_2112, n_3250, n_1739, n_3181, n_270, n_2958, n_616, n_2278, n_81, n_2594, n_3114, n_3125, n_2394, n_3234, n_1914, n_3612, n_2954, n_2135, n_2335, n_2904, n_3493, n_745, n_2381, n_3303, n_1654, n_3004, n_3323, n_2569, n_3112, n_2349, n_1103, n_3132, n_3556, n_648, n_1379, n_2734, n_312, n_2196, n_3591, n_3024, n_2170, n_1076, n_2823, n_1091, n_1408, n_3512, n_494, n_1761, n_641, n_3238, n_3210, n_730, n_3175, n_3522, n_2036, n_1325, n_3267, n_1595, n_2161, n_354, n_575, n_480, n_425, n_795, n_2404, n_2083, n_695, n_180, n_3281, n_656, n_3307, n_1606, n_2503, n_1220, n_37, n_1694, n_1540, n_3266, n_2485, n_229, n_1936, n_1956, n_437, n_1642, n_2279, n_3373, n_2655, n_2027, n_60, n_403, n_453, n_2642, n_1130, n_720, n_0, n_2500, n_2366, n_1918, n_1526, n_863, n_2210, n_805, n_3247, n_1604, n_1275, n_2513, n_2525, n_3091, n_2695, n_1764, n_3480, n_2892, n_3057, n_3194, n_3582, n_3066, n_113, n_712, n_2414, n_2907, n_246, n_1583, n_2426, n_2826, n_3577, n_3539, n_1042, n_1402, n_2820, n_269, n_2049, n_2273, n_285, n_412, n_2719, n_1493, n_657, n_644, n_1741, n_2229, n_1160, n_1397, n_491, n_1258, n_1074, n_3347, n_2004, n_3216, n_1621, n_2708, n_2113, n_251, n_160, n_566, n_565, n_2586, n_1448, n_2225, n_3567, n_3613, n_1507, n_1398, n_2383, n_1879, n_597, n_1996, n_3406, n_3604, n_3444, n_1181, n_1505, n_1634, n_1196, n_2019, n_651, n_1340, n_2274, n_2972, n_334, n_811, n_1558, n_3225, n_807, n_3321, n_2166, n_2938, n_3212, n_835, n_175, n_666, n_3319, n_262, n_1433, n_3594, n_1704, n_2256, n_3152, n_3335, n_99, n_1254, n_1026, n_3413, n_2026, n_1969, n_1234, n_2109, n_319, n_364, n_1138, n_927, n_20, n_1089, n_2013, n_1990, n_2044, n_2689, n_2920, n_3259, n_1004, n_1186, n_1032, n_242, n_2614, n_2511, n_1681, n_2010, n_2991, n_3383, n_1018, n_2242, n_2247, n_2752, n_2894, n_3016, n_1693, n_3585, n_2975, n_3473, n_438, n_2599, n_713, n_2704, n_904, n_2839, n_3338, n_1588, n_1622, n_2237, n_3414, n_3463, n_166, n_1180, n_1827, n_3360, n_2524, n_1271, n_2802, n_533, n_1542, n_1251, n_3159, n_278, n_2728, n_2268, n_15103);

input n_924;
input n_1263;
input n_3304;
input n_977;
input n_1378;
input n_2253;
input n_2417;
input n_611;
input n_2756;
input n_1126;
input n_1423;
input n_1729;
input n_2739;
input n_1166;
input n_2380;
input n_1751;
input n_469;
input n_1508;
input n_82;
input n_2771;
input n_785;
input n_3241;
input n_549;
input n_2617;
input n_2200;
input n_3261;
input n_3006;
input n_532;
input n_1161;
input n_3027;
input n_1859;
input n_2746;
input n_1677;
input n_1150;
input n_2327;
input n_3179;
input n_3127;
input n_226;
input n_1780;
input n_3256;
input n_1488;
input n_667;
input n_2899;
input n_2955;
input n_790;
input n_3619;
input n_1055;
input n_3541;
input n_3622;
input n_2386;
input n_3596;
input n_1501;
input n_111;
input n_2395;
input n_880;
input n_3086;
input n_3297;
input n_544;
input n_1007;
input n_2369;
input n_155;
input n_2927;
input n_552;
input n_1528;
input n_2683;
input n_1370;
input n_1292;
input n_2347;
input n_2520;
input n_2821;
input n_1198;
input n_1360;
input n_2388;
input n_1099;
input n_2568;
input n_956;
input n_564;
input n_423;
input n_1738;
input n_2021;
input n_21;
input n_2134;
input n_3064;
input n_2391;
input n_105;
input n_3088;
input n_1021;
input n_1960;
input n_2843;
input n_2185;
input n_4;
input n_3270;
input n_551;
input n_2143;
input n_2853;
input n_3615;
input n_2059;
input n_1323;
input n_1466;
input n_688;
input n_1695;
input n_2487;
input n_1353;
input n_800;
input n_3595;
input n_3246;
input n_3202;
input n_1347;
input n_2495;
input n_2880;
input n_1535;
input n_1789;
input n_1666;
input n_3350;
input n_2389;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_2302;
input n_915;
input n_1545;
input n_2374;
input n_864;
input n_173;
input n_859;
input n_951;
input n_3341;
input n_1947;
input n_1264;
input n_3587;
input n_2114;
input n_3445;
input n_447;
input n_247;
input n_2001;
input n_1494;
input n_3407;
input n_3571;
input n_3599;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1799;
input n_2069;
input n_2396;
input n_3621;
input n_1580;
input n_674;
input n_417;
input n_1939;
input n_2486;
input n_3434;
input n_1806;
input n_516;
input n_933;
input n_2244;
input n_2257;
input n_1152;
input n_3501;
input n_3448;
input n_497;
input n_1869;
input n_1607;
input n_1563;
input n_606;
input n_3019;
input n_275;
input n_3039;
input n_2011;
input n_2096;
input n_26;
input n_877;
input n_2105;
input n_2538;
input n_2024;
input n_2;
input n_2530;
input n_1696;
input n_2483;
input n_3163;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1860;
input n_2543;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_2031;
input n_2076;
input n_2482;
input n_3036;
input n_2677;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_1896;
input n_2165;
input n_2147;
input n_929;
input n_3010;
input n_3180;
input n_3379;
input n_3532;
input n_2770;
input n_1124;
input n_1818;
input n_2127;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_2584;
input n_1257;
input n_2639;
input n_171;
input n_1182;
input n_3188;
input n_3325;
input n_3107;
input n_3531;
input n_3403;
input n_579;
input n_1698;
input n_1261;
input n_2329;
input n_938;
input n_1098;
input n_2963;
input n_3624;
input n_2142;
input n_3186;
input n_3461;
input n_3082;
input n_320;
input n_1154;
input n_2189;
input n_3332;
input n_1242;
input n_3283;
input n_1135;
input n_3048;
input n_3258;
input n_24;
input n_406;
input n_519;
input n_2323;
input n_2203;
input n_2597;
input n_1016;
input n_1243;
input n_546;
input n_2959;
input n_101;
input n_3340;
input n_2047;
input n_1280;
input n_3277;
input n_1845;
input n_281;
input n_240;
input n_2052;
input n_2193;
input n_2978;
input n_2058;
input n_2458;
input n_2478;
input n_291;
input n_231;
input n_257;
input n_2761;
input n_731;
input n_371;
input n_1483;
input n_2888;
input n_1314;
input n_1512;
input n_3157;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_2537;
input n_2983;
input n_569;
input n_2669;
input n_2144;
input n_1778;
input n_3214;
input n_227;
input n_2306;
input n_920;
input n_2515;
input n_3022;
input n_1289;
input n_1517;
input n_2091;
input n_2466;
input n_2635;
input n_2652;
input n_94;
input n_335;
input n_3631;
input n_2715;
input n_3087;
input n_2085;
input n_3489;
input n_1669;
input n_2566;
input n_370;
input n_976;
input n_1949;
input n_343;
input n_1449;
input n_308;
input n_1946;
input n_2936;
input n_1566;
input n_2032;
input n_297;
input n_2587;
input n_156;
input n_2149;
input n_1078;
input n_2782;
input n_1670;
input n_2672;
input n_775;
input n_219;
input n_3060;
input n_157;
input n_2651;
input n_3490;
input n_600;
input n_1484;
input n_2071;
input n_2561;
input n_1374;
input n_1328;
input n_2643;
input n_223;
input n_2141;
input n_1948;
input n_3013;
input n_3183;
input n_1984;
input n_3437;
input n_2099;
input n_2408;
input n_3446;
input n_3353;
input n_264;
input n_1877;
input n_1831;
input n_1598;
input n_3049;
input n_1723;
input n_955;
input n_1850;
input n_163;
input n_3028;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_2384;
input n_1036;
input n_1097;
input n_1749;
input n_347;
input n_3156;
input n_59;
input n_550;
input n_696;
input n_3101;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_3376;
input n_646;
input n_1428;
input n_2663;
input n_436;
input n_1394;
input n_2659;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_2693;
input n_1040;
input n_2202;
input n_2648;
input n_1872;
input n_3389;
input n_1852;
input n_2159;
input n_578;
input n_2976;
input n_926;
input n_2180;
input n_2249;
input n_344;
input n_2353;
input n_1218;
input n_1931;
input n_2439;
input n_2632;
input n_2276;
input n_3089;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_2089;
input n_3420;
input n_1030;
input n_72;
input n_2470;
input n_1755;
input n_3222;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1801;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_2908;
input n_2970;
input n_3361;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_2235;
input n_1862;
input n_673;
input n_837;
input n_1239;
input n_2915;
input n_528;
input n_2300;
input n_2791;
input n_1796;
input n_2551;
input n_3291;
input n_680;
input n_1473;
input n_1587;
input n_2682;
input n_395;
input n_164;
input n_553;
input n_901;
input n_2432;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_3440;
input n_3405;
input n_214;
input n_2174;
input n_2714;
input n_1748;
input n_3563;
input n_2934;
input n_1672;
input n_2506;
input n_675;
input n_2699;
input n_888;
input n_1880;
input n_2769;
input n_3542;
input n_2337;
input n_3436;
input n_1167;
input n_1626;
input n_3550;
input n_637;
input n_2615;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1863;
input n_1064;
input n_144;
input n_858;
input n_2079;
input n_2238;
input n_114;
input n_96;
input n_923;
input n_2118;
input n_691;
input n_1151;
input n_2985;
input n_2944;
input n_881;
input n_1405;
input n_2407;
input n_1706;
input n_468;
input n_3418;
input n_213;
input n_129;
input n_342;
input n_2932;
input n_2753;
input n_464;
input n_2980;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_3306;
input n_1784;
input n_2859;
input n_2842;
input n_1075;
input n_3262;
input n_3136;
input n_1836;
input n_2868;
input n_3395;
input n_1450;
input n_3141;
input n_1322;
input n_2101;
input n_1471;
input n_1986;
input n_2863;
input n_2072;
input n_3164;
input n_2738;
input n_1750;
input n_3570;
input n_1459;
input n_460;
input n_889;
input n_2358;
input n_973;
input n_2968;
input n_1700;
input n_2833;
input n_477;
input n_3191;
input n_571;
input n_1585;
input n_461;
input n_2684;
input n_2712;
input n_3593;
input n_3193;
input n_1971;
input n_1599;
input n_3252;
input n_2275;
input n_2855;
input n_3507;
input n_3273;
input n_2713;
input n_3544;
input n_2644;
input n_2700;
input n_1211;
input n_1197;
input n_3367;
input n_2951;
input n_1523;
input n_2730;
input n_1950;
input n_3008;
input n_907;
input n_1447;
input n_2251;
input n_3096;
input n_1377;
input n_2370;
input n_190;
input n_3496;
input n_989;
input n_2544;
input n_1039;
input n_2214;
input n_3339;
input n_34;
input n_2055;
input n_3427;
input n_228;
input n_283;
input n_3025;
input n_3349;
input n_1403;
input n_2248;
input n_2356;
input n_488;
input n_736;
input n_892;
input n_3320;
input n_3007;
input n_2688;
input n_1000;
input n_1202;
input n_2750;
input n_2620;
input n_1278;
input n_2622;
input n_2062;
input n_2668;
input n_1002;
input n_1463;
input n_1581;
input n_2100;
input n_49;
input n_3071;
input n_310;
input n_3310;
input n_54;
input n_593;
input n_3487;
input n_2258;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_3359;
input n_838;
input n_2784;
input n_2919;
input n_332;
input n_3092;
input n_1053;
input n_3470;
input n_1224;
input n_2865;
input n_349;
input n_2557;
input n_1926;
input n_2706;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_2150;
input n_3146;
input n_2241;
input n_2757;
input n_2152;
input n_3598;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_2590;
input n_2776;
input n_2140;
input n_2385;
input n_3580;
input n_1819;
input n_2330;
input n_2139;
input n_2942;
input n_476;
input n_2987;
input n_1527;
input n_2042;
input n_534;
input n_3106;
input n_1882;
input n_884;
input n_3328;
input n_345;
input n_944;
input n_1754;
input n_3611;
input n_1623;
input n_2862;
input n_2175;
input n_2921;
input n_2720;
input n_2324;
input n_1854;
input n_91;
input n_2606;
input n_2674;
input n_3187;
input n_1565;
input n_3508;
input n_2828;
input n_3371;
input n_1809;
input n_1856;
input n_182;
input n_143;
input n_647;
input n_3433;
input n_237;
input n_407;
input n_1072;
input n_2218;
input n_2267;
input n_832;
input n_857;
input n_2305;
input n_3392;
input n_3430;
input n_2636;
input n_2450;
input n_3208;
input n_207;
input n_561;
input n_1319;
input n_2379;
input n_3331;
input n_3447;
input n_2616;
input n_2911;
input n_3305;
input n_2154;
input n_1825;
input n_1951;
input n_1883;
input n_1906;
input n_2759;
input n_1712;
input n_1387;
input n_3528;
input n_2262;
input n_2462;
input n_2514;
input n_1532;
input n_2322;
input n_2271;
input n_2625;
input n_18;
input n_3257;
input n_3625;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_2798;
input n_2331;
input n_2945;
input n_2293;
input n_686;
input n_2837;
input n_847;
input n_1393;
input n_2319;
input n_596;
input n_1775;
input n_2979;
input n_3296;
input n_2028;
input n_1368;
input n_3481;
input n_2762;
input n_558;
input n_2808;
input n_702;
input n_1276;
input n_3009;
input n_2548;
input n_822;
input n_1412;
input n_2676;
input n_1709;
input n_2679;
input n_2108;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_2930;
input n_1838;
input n_1199;
input n_1847;
input n_1779;
input n_2767;
input n_2777;
input n_2603;
input n_3514;
input n_3116;
input n_352;
input n_1884;
input n_2434;
input n_2660;
input n_53;
input n_3602;
input n_1038;
input n_2967;
input n_520;
input n_1369;
input n_409;
input n_2611;
input n_1841;
input n_1660;
input n_887;
input n_1905;
input n_2553;
input n_154;
input n_3207;
input n_2581;
input n_71;
input n_2195;
input n_2529;
input n_3224;
input n_300;
input n_2698;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1891;
input n_1481;
input n_2626;
input n_3441;
input n_3042;
input n_1942;
input n_434;
input n_1978;
input n_1544;
input n_2510;
input n_3047;
input n_3526;
input n_868;
input n_2454;
input n_639;
input n_2804;
input n_914;
input n_2120;
input n_411;
input n_414;
input n_2546;
input n_1629;
input n_1293;
input n_2801;
input n_3120;
input n_965;
input n_1876;
input n_1743;
input n_3491;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_2763;
input n_360;
input n_36;
input n_1479;
input n_1810;
input n_2350;
input n_2813;
input n_64;
input n_2825;
input n_1888;
input n_2009;
input n_759;
input n_2222;
input n_1892;
input n_3510;
input n_28;
input n_806;
input n_2990;
input n_1997;
input n_2667;
input n_1766;
input n_3218;
input n_1477;
input n_3142;
input n_324;
input n_1635;
input n_1963;
input n_2226;
input n_1571;
input n_2891;
input n_3119;
input n_187;
input n_1189;
input n_2690;
input n_103;
input n_97;
input n_3370;
input n_11;
input n_2215;
input n_3479;
input n_7;
input n_1259;
input n_1690;
input n_706;
input n_746;
input n_1649;
input n_3150;
input n_747;
input n_2064;
input n_52;
input n_784;
input n_110;
input n_2449;
input n_1733;
input n_1244;
input n_3500;
input n_2413;
input n_431;
input n_1194;
input n_1925;
input n_2297;
input n_1815;
input n_3279;
input n_2621;
input n_615;
input n_851;
input n_1759;
input n_843;
input n_1788;
input n_2177;
input n_2491;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_2227;
input n_678;
input n_2671;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_2190;
input n_3346;
input n_776;
input n_1798;
input n_2022;
input n_1790;
input n_2518;
input n_2876;
input n_1415;
input n_367;
input n_2629;
input n_2592;
input n_3416;
input n_452;
input n_525;
input n_3484;
input n_3620;
input n_1260;
input n_1746;
input n_1647;
input n_2181;
input n_2479;
input n_2838;
input n_1829;
input n_1464;
input n_3133;
input n_3513;
input n_649;
input n_547;
input n_2563;
input n_43;
input n_1444;
input n_1191;
input n_2387;
input n_2992;
input n_1674;
input n_1833;
input n_116;
input n_3138;
input n_1830;
input n_2517;
input n_2073;
input n_1710;
input n_284;
input n_1128;
input n_2928;
input n_3128;
input n_139;
input n_1734;
input n_3038;
input n_744;
input n_590;
input n_629;
input n_2631;
input n_1308;
input n_2871;
input n_2178;
input n_3068;
input n_1767;
input n_3144;
input n_2943;
input n_2913;
input n_2336;
input n_3143;
input n_3168;
input n_254;
input n_1680;
input n_1233;
input n_3469;
input n_2607;
input n_23;
input n_1615;
input n_1529;
input n_2005;
input n_526;
input n_1916;
input n_3317;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_2469;
input n_1121;
input n_2723;
input n_3355;
input n_314;
input n_368;
input n_433;
input n_604;
input n_2007;
input n_8;
input n_3220;
input n_949;
input n_2539;
input n_3263;
input n_100;
input n_2582;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_2736;
input n_1001;
input n_1503;
input n_2054;
input n_498;
input n_1468;
input n_1559;
input n_1765;
input n_3455;
input n_1866;
input n_689;
input n_3158;
input n_738;
input n_1624;
input n_3000;
input n_640;
input n_3452;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1744;
input n_2623;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1994;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_3108;
input n_3113;
input n_3111;
input n_2718;
input n_1195;
input n_1837;
input n_1839;
input n_610;
input n_2577;
input n_1760;
input n_2875;
input n_936;
input n_568;
input n_1500;
input n_2960;
input n_39;
input n_1090;
input n_2796;
input n_757;
input n_3280;
input n_2342;
input n_633;
input n_2856;
input n_439;
input n_3471;
input n_106;
input n_1832;
input n_259;
input n_448;
input n_1851;
input n_758;
input n_999;
input n_3205;
input n_2046;
input n_2848;
input n_2741;
input n_2937;
input n_3003;
input n_3610;
input n_1933;
input n_2290;
input n_93;
input n_1656;
input n_3564;
input n_3288;
input n_1158;
input n_3095;
input n_2045;
input n_3369;
input n_1509;
input n_1874;
input n_2040;
input n_563;
input n_2060;
input n_3199;
input n_2613;
input n_1987;
input n_2805;
input n_1145;
input n_878;
input n_524;
input n_3457;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_2145;
input n_741;
input n_1639;
input n_1306;
input n_1068;
input n_3030;
input n_3558;
input n_1871;
input n_2580;
input n_3630;
input n_2545;
input n_2787;
input n_2914;
input n_1964;
input n_2869;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_3271;
input n_2039;
input n_1207;
input n_919;
input n_908;
input n_2412;
input n_2406;
input n_3623;
input n_90;
input n_2846;
input n_724;
input n_1781;
input n_2084;
input n_2925;
input n_2035;
input n_658;
input n_2061;
input n_3555;
input n_3579;
input n_3075;
input n_3173;
input n_2378;
input n_2509;
input n_1740;
input n_3236;
input n_2398;
input n_1362;
input n_2857;
input n_1586;
input n_456;
input n_959;
input n_2459;
input n_3031;
input n_535;
input n_152;
input n_3396;
input n_940;
input n_1445;
input n_9;
input n_3516;
input n_1492;
input n_2155;
input n_2516;
input n_1923;
input n_1773;
input n_592;
input n_3243;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_2666;
input n_2982;
input n_3385;
input n_1017;
input n_2481;
input n_2947;
input n_3545;
input n_2171;
input n_123;
input n_978;
input n_2768;
input n_2116;
input n_2314;
input n_1434;
input n_1054;
input n_2507;
input n_1474;
input n_1665;
input n_1269;
input n_2420;
input n_2900;
input n_1095;
input n_3343;
input n_3515;
input n_1828;
input n_1614;
input n_2886;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_2093;
input n_2038;
input n_2320;
input n_2339;
input n_2473;
input n_3287;
input n_2137;
input n_3378;
input n_603;
input n_1431;
input n_2583;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_3426;
input n_3454;
input n_2299;
input n_131;
input n_2540;
input n_2873;
input n_636;
input n_660;
input n_3410;
input n_2087;
input n_1640;
input n_2162;
input n_1732;
input n_1009;
input n_2847;
input n_1148;
input n_2051;
input n_109;
input n_742;
input n_750;
input n_2029;
input n_995;
input n_454;
input n_3221;
input n_2168;
input n_2790;
input n_1609;
input n_374;
input n_3629;
input n_3021;
input n_1989;
input n_185;
input n_2359;
input n_2941;
input n_396;
input n_1887;
input n_3502;
input n_2523;
input n_1383;
input n_3098;
input n_1073;
input n_255;
input n_2346;
input n_2457;
input n_662;
input n_459;
input n_2312;
input n_218;
input n_962;
input n_3475;
input n_1215;
input n_3015;
input n_1171;
input n_1578;
input n_723;
input n_1920;
input n_1065;
input n_1592;
input n_2536;
input n_1336;
input n_2882;
input n_1721;
input n_1959;
input n_1758;
input n_2338;
input n_2952;
input n_2737;
input n_1574;
input n_2399;
input n_3058;
input n_2812;
input n_473;
input n_2048;
input n_3197;
input n_3109;
input n_3607;
input n_2355;
input n_2133;
input n_1921;
input n_2721;
input n_1309;
input n_1878;
input n_1426;
input n_1043;
input n_2585;
input n_355;
input n_3505;
input n_486;
input n_3002;
input n_1800;
input n_1548;
input n_2725;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_2571;
input n_1286;
input n_1177;
input n_3276;
input n_1355;
input n_168;
input n_974;
input n_2565;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_2124;
input n_743;
input n_3001;
input n_2081;
input n_299;
input n_303;
input n_3149;
input n_296;
input n_613;
input n_1119;
input n_2156;
input n_1240;
input n_2261;
input n_1820;
input n_2729;
input n_3268;
input n_3597;
input n_2418;
input n_65;
input n_829;
input n_2519;
input n_3354;
input n_2724;
input n_1612;
input n_2179;
input n_1416;
input n_2077;
input n_2897;
input n_3614;
input n_2909;
input n_1724;
input n_2111;
input n_2521;
input n_3301;
input n_361;
input n_3466;
input n_3458;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_3185;
input n_1132;
input n_3330;
input n_388;
input n_1366;
input n_1300;
input n_2595;
input n_1127;
input n_3248;
input n_2277;
input n_761;
input n_2477;
input n_3523;
input n_1785;
input n_1568;
input n_2829;
input n_1006;
input n_3411;
input n_2110;
input n_329;
input n_274;
input n_1270;
input n_1664;
input n_3200;
input n_1486;
input n_582;
input n_3586;
input n_1332;
input n_3519;
input n_2231;
input n_1390;
input n_2017;
input n_73;
input n_2474;
input n_2879;
input n_2604;
input n_19;
input n_2090;
input n_3374;
input n_3153;
input n_3045;
input n_1870;
input n_309;
input n_30;
input n_512;
input n_2367;
input n_1591;
input n_2033;
input n_84;
input n_3453;
input n_130;
input n_322;
input n_1682;
input n_1980;
input n_2390;
input n_2628;
input n_1249;
input n_3399;
input n_2896;
input n_652;
input n_1111;
input n_3213;
input n_1365;
input n_1927;
input n_25;
input n_3065;
input n_2132;
input n_1349;
input n_1093;
input n_288;
input n_2400;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_3223;
input n_1909;
input n_44;
input n_224;
input n_3077;
input n_2681;
input n_1562;
input n_383;
input n_3103;
input n_834;
input n_3474;
input n_112;
input n_765;
input n_2255;
input n_2424;
input n_2272;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_1965;
input n_239;
input n_3387;
input n_630;
input n_1902;
input n_2151;
input n_1941;
input n_55;
input n_2106;
input n_2775;
input n_2716;
input n_1913;
input n_2878;
input n_504;
input n_1823;
input n_511;
input n_874;
input n_2464;
input n_358;
input n_3422;
input n_1101;
input n_2831;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_3557;
input n_2230;
input n_3498;
input n_2015;
input n_2365;
input n_1875;
input n_1982;
input n_1304;
input n_2803;
input n_1324;
input n_2851;
input n_987;
input n_3189;
input n_1846;
input n_3037;
input n_261;
input n_174;
input n_2066;
input n_1885;
input n_1455;
input n_3429;
input n_767;
input n_993;
input n_1903;
input n_2490;
input n_1407;
input n_2452;
input n_1551;
input n_3154;
input n_545;
input n_441;
input n_860;
input n_3229;
input n_450;
input n_2849;
input n_1805;
input n_2176;
input n_2204;
input n_2905;
input n_1816;
input n_429;
input n_948;
input n_3566;
input n_1217;
input n_2220;
input n_2455;
input n_628;
input n_365;
input n_1849;
input n_2410;
input n_729;
input n_1131;
input n_1084;
input n_1961;
input n_970;
input n_1935;
input n_911;
input n_2922;
input n_1430;
input n_83;
input n_3275;
input n_3499;
input n_2645;
input n_2467;
input n_513;
input n_3366;
input n_2727;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_2288;
input n_3421;
input n_1351;
input n_2240;
input n_2696;
input n_1044;
input n_1205;
input n_2436;
input n_346;
input n_1209;
input n_3029;
input n_1552;
input n_2508;
input n_3242;
input n_3592;
input n_3618;
input n_495;
input n_602;
input n_3525;
input n_574;
input n_2593;
input n_3486;
input n_1435;
input n_879;
input n_3394;
input n_16;
input n_2416;
input n_58;
input n_2405;
input n_623;
input n_3286;
input n_2088;
input n_405;
input n_2953;
input n_824;
input n_359;
input n_1645;
input n_2461;
input n_490;
input n_1327;
input n_2858;
input n_2243;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_2658;
input n_3590;
input n_1717;
input n_572;
input n_366;
input n_2895;
input n_815;
input n_1795;
input n_2128;
input n_2578;
input n_3097;
input n_3483;
input n_128;
input n_1821;
input n_120;
input n_2929;
input n_3424;
input n_327;
input n_3478;
input n_135;
input n_1381;
input n_2555;
input n_2662;
input n_2740;
input n_1611;
input n_1037;
input n_2368;
input n_3388;
input n_2656;
input n_1080;
input n_2301;
input n_1274;
input n_3583;
input n_2890;
input n_3560;
input n_3059;
input n_3524;
input n_2554;
input n_3465;
input n_1316;
input n_1708;
input n_2419;
input n_3215;
input n_426;
input n_1438;
input n_1082;
input n_1840;
input n_589;
input n_716;
input n_1630;
input n_2122;
input n_2512;
input n_3589;
input n_562;
input n_1436;
input n_62;
input n_3549;
input n_1691;
input n_952;
input n_2786;
input n_2534;
input n_2092;
input n_3171;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_2075;
input n_645;
input n_539;
input n_3449;
input n_803;
input n_1092;
input n_2694;
input n_238;
input n_1776;
input n_3559;
input n_2198;
input n_2610;
input n_2661;
input n_2572;
input n_2989;
input n_2281;
input n_2131;
input n_2789;
input n_3026;
input n_2216;
input n_531;
input n_3020;
input n_1757;
input n_890;
input n_1897;
input n_764;
input n_1919;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_3462;
input n_3588;
input n_2933;
input n_2308;
input n_3468;
input n_1893;
input n_2910;
input n_222;
input n_3419;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_2053;
input n_2163;
input n_634;
input n_2328;
input n_199;
input n_1958;
input n_32;
input n_2254;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_3546;
input n_1206;
input n_424;
input n_2647;
input n_3160;
input n_1311;
input n_2191;
input n_2864;
input n_2969;
input n_3195;
input n_1519;
input n_256;
input n_950;
input n_3190;
input n_2428;
input n_1553;
input n_2664;
input n_1811;
input n_2443;
input n_2624;
input n_3012;
input n_3456;
input n_380;
input n_419;
input n_1346;
input n_3053;
input n_444;
input n_1299;
input n_3244;
input n_2158;
input n_1808;
input n_3290;
input n_1060;
input n_1141;
input n_316;
input n_2266;
input n_389;
input n_3130;
input n_2465;
input n_2824;
input n_3033;
input n_2650;
input n_3298;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_3548;
input n_451;
input n_619;
input n_408;
input n_2440;
input n_1386;
input n_1699;
input n_376;
input n_3334;
input n_967;
input n_1442;
input n_2923;
input n_3494;
input n_2541;
input n_74;
input n_1139;
input n_2731;
input n_3264;
input n_515;
input n_2333;
input n_57;
input n_351;
input n_885;
input n_2916;
input n_3166;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_2125;
input n_683;
input n_1632;
input n_3110;
input n_2998;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_2402;
input n_1157;
input n_3073;
input n_2403;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_1954;
input n_2265;
input n_46;
input n_3162;
input n_1608;
input n_983;
input n_1844;
input n_2760;
input n_2792;
input n_3554;
input n_38;
input n_3377;
input n_2870;
input n_280;
input n_1305;
input n_3178;
input n_873;
input n_1826;
input n_378;
input n_1112;
input n_3134;
input n_2304;
input n_2999;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_2334;
input n_2637;
input n_690;
input n_33;
input n_1974;
input n_2463;
input n_583;
input n_2086;
input n_3537;
input n_2289;
input n_3080;
input n_3051;
input n_302;
input n_1343;
input n_2701;
input n_2783;
input n_2263;
input n_3362;
input n_2881;
input n_1203;
input n_1631;
input n_3282;
input n_2472;
input n_821;
input n_1763;
input n_2341;
input n_3105;
input n_3231;
input n_1966;
input n_1768;
input n_321;
input n_2294;
input n_1179;
input n_621;
input n_753;
input n_2475;
input n_2733;
input n_455;
input n_1048;
input n_1719;
input n_2993;
input n_1288;
input n_212;
input n_385;
input n_2785;
input n_2556;
input n_507;
input n_2269;
input n_2732;
input n_3569;
input n_2309;
input n_2415;
input n_2948;
input n_3274;
input n_3041;
input n_3299;
input n_2646;
input n_1560;
input n_1605;
input n_2236;
input n_330;
input n_1228;
input n_2816;
input n_2123;
input n_3209;
input n_972;
input n_3504;
input n_692;
input n_2037;
input n_2685;
input n_3040;
input n_1953;
input n_1938;
input n_820;
input n_1200;
input n_2499;
input n_1911;
input n_3616;
input n_2460;
input n_3568;
input n_2589;
input n_3203;
input n_1301;
input n_1363;
input n_1668;
input n_1185;
input n_991;
input n_2903;
input n_3417;
input n_3482;
input n_828;
input n_1967;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_2233;
input n_1329;
input n_2743;
input n_2675;
input n_3255;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_2827;
input n_1688;
input n_3052;
input n_945;
input n_2997;
input n_492;
input n_3327;
input n_153;
input n_1504;
input n_943;
input n_3326;
input n_341;
input n_3572;
input n_250;
input n_992;
input n_3067;
input n_1932;
input n_3375;
input n_2755;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_3237;
input n_2082;
input n_286;
input n_1992;
input n_2429;
input n_1643;
input n_883;
input n_1983;
input n_3167;
input n_3400;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_3423;
input n_900;
input n_2362;
input n_856;
input n_2609;
input n_1793;
input n_3382;
input n_1976;
input n_2223;
input n_3044;
input n_3574;
input n_918;
input n_3529;
input n_942;
input n_2169;
input n_1804;
input n_189;
input n_1147;
input n_1557;
input n_1977;
input n_2153;
input n_2468;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_3196;
input n_3078;
input n_2364;
input n_2533;
input n_540;
input n_3492;
input n_618;
input n_3094;
input n_896;
input n_2310;
input n_2780;
input n_323;
input n_2287;
input n_2860;
input n_3316;
input n_195;
input n_356;
input n_2291;
input n_3099;
input n_2596;
input n_894;
input n_1636;
input n_2056;
input n_3253;
input n_1730;
input n_3601;
input n_3603;
input n_831;
input n_2280;
input n_2192;
input n_964;
input n_3363;
input n_1373;
input n_1350;
input n_1511;
input n_1865;
input n_2973;
input n_1470;
input n_1096;
input n_2094;
input n_2670;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_2318;
input n_2393;
input n_2020;
input n_5;
input n_1646;
input n_2502;
input n_225;
input n_2504;
input n_1307;
input n_1881;
input n_2974;
input n_988;
input n_2749;
input n_2043;
input n_2901;
input n_1940;
input n_814;
input n_2707;
input n_2751;
input n_2793;
input n_3372;
input n_3451;
input n_192;
input n_2971;
input n_3442;
input n_1549;
input n_1934;
input n_2311;
input n_1201;
input n_1114;
input n_655;
input n_3240;
input n_2025;
input n_1616;
input n_1446;
input n_2285;
input n_3147;
input n_2758;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_2298;
input n_2471;
input n_1807;
input n_387;
input n_1149;
input n_2618;
input n_398;
input n_1671;
input n_635;
input n_2559;
input n_763;
input n_3230;
input n_1020;
input n_1062;
input n_3342;
input n_211;
input n_2303;
input n_1824;
input n_1917;
input n_2295;
input n_1219;
input n_3386;
input n_3;
input n_1204;
input n_2840;
input n_2810;
input n_2325;
input n_178;
input n_2747;
input n_2446;
input n_3488;
input n_1814;
input n_1035;
input n_2822;
input n_287;
input n_555;
input n_783;
input n_1848;
input n_1928;
input n_2126;
input n_2893;
input n_1188;
input n_2588;
input n_2962;
input n_1722;
input n_661;
input n_2441;
input n_41;
input n_1802;
input n_3083;
input n_2600;
input n_849;
input n_2795;
input n_15;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_1786;
input n_2981;
input n_50;
input n_430;
input n_2002;
input n_2282;
input n_3608;
input n_510;
input n_2800;
input n_216;
input n_2371;
input n_2935;
input n_311;
input n_3233;
input n_3380;
input n_3177;
input n_830;
input n_2098;
input n_1296;
input n_2627;
input n_3409;
input n_3460;
input n_2352;
input n_3538;
input n_1413;
input n_801;
input n_2207;
input n_2080;
input n_2377;
input n_2619;
input n_2340;
input n_3085;
input n_2444;
input n_2068;
input n_241;
input n_3552;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_2641;
input n_3198;
input n_749;
input n_1895;
input n_3123;
input n_3137;
input n_2574;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_2361;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_3393;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_2638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_3520;
input n_2492;
input n_1019;
input n_1105;
input n_249;
input n_1998;
input n_304;
input n_1338;
input n_577;
input n_2016;
input n_1522;
input n_2949;
input n_1687;
input n_1637;
input n_2034;
input n_1419;
input n_2711;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_2270;
input n_1506;
input n_3206;
input n_2653;
input n_3578;
input n_14;
input n_836;
input n_990;
input n_2867;
input n_2496;
input n_1886;
input n_1389;
input n_1894;
input n_975;
input n_1908;
input n_1256;
input n_1702;
input n_2259;
input n_2794;
input n_567;
input n_1465;
input n_3145;
input n_3124;
input n_778;
input n_1122;
input n_151;
input n_3192;
input n_2608;
input n_306;
input n_2657;
input n_458;
input n_770;
input n_2995;
input n_1375;
input n_2494;
input n_3547;
input n_2649;
input n_1102;
input n_2852;
input n_2392;
input n_3459;
input n_3093;
input n_1843;
input n_711;
input n_1499;
input n_3061;
input n_3155;
input n_85;
input n_1187;
input n_3517;
input n_2633;
input n_1441;
input n_3100;
input n_2522;
input n_2435;
input n_1392;
input n_1597;
input n_1929;
input n_2807;
input n_1164;
input n_1659;
input n_1834;
input n_2097;
input n_2313;
input n_2542;
input n_489;
input n_1174;
input n_2431;
input n_3324;
input n_3356;
input n_2835;
input n_2558;
input n_1371;
input n_617;
input n_1303;
input n_2206;
input n_2063;
input n_3182;
input n_1572;
input n_1968;
input n_3269;
input n_2564;
input n_2252;
input n_876;
input n_1516;
input n_1190;
input n_3506;
input n_1736;
input n_3605;
input n_1685;
input n_118;
input n_2409;
input n_601;
input n_917;
input n_3450;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_2000;
input n_1661;
input n_3402;
input n_1212;
input n_2074;
input n_1541;
input n_2576;
input n_3565;
input n_172;
input n_206;
input n_217;
input n_726;
input n_3174;
input n_982;
input n_2575;
input n_2988;
input n_3390;
input n_1573;
input n_1453;
input n_1731;
input n_2217;
input n_818;
input n_2373;
input n_1970;
input n_861;
input n_1713;
input n_1183;
input n_3398;
input n_2307;
input n_2766;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_2201;
input n_2722;
input n_2117;
input n_2745;
input n_3408;
input n_1904;
input n_2640;
input n_1993;
input n_774;
input n_1628;
input n_2493;
input n_2205;
input n_3432;
input n_1335;
input n_1514;
input n_1777;
input n_1957;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_1771;
input n_1912;
input n_3401;
input n_1899;
input n_3226;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_3090;
input n_2067;
input n_527;
input n_1168;
input n_707;
input n_2219;
input n_2437;
input n_2885;
input n_3533;
input n_2877;
input n_3318;
input n_2148;
input n_937;
input n_2445;
input n_1427;
input n_2779;
input n_3485;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_1835;
input n_3035;
input n_66;
input n_1440;
input n_177;
input n_2164;
input n_421;
input n_1988;
input n_3333;
input n_2115;
input n_1853;
input n_1356;
input n_2845;
input n_1787;
input n_2634;
input n_910;
input n_2232;
input n_3034;
input n_2212;
input n_2602;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1774;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_2811;
input n_1496;
input n_3348;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_2547;
input n_3014;
input n_708;
input n_529;
input n_1812;
input n_735;
input n_2501;
input n_3079;
input n_232;
input n_1915;
input n_1109;
input n_126;
input n_895;
input n_2532;
input n_1310;
input n_2605;
input n_3358;
input n_2121;
input n_1803;
input n_202;
input n_3308;
input n_2665;
input n_427;
input n_1399;
input n_1543;
input n_1991;
input n_1979;
input n_791;
input n_732;
input n_1533;
input n_2224;
input n_193;
input n_3368;
input n_2924;
input n_3467;
input n_808;
input n_2484;
input n_797;
input n_3530;
input n_1025;
input n_1930;
input n_1955;
input n_2765;
input n_3329;
input n_500;
input n_2994;
input n_1067;
input n_2946;
input n_1720;
input n_148;
input n_2830;
input n_2401;
input n_3135;
input n_435;
input n_2003;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_2692;
input n_3573;
input n_3148;
input n_538;
input n_2354;
input n_2246;
input n_2008;
input n_1117;
input n_799;
input n_2264;
input n_2754;
input n_687;
input n_3534;
input n_715;
input n_1742;
input n_1480;
input n_1482;
input n_1213;
input n_2489;
input n_1266;
input n_536;
input n_3438;
input n_872;
input n_2012;
input n_594;
input n_200;
input n_1291;
input n_3381;
input n_3503;
input n_1297;
input n_1753;
input n_2283;
input n_2866;
input n_3278;
input n_1782;
input n_2245;
input n_3561;
input n_1155;
input n_1418;
input n_89;
input n_1972;
input n_1524;
input n_1689;
input n_1485;
input n_2806;
input n_115;
input n_1011;
input n_1184;
input n_2184;
input n_985;
input n_1855;
input n_2425;
input n_2917;
input n_869;
input n_810;
input n_2965;
input n_3536;
input n_416;
input n_827;
input n_3217;
input n_3404;
input n_3425;
input n_401;
input n_1703;
input n_3312;
input n_1352;
input n_2926;
input n_626;
input n_2197;
input n_2199;
input n_3540;
input n_1650;
input n_1144;
input n_1137;
input n_1570;
input n_2814;
input n_3046;
input n_1170;
input n_305;
input n_2023;
input n_2213;
input n_3249;
input n_3211;
input n_3285;
input n_2351;
input n_2211;
input n_2095;
input n_3121;
input n_137;
input n_676;
input n_294;
input n_318;
input n_2103;
input n_653;
input n_2160;
input n_642;
input n_3337;
input n_2228;
input n_2527;
input n_1602;
input n_2498;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_2697;
input n_850;
input n_684;
input n_3074;
input n_124;
input n_3204;
input n_268;
input n_2421;
input n_2286;
input n_2902;
input n_664;
input n_1999;
input n_503;
input n_2372;
input n_2065;
input n_2136;
input n_2480;
input n_235;
input n_1372;
input n_2861;
input n_605;
input n_2630;
input n_1273;
input n_1822;
input n_3397;
input n_353;
input n_620;
input n_643;
input n_2363;
input n_2430;
input n_916;
input n_1081;
input n_2549;
input n_493;
input n_2705;
input n_3005;
input n_2332;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_2433;
input n_3293;
input n_3129;
input n_1282;
input n_1318;
input n_1783;
input n_780;
input n_2977;
input n_3606;
input n_2601;
input n_3043;
input n_998;
input n_2375;
input n_2550;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_1907;
input n_3600;
input n_501;
input n_823;
input n_245;
input n_2686;
input n_2528;
input n_725;
input n_2344;
input n_1388;
input n_1417;
input n_1295;
input n_2836;
input n_2316;
input n_672;
input n_1985;
input n_3055;
input n_1898;
input n_2107;
input n_3294;
input n_3219;
input n_3315;
input n_581;
input n_2906;
input n_382;
input n_554;
input n_1625;
input n_2130;
input n_3415;
input n_2187;
input n_2284;
input n_898;
input n_2817;
input n_3172;
input n_3139;
input n_2773;
input n_3239;
input n_3292;
input n_2598;
input n_1762;
input n_1013;
input n_3365;
input n_3476;
input n_1452;
input n_718;
input n_2687;
input n_265;
input n_3023;
input n_3553;
input n_1120;
input n_719;
input n_443;
input n_1791;
input n_198;
input n_1890;
input n_1747;
input n_714;
input n_2850;
input n_1683;
input n_1817;
input n_909;
input n_1944;
input n_1497;
input n_1530;
input n_2654;
input n_997;
input n_3431;
input n_3104;
input n_932;
input n_3169;
input n_3151;
input n_612;
input n_3131;
input n_2078;
input n_1409;
input n_788;
input n_1326;
input n_3070;
input n_3284;
input n_119;
input n_3176;
input n_2884;
input n_1268;
input n_2996;
input n_559;
input n_825;
input n_2819;
input n_3126;
input n_1981;
input n_508;
input n_2186;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_3609;
input n_986;
input n_2315;
input n_509;
input n_3228;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_2102;
input n_3581;
input n_2562;
input n_1281;
input n_67;
input n_1952;
input n_1192;
input n_2221;
input n_1024;
input n_3576;
input n_1063;
input n_1889;
input n_209;
input n_1792;
input n_1564;
input n_1868;
input n_1613;
input n_733;
input n_1489;
input n_1922;
input n_2966;
input n_1376;
input n_941;
input n_2326;
input n_981;
input n_2560;
input n_1569;
input n_2188;
input n_68;
input n_3495;
input n_867;
input n_186;
input n_2348;
input n_2422;
input n_134;
input n_2239;
input n_587;
input n_2950;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_2448;
input n_3140;
input n_548;
input n_3170;
input n_812;
input n_298;
input n_2104;
input n_2748;
input n_3311;
input n_518;
input n_505;
input n_2057;
input n_3272;
input n_3011;
input n_1772;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_2898;
input n_782;
input n_2717;
input n_2818;
input n_1100;
input n_1861;
input n_2129;
input n_1395;
input n_3345;
input n_862;
input n_3584;
input n_1425;
input n_760;
input n_1901;
input n_3069;
input n_1900;
input n_1620;
input n_3032;
input n_381;
input n_3628;
input n_2889;
input n_220;
input n_390;
input n_1330;
input n_1867;
input n_31;
input n_1945;
input n_2772;
input n_481;
input n_3018;
input n_1675;
input n_3072;
input n_1924;
input n_2573;
input n_3084;
input n_3081;
input n_3313;
input n_1727;
input n_2710;
input n_1554;
input n_2939;
input n_1745;
input n_2735;
input n_769;
input n_2497;
input n_2006;
input n_3412;
input n_42;
input n_2844;
input n_1995;
input n_2411;
input n_2138;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_2260;
input n_826;
input n_2343;
input n_1813;
input n_2447;
input n_886;
input n_3439;
input n_2014;
input n_3056;
input n_1221;
input n_2345;
input n_2986;
input n_654;
input n_1172;
input n_167;
input n_2535;
input n_379;
input n_428;
input n_1341;
input n_2726;
input n_570;
input n_2774;
input n_3295;
input n_1641;
input n_1361;
input n_3184;
input n_2382;
input n_1707;
input n_853;
input n_3062;
input n_3161;
input n_377;
input n_2317;
input n_751;
input n_3289;
input n_2799;
input n_2172;
input n_1973;
input n_786;
input n_1083;
input n_1142;
input n_2376;
input n_2488;
input n_1129;
input n_392;
input n_2579;
input n_3477;
input n_3017;
input n_158;
input n_3626;
input n_2476;
input n_704;
input n_787;
input n_1770;
input n_138;
input n_2781;
input n_2456;
input n_961;
input n_2250;
input n_2678;
input n_1756;
input n_771;
input n_2778;
input n_276;
input n_95;
input n_1716;
input n_2788;
input n_2872;
input n_1225;
input n_2984;
input n_1520;
input n_2451;
input n_169;
input n_2887;
input n_522;
input n_3364;
input n_1287;
input n_1262;
input n_2691;
input n_400;
input n_930;
input n_181;
input n_1873;
input n_1411;
input n_3201;
input n_3054;
input n_221;
input n_622;
input n_1962;
input n_1577;
input n_2423;
input n_1087;
input n_3472;
input n_2526;
input n_2854;
input n_386;
input n_994;
input n_1701;
input n_3344;
input n_2194;
input n_848;
input n_1550;
input n_2874;
input n_2764;
input n_2703;
input n_1498;
input n_2167;
input n_3302;
input n_3235;
input n_1223;
input n_1272;
input n_2680;
input n_3391;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_2567;
input n_3543;
input n_1247;
input n_2709;
input n_3102;
input n_922;
input n_3122;
input n_816;
input n_1648;
input n_591;
input n_145;
input n_1536;
input n_3050;
input n_3265;
input n_1857;
input n_1344;
input n_2041;
input n_313;
input n_631;
input n_3627;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_1797;
input n_432;
input n_1769;
input n_2957;
input n_839;
input n_3551;
input n_1210;
input n_3518;
input n_2964;
input n_1364;
input n_2956;
input n_2357;
input n_2183;
input n_2673;
input n_2742;
input n_3314;
input n_2360;
input n_3254;
input n_328;
input n_140;
input n_2292;
input n_1250;
input n_2173;
input n_369;
input n_1842;
input n_871;
input n_2442;
input n_3309;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1943;
input n_1460;
input n_772;
input n_2018;
input n_3464;
input n_3260;
input n_1555;
input n_3117;
input n_2834;
input n_3245;
input n_3357;
input n_499;
input n_2531;
input n_1589;
input n_517;
input n_3428;
input n_98;
input n_2961;
input n_402;
input n_413;
input n_1086;
input n_2570;
input n_2702;
input n_796;
input n_1858;
input n_3351;
input n_1619;
input n_3527;
input n_2815;
input n_236;
input n_2119;
input n_1502;
input n_2157;
input n_2552;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_2744;
input n_1348;
input n_2030;
input n_903;
input n_2453;
input n_1525;
input n_1752;
input n_2397;
input n_740;
input n_2883;
input n_3115;
input n_203;
input n_3509;
input n_3352;
input n_384;
input n_2208;
input n_3076;
input n_1404;
input n_80;
input n_3063;
input n_3617;
input n_2912;
input n_1794;
input n_3535;
input n_2182;
input n_35;
input n_1315;
input n_2234;
input n_277;
input n_1061;
input n_3251;
input n_92;
input n_1910;
input n_333;
input n_1298;
input n_2931;
input n_1652;
input n_2209;
input n_462;
input n_2050;
input n_2809;
input n_1193;
input n_2797;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_3118;
input n_29;
input n_79;
input n_3227;
input n_3300;
input n_2321;
input n_3511;
input n_1226;
input n_722;
input n_1277;
input n_2591;
input n_3443;
input n_188;
input n_2146;
input n_844;
input n_201;
input n_3384;
input n_471;
input n_852;
input n_3497;
input n_1487;
input n_40;
input n_1864;
input n_1028;
input n_1601;
input n_3336;
input n_781;
input n_474;
input n_2940;
input n_542;
input n_3435;
input n_3521;
input n_463;
input n_3575;
input n_1546;
input n_595;
input n_502;
input n_3562;
input n_466;
input n_2612;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_2841;
input n_3165;
input n_1627;
input n_2918;
input n_3232;
input n_3322;
input n_1245;
input n_846;
input n_2427;
input n_2438;
input n_2505;
input n_1673;
input n_465;
input n_2832;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_1975;
input n_27;
input n_2296;
input n_2070;
input n_161;
input n_273;
input n_1937;
input n_585;
input n_2112;
input n_3250;
input n_1739;
input n_3181;
input n_270;
input n_2958;
input n_616;
input n_2278;
input n_81;
input n_2594;
input n_3114;
input n_3125;
input n_2394;
input n_3234;
input n_1914;
input n_3612;
input n_2954;
input n_2135;
input n_2335;
input n_2904;
input n_3493;
input n_745;
input n_2381;
input n_3303;
input n_1654;
input n_3004;
input n_3323;
input n_2569;
input n_3112;
input n_2349;
input n_1103;
input n_3132;
input n_3556;
input n_648;
input n_1379;
input n_2734;
input n_312;
input n_2196;
input n_3591;
input n_3024;
input n_2170;
input n_1076;
input n_2823;
input n_1091;
input n_1408;
input n_3512;
input n_494;
input n_1761;
input n_641;
input n_3238;
input n_3210;
input n_730;
input n_3175;
input n_3522;
input n_2036;
input n_1325;
input n_3267;
input n_1595;
input n_2161;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_2404;
input n_2083;
input n_695;
input n_180;
input n_3281;
input n_656;
input n_3307;
input n_1606;
input n_2503;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_3266;
input n_2485;
input n_229;
input n_1936;
input n_1956;
input n_437;
input n_1642;
input n_2279;
input n_3373;
input n_2655;
input n_2027;
input n_60;
input n_403;
input n_453;
input n_2642;
input n_1130;
input n_720;
input n_0;
input n_2500;
input n_2366;
input n_1918;
input n_1526;
input n_863;
input n_2210;
input n_805;
input n_3247;
input n_1604;
input n_1275;
input n_2513;
input n_2525;
input n_3091;
input n_2695;
input n_1764;
input n_3480;
input n_2892;
input n_3057;
input n_3194;
input n_3582;
input n_3066;
input n_113;
input n_712;
input n_2414;
input n_2907;
input n_246;
input n_1583;
input n_2426;
input n_2826;
input n_3577;
input n_3539;
input n_1042;
input n_1402;
input n_2820;
input n_269;
input n_2049;
input n_2273;
input n_285;
input n_412;
input n_2719;
input n_1493;
input n_657;
input n_644;
input n_1741;
input n_2229;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_3347;
input n_2004;
input n_3216;
input n_1621;
input n_2708;
input n_2113;
input n_251;
input n_160;
input n_566;
input n_565;
input n_2586;
input n_1448;
input n_2225;
input n_3567;
input n_3613;
input n_1507;
input n_1398;
input n_2383;
input n_1879;
input n_597;
input n_1996;
input n_3406;
input n_3604;
input n_3444;
input n_1181;
input n_1505;
input n_1634;
input n_1196;
input n_2019;
input n_651;
input n_1340;
input n_2274;
input n_2972;
input n_334;
input n_811;
input n_1558;
input n_3225;
input n_807;
input n_3321;
input n_2166;
input n_2938;
input n_3212;
input n_835;
input n_175;
input n_666;
input n_3319;
input n_262;
input n_1433;
input n_3594;
input n_1704;
input n_2256;
input n_3152;
input n_3335;
input n_99;
input n_1254;
input n_1026;
input n_3413;
input n_2026;
input n_1969;
input n_1234;
input n_2109;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_2013;
input n_1990;
input n_2044;
input n_2689;
input n_2920;
input n_3259;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_2614;
input n_2511;
input n_1681;
input n_2010;
input n_2991;
input n_3383;
input n_1018;
input n_2242;
input n_2247;
input n_2752;
input n_2894;
input n_3016;
input n_1693;
input n_3585;
input n_2975;
input n_3473;
input n_438;
input n_2599;
input n_713;
input n_2704;
input n_904;
input n_2839;
input n_3338;
input n_1588;
input n_1622;
input n_2237;
input n_3414;
input n_3463;
input n_166;
input n_1180;
input n_1827;
input n_3360;
input n_2524;
input n_1271;
input n_2802;
input n_533;
input n_1542;
input n_1251;
input n_3159;
input n_278;
input n_2728;
input n_2268;

output n_15103;

wire n_13115;
wire n_6643;
wire n_6122;
wire n_10564;
wire n_13903;
wire n_7981;
wire n_9936;
wire n_5567;
wire n_4706;
wire n_12148;
wire n_14870;
wire n_9194;
wire n_12407;
wire n_6579;
wire n_9325;
wire n_7164;
wire n_10794;
wire n_5287;
wire n_6546;
wire n_12872;
wire n_13683;
wire n_14881;
wire n_9655;
wire n_14101;
wire n_5484;
wire n_10515;
wire n_11207;
wire n_11326;
wire n_5978;
wire n_8174;
wire n_5161;
wire n_5776;
wire n_14036;
wire n_13241;
wire n_6551;
wire n_13217;
wire n_5512;
wire n_14764;
wire n_10793;
wire n_14635;
wire n_5207;
wire n_12853;
wire n_9044;
wire n_6786;
wire n_12327;
wire n_13927;
wire n_7206;
wire n_7303;
wire n_10552;
wire n_9083;
wire n_12215;
wire n_4963;
wire n_13112;
wire n_14631;
wire n_4240;
wire n_4508;
wire n_8363;
wire n_9408;
wire n_13779;
wire n_12975;
wire n_11802;
wire n_7710;
wire n_8383;
wire n_5035;
wire n_5282;
wire n_10885;
wire n_11583;
wire n_11349;
wire n_8328;
wire n_13499;
wire n_7461;
wire n_12641;
wire n_6649;
wire n_8060;
wire n_9331;
wire n_14203;
wire n_14939;
wire n_7154;
wire n_8551;
wire n_14264;
wire n_13768;
wire n_8002;
wire n_12924;
wire n_4977;
wire n_3813;
wire n_10108;
wire n_8594;
wire n_6810;
wire n_13386;
wire n_7660;
wire n_14070;
wire n_12071;
wire n_6276;
wire n_11016;
wire n_6072;
wire n_12738;
wire n_4128;
wire n_8976;
wire n_4145;
wire n_8617;
wire n_14144;
wire n_5033;
wire n_3785;
wire n_10883;
wire n_7686;
wire n_4211;
wire n_10117;
wire n_12139;
wire n_9846;
wire n_12328;
wire n_8603;
wire n_7024;
wire n_12493;
wire n_14762;
wire n_7205;
wire n_9204;
wire n_6742;
wire n_9769;
wire n_11342;
wire n_9312;
wire n_13493;
wire n_10363;
wire n_8319;
wire n_6694;
wire n_9610;
wire n_3776;
wire n_7616;
wire n_7486;
wire n_4517;
wire n_13220;
wire n_13822;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_11450;
wire n_14287;
wire n_8244;
wire n_12028;
wire n_9273;
wire n_12357;
wire n_4615;
wire n_6090;
wire n_6580;
wire n_12515;
wire n_7010;
wire n_11678;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_14471;
wire n_6913;
wire n_7867;
wire n_13158;
wire n_10756;
wire n_7315;
wire n_11801;
wire n_14435;
wire n_13516;
wire n_11653;
wire n_7004;
wire n_8961;
wire n_13415;
wire n_4131;
wire n_7772;
wire n_10761;
wire n_11299;
wire n_5402;
wire n_13146;
wire n_5851;
wire n_13889;
wire n_5509;
wire n_13775;
wire n_9773;
wire n_8574;
wire n_11089;
wire n_14045;
wire n_11077;
wire n_8864;
wire n_12861;
wire n_9173;
wire n_12709;
wire n_7641;
wire n_11296;
wire n_3796;
wire n_5154;
wire n_9363;
wire n_8681;
wire n_7468;
wire n_9796;
wire n_5469;
wire n_6431;
wire n_11800;
wire n_13906;
wire n_14721;
wire n_12012;
wire n_12462;
wire n_5744;
wire n_14714;
wire n_12266;
wire n_9049;
wire n_11947;
wire n_5453;
wire n_14411;
wire n_11917;
wire n_14537;
wire n_7861;
wire n_9907;
wire n_4499;
wire n_4927;
wire n_8413;
wire n_9738;
wire n_5202;
wire n_5648;
wire n_10745;
wire n_13748;
wire n_14898;
wire n_13178;
wire n_7667;
wire n_13072;
wire n_6931;
wire n_9539;
wire n_14270;
wire n_8114;
wire n_9811;
wire n_12970;
wire n_6618;
wire n_13771;
wire n_6408;
wire n_9993;
wire n_9208;
wire n_14729;
wire n_10421;
wire n_7523;
wire n_4311;
wire n_14800;
wire n_8706;
wire n_3806;
wire n_4691;
wire n_13000;
wire n_5922;
wire n_8158;
wire n_11594;
wire n_12100;
wire n_14959;
wire n_6698;
wire n_4678;
wire n_9500;
wire n_8104;
wire n_10399;
wire n_5848;
wire n_10420;
wire n_12575;
wire n_11635;
wire n_5406;
wire n_12501;
wire n_6085;
wire n_14408;
wire n_3947;
wire n_12819;
wire n_7421;
wire n_7306;
wire n_11505;
wire n_14403;
wire n_8819;
wire n_10535;
wire n_6214;
wire n_7493;
wire n_10360;
wire n_3868;
wire n_9420;
wire n_12027;
wire n_7804;
wire n_8089;
wire n_12111;
wire n_12075;
wire n_12078;
wire n_13401;
wire n_9557;
wire n_4203;
wire n_3687;
wire n_13708;
wire n_9382;
wire n_5241;
wire n_12175;
wire n_6939;
wire n_12604;
wire n_7528;
wire n_11615;
wire n_10307;
wire n_14519;
wire n_10781;
wire n_8262;
wire n_8290;
wire n_9206;
wire n_11507;
wire n_7562;
wire n_12626;
wire n_11497;
wire n_5037;
wire n_9388;
wire n_10193;
wire n_14611;
wire n_11541;
wire n_5661;
wire n_4468;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_8885;
wire n_9772;
wire n_10437;
wire n_12142;
wire n_10430;
wire n_3702;
wire n_8147;
wire n_4976;
wire n_6586;
wire n_11111;
wire n_11354;
wire n_5008;
wire n_10177;
wire n_13782;
wire n_3876;
wire n_8310;
wire n_11052;
wire n_4811;
wire n_5398;
wire n_13875;
wire n_6096;
wire n_6707;
wire n_14170;
wire n_10175;
wire n_5852;
wire n_12767;
wire n_6920;
wire n_13110;
wire n_6868;
wire n_9311;
wire n_12754;
wire n_5144;
wire n_9422;
wire n_14892;
wire n_4758;
wire n_10672;
wire n_9040;
wire n_9795;
wire n_14336;
wire n_8380;
wire n_9027;
wire n_8962;
wire n_12225;
wire n_7402;
wire n_4255;
wire n_5577;
wire n_10626;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_11316;
wire n_7152;
wire n_14579;
wire n_6512;
wire n_9966;
wire n_11272;
wire n_13571;
wire n_13096;
wire n_4237;
wire n_8126;
wire n_5689;
wire n_13087;
wire n_13309;
wire n_10392;
wire n_5894;
wire n_12670;
wire n_12152;
wire n_7801;
wire n_7992;
wire n_11588;
wire n_11689;
wire n_9161;
wire n_10231;
wire n_7463;
wire n_12101;
wire n_8556;
wire n_10316;
wire n_9369;
wire n_13753;
wire n_13147;
wire n_4901;
wire n_9033;
wire n_13542;
wire n_8305;
wire n_10683;
wire n_6725;
wire n_14109;
wire n_7613;
wire n_9429;
wire n_12576;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_14458;
wire n_13610;
wire n_10514;
wire n_6464;
wire n_8317;
wire n_10730;
wire n_10958;
wire n_13095;
wire n_10562;
wire n_11273;
wire n_11962;
wire n_14856;
wire n_15008;
wire n_13706;
wire n_8653;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_14792;
wire n_11303;
wire n_14711;
wire n_7316;
wire n_6820;
wire n_12224;
wire n_5343;
wire n_9780;
wire n_10252;
wire n_4421;
wire n_10438;
wire n_9824;
wire n_6098;
wire n_12237;
wire n_7019;
wire n_12751;
wire n_13612;
wire n_6686;
wire n_11664;
wire n_10523;
wire n_4836;
wire n_11720;
wire n_5062;
wire n_4020;
wire n_10202;
wire n_11398;
wire n_11659;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_8939;
wire n_4532;
wire n_12824;
wire n_9489;
wire n_8604;
wire n_3735;
wire n_7323;
wire n_14405;
wire n_14605;
wire n_11365;
wire n_13755;
wire n_12269;
wire n_7195;
wire n_6701;
wire n_13243;
wire n_10988;
wire n_7478;
wire n_11836;
wire n_6769;
wire n_7683;
wire n_13131;
wire n_6592;
wire n_11150;
wire n_5686;
wire n_12298;
wire n_12019;
wire n_13457;
wire n_5463;
wire n_14263;
wire n_14824;
wire n_5236;
wire n_6062;
wire n_6191;
wire n_7903;
wire n_11003;
wire n_12299;
wire n_9625;
wire n_8440;
wire n_3983;
wire n_10980;
wire n_5433;
wire n_4405;
wire n_10367;
wire n_8525;
wire n_4195;
wire n_8416;
wire n_13734;
wire n_13219;
wire n_4969;
wire n_4504;
wire n_9570;
wire n_12232;
wire n_9368;
wire n_15040;
wire n_8064;
wire n_13547;
wire n_5909;
wire n_7575;
wire n_8879;
wire n_10664;
wire n_4408;
wire n_13458;
wire n_9115;
wire n_9694;
wire n_9367;
wire n_4531;
wire n_6043;
wire n_11520;
wire n_13747;
wire n_12812;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_11099;
wire n_7701;
wire n_4164;
wire n_13223;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_11859;
wire n_13416;
wire n_8931;
wire n_5348;
wire n_8214;
wire n_5055;
wire n_9072;
wire n_14973;
wire n_6793;
wire n_7873;
wire n_9612;
wire n_12777;
wire n_9971;
wire n_13620;
wire n_8729;
wire n_14886;
wire n_7127;
wire n_5397;
wire n_6550;
wire n_4471;
wire n_5031;
wire n_10575;
wire n_11746;
wire n_3975;
wire n_5709;
wire n_4444;
wire n_7568;
wire n_10803;
wire n_6021;
wire n_9720;
wire n_4983;
wire n_5695;
wire n_7814;
wire n_9213;
wire n_10187;
wire n_10400;
wire n_14227;
wire n_14345;
wire n_11330;
wire n_14698;
wire n_10778;
wire n_5860;
wire n_6926;
wire n_4916;
wire n_11121;
wire n_3649;
wire n_9607;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_13283;
wire n_5862;
wire n_6304;
wire n_8228;
wire n_8210;
wire n_5189;
wire n_10586;
wire n_6956;
wire n_10040;
wire n_5381;
wire n_13555;
wire n_4786;
wire n_7026;
wire n_4160;
wire n_6782;
wire n_13582;
wire n_5854;
wire n_11911;
wire n_5516;
wire n_4051;
wire n_9554;
wire n_9262;
wire n_11599;
wire n_12412;
wire n_8387;
wire n_7002;
wire n_12782;
wire n_3981;
wire n_8898;
wire n_8410;
wire n_14852;
wire n_7141;
wire n_14019;
wire n_10935;
wire n_13809;
wire n_5936;
wire n_6126;
wire n_9761;
wire n_12284;
wire n_12612;
wire n_11102;
wire n_8795;
wire n_9649;
wire n_10269;
wire n_10164;
wire n_11039;
wire n_8501;
wire n_12567;
wire n_10401;
wire n_14228;
wire n_6027;
wire n_6598;
wire n_9254;
wire n_9529;
wire n_11535;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_14854;
wire n_14627;
wire n_6638;
wire n_10651;
wire n_7308;
wire n_5254;
wire n_12180;
wire n_6900;
wire n_8953;
wire n_14016;
wire n_13295;
wire n_12731;
wire n_13644;
wire n_9726;
wire n_11686;
wire n_8823;
wire n_12153;
wire n_3790;
wire n_10851;
wire n_7264;
wire n_11730;
wire n_12608;
wire n_7457;
wire n_4613;
wire n_12383;
wire n_7718;
wire n_10918;
wire n_4649;
wire n_7617;
wire n_13629;
wire n_14671;
wire n_15041;
wire n_13360;
wire n_9197;
wire n_14265;
wire n_13351;
wire n_6269;
wire n_8843;
wire n_11942;
wire n_14709;
wire n_5615;
wire n_4795;
wire n_12057;
wire n_14098;
wire n_5902;
wire n_4028;
wire n_7768;
wire n_13083;
wire n_5479;
wire n_10964;
wire n_13294;
wire n_14143;
wire n_13234;
wire n_3819;
wire n_7974;
wire n_13896;
wire n_12902;
wire n_9106;
wire n_6013;
wire n_7357;
wire n_5083;
wire n_8247;
wire n_9564;
wire n_6927;
wire n_9627;
wire n_7975;
wire n_10864;
wire n_13380;
wire n_6503;
wire n_5888;
wire n_8172;
wire n_4186;
wire n_8940;
wire n_8941;
wire n_7310;
wire n_9739;
wire n_10598;
wire n_11835;
wire n_12070;
wire n_13021;
wire n_14797;
wire n_4731;
wire n_11444;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_12430;
wire n_4618;
wire n_7593;
wire n_4742;
wire n_6256;
wire n_7716;
wire n_13971;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_11353;
wire n_10223;
wire n_5870;
wire n_13884;
wire n_9812;
wire n_14905;
wire n_4295;
wire n_14415;
wire n_11823;
wire n_9646;
wire n_5303;
wire n_13686;
wire n_10451;
wire n_10553;
wire n_12718;
wire n_12393;
wire n_10201;
wire n_12249;
wire n_7076;
wire n_11814;
wire n_12719;
wire n_8780;
wire n_10215;
wire n_11205;
wire n_9465;
wire n_12932;
wire n_14093;
wire n_9928;
wire n_14150;
wire n_4694;
wire n_8456;
wire n_9970;
wire n_13719;
wire n_4533;
wire n_11138;
wire n_14238;
wire n_5081;
wire n_9894;
wire n_10100;
wire n_10278;
wire n_5124;
wire n_10436;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_11048;
wire n_4254;
wire n_9129;
wire n_14641;
wire n_6982;
wire n_14616;
wire n_4697;
wire n_14842;
wire n_7286;
wire n_7137;
wire n_12625;
wire n_9957;
wire n_10915;
wire n_13172;
wire n_4190;
wire n_3994;
wire n_9558;
wire n_11292;
wire n_13167;
wire n_11487;
wire n_11753;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_11782;
wire n_8218;
wire n_10689;
wire n_9267;
wire n_12371;
wire n_7539;
wire n_8769;
wire n_7229;
wire n_4391;
wire n_10538;
wire n_8514;
wire n_14628;
wire n_14117;
wire n_13487;
wire n_5954;
wire n_11865;
wire n_12258;
wire n_4157;
wire n_4283;
wire n_8368;
wire n_4681;
wire n_12163;
wire n_8334;
wire n_9918;
wire n_4638;
wire n_8159;
wire n_6097;
wire n_10773;
wire n_11397;
wire n_8639;
wire n_10621;
wire n_5047;
wire n_11600;
wire n_14116;
wire n_12516;
wire n_14342;
wire n_5346;
wire n_14916;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_7797;
wire n_8216;
wire n_4707;
wire n_14979;
wire n_13887;
wire n_4527;
wire n_14740;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_10924;
wire n_11844;
wire n_10874;
wire n_7869;
wire n_6466;
wire n_12871;
wire n_10942;
wire n_12602;
wire n_12295;
wire n_13912;
wire n_14171;
wire n_14830;
wire n_4156;
wire n_9956;
wire n_4848;
wire n_9095;
wire n_9715;
wire n_14975;
wire n_6008;
wire n_15048;
wire n_12198;
wire n_8337;
wire n_11201;
wire n_14141;
wire n_8257;
wire n_11781;
wire n_10292;
wire n_7983;
wire n_11550;
wire n_12077;
wire n_7781;
wire n_8125;
wire n_12166;
wire n_12786;
wire n_13467;
wire n_14677;
wire n_5624;
wire n_14860;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_9246;
wire n_13675;
wire n_7624;
wire n_10653;
wire n_9683;
wire n_12117;
wire n_12110;
wire n_11945;
wire n_14716;
wire n_4898;
wire n_12216;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_8063;
wire n_9931;
wire n_6805;
wire n_12098;
wire n_6185;
wire n_5010;
wire n_7762;
wire n_13097;
wire n_13749;
wire n_15064;
wire n_8731;
wire n_14334;
wire n_14683;
wire n_12102;
wire n_13009;
wire n_14373;
wire n_14325;
wire n_3773;
wire n_8950;
wire n_3918;
wire n_13535;
wire n_14955;
wire n_10624;
wire n_12802;
wire n_13982;
wire n_6568;
wire n_9011;
wire n_9899;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_8295;
wire n_13668;
wire n_12570;
wire n_13577;
wire n_14836;
wire n_4619;
wire n_4673;
wire n_13034;
wire n_6004;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_14292;
wire n_4822;
wire n_8995;
wire n_8146;
wire n_3797;
wire n_11502;
wire n_14583;
wire n_6901;
wire n_8082;
wire n_11965;
wire n_13046;
wire n_11997;
wire n_9094;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_14589;
wire n_4801;
wire n_7183;
wire n_13300;
wire n_12456;
wire n_11424;
wire n_6411;
wire n_8339;
wire n_13405;
wire n_11816;
wire n_9195;
wire n_7746;
wire n_13641;
wire n_5435;
wire n_12768;
wire n_10867;
wire n_11361;
wire n_10701;
wire n_14735;
wire n_14233;
wire n_11062;
wire n_14068;
wire n_6873;
wire n_14610;
wire n_4279;
wire n_4769;
wire n_14584;
wire n_4632;
wire n_10741;
wire n_5373;
wire n_5745;
wire n_8032;
wire n_14505;
wire n_7139;
wire n_14655;
wire n_12710;
wire n_12483;
wire n_8640;
wire n_4294;
wire n_9332;
wire n_10016;
wire n_10070;
wire n_5279;
wire n_14121;
wire n_4125;
wire n_4232;
wire n_8351;
wire n_4949;
wire n_10190;
wire n_14673;
wire n_11499;
wire n_8196;
wire n_11580;
wire n_15084;
wire n_12128;
wire n_6594;
wire n_5493;
wire n_4790;
wire n_7857;
wire n_9054;
wire n_10812;
wire n_10150;
wire n_9460;
wire n_9638;
wire n_12682;
wire n_13028;
wire n_6387;
wire n_14896;
wire n_13613;
wire n_12389;
wire n_7223;
wire n_7890;
wire n_12464;
wire n_4847;
wire n_6179;
wire n_9281;
wire n_7338;
wire n_5321;
wire n_10134;
wire n_11379;
wire n_13700;
wire n_7964;
wire n_13135;
wire n_5096;
wire n_9740;
wire n_4365;
wire n_9475;
wire n_8865;
wire n_9661;
wire n_13721;
wire n_13056;
wire n_10861;
wire n_6019;
wire n_12313;
wire n_12147;
wire n_11070;
wire n_9190;
wire n_6222;
wire n_7165;
wire n_8110;
wire n_11245;
wire n_10635;
wire n_12874;
wire n_14749;
wire n_6223;
wire n_8475;
wire n_8838;
wire n_4610;
wire n_6435;
wire n_12909;
wire n_9143;
wire n_4489;
wire n_3730;
wire n_12990;
wire n_14871;
wire n_7235;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_8488;
wire n_11286;
wire n_5657;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_8766;
wire n_6844;
wire n_13628;
wire n_7795;
wire n_8969;
wire n_12240;
wire n_11631;
wire n_7404;
wire n_3945;
wire n_13326;
wire n_9891;
wire n_10555;
wire n_4542;
wire n_6295;
wire n_10897;
wire n_11147;
wire n_9087;
wire n_11700;
wire n_9804;
wire n_10287;
wire n_8087;
wire n_8119;
wire n_10135;
wire n_9321;
wire n_7885;
wire n_12468;
wire n_4198;
wire n_5857;
wire n_10983;
wire n_8173;
wire n_4534;
wire n_4500;
wire n_11833;
wire n_9800;
wire n_7437;
wire n_5014;
wire n_11053;
wire n_6241;
wire n_8420;
wire n_6087;
wire n_14035;
wire n_8019;
wire n_9186;
wire n_13307;
wire n_9951;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_4087;
wire n_9243;
wire n_11335;
wire n_14346;
wire n_14921;
wire n_3811;
wire n_13509;
wire n_14902;
wire n_5756;
wire n_12294;
wire n_11336;
wire n_11057;
wire n_11247;
wire n_6041;
wire n_7822;
wire n_12186;
wire n_8851;
wire n_14949;
wire n_6994;
wire n_15069;
wire n_10987;
wire n_4257;
wire n_7449;
wire n_11262;
wire n_7329;
wire n_9359;
wire n_5708;
wire n_10402;
wire n_15083;
wire n_13238;
wire n_8687;
wire n_6790;
wire n_14813;
wire n_12860;
wire n_10001;
wire n_13598;
wire n_10666;
wire n_7194;
wire n_11363;
wire n_6273;
wire n_14482;
wire n_11783;
wire n_8740;
wire n_11661;
wire n_14450;
wire n_11026;
wire n_3984;
wire n_6807;
wire n_11889;
wire n_15066;
wire n_14806;
wire n_14990;
wire n_5927;
wire n_10189;
wire n_12939;
wire n_9879;
wire n_4665;
wire n_8221;
wire n_8468;
wire n_7708;
wire n_7696;
wire n_14708;
wire n_11756;
wire n_3679;
wire n_13153;
wire n_11419;
wire n_11232;
wire n_13211;
wire n_3888;
wire n_5638;
wire n_9975;
wire n_10997;
wire n_7115;
wire n_9335;
wire n_13763;
wire n_4189;
wire n_5670;
wire n_9171;
wire n_12778;
wire n_8815;
wire n_14994;
wire n_9942;
wire n_11081;
wire n_13304;
wire n_3707;
wire n_12813;
wire n_13391;
wire n_13711;
wire n_11407;
wire n_5584;
wire n_8952;
wire n_14102;
wire n_11654;
wire n_3849;
wire n_3946;
wire n_9247;
wire n_9933;
wire n_5965;
wire n_12907;
wire n_4463;
wire n_7958;
wire n_10209;
wire n_8128;
wire n_11519;
wire n_4687;
wire n_5751;
wire n_13475;
wire n_10434;
wire n_5664;
wire n_12011;
wire n_9441;
wire n_11668;
wire n_11913;
wire n_4670;
wire n_11978;
wire n_15013;
wire n_4084;
wire n_4703;
wire n_15014;
wire n_10829;
wire n_5641;
wire n_8667;
wire n_4037;
wire n_6218;
wire n_8863;
wire n_7281;
wire n_10233;
wire n_11810;
wire n_8106;
wire n_9362;
wire n_10690;
wire n_14212;
wire n_10311;
wire n_14001;
wire n_6824;
wire n_11198;
wire n_11767;
wire n_8717;
wire n_14712;
wire n_6189;
wire n_11595;
wire n_13305;
wire n_9216;
wire n_11168;
wire n_8299;
wire n_5262;
wire n_9200;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_11872;
wire n_13787;
wire n_5963;
wire n_3808;
wire n_5980;
wire n_8892;
wire n_11235;
wire n_12007;
wire n_10146;
wire n_4763;
wire n_14445;
wire n_14550;
wire n_9067;
wire n_12712;
wire n_5310;
wire n_9152;
wire n_12846;
wire n_8287;
wire n_11906;
wire n_13837;
wire n_14604;
wire n_4594;
wire n_6153;
wire n_9074;
wire n_13550;
wire n_7989;
wire n_14528;
wire n_13908;
wire n_15019;
wire n_10790;
wire n_5970;
wire n_6418;
wire n_12908;
wire n_6564;
wire n_13461;
wire n_13955;
wire n_8657;
wire n_12505;
wire n_12747;
wire n_12577;
wire n_4076;
wire n_4714;
wire n_12426;
wire n_5146;
wire n_4776;
wire n_11122;
wire n_9287;
wire n_4102;
wire n_8197;
wire n_9511;
wire n_14500;
wire n_13733;
wire n_10052;
wire n_13067;
wire n_8081;
wire n_7192;
wire n_12309;
wire n_13974;
wire n_6671;
wire n_10407;
wire n_10449;
wire n_11324;
wire n_12164;
wire n_6591;
wire n_6266;
wire n_10950;
wire n_14235;
wire n_14425;
wire n_7161;
wire n_11566;
wire n_14352;
wire n_7580;
wire n_7153;
wire n_9880;
wire n_10072;
wire n_14929;
wire n_9843;
wire n_5213;
wire n_8609;
wire n_3677;
wire n_11869;
wire n_14609;
wire n_5441;
wire n_6517;
wire n_14326;
wire n_11579;
wire n_14196;
wire n_8559;
wire n_7350;
wire n_10838;
wire n_5690;
wire n_12140;
wire n_13312;
wire n_10369;
wire n_14075;
wire n_6967;
wire n_5885;
wire n_10920;
wire n_9248;
wire n_6433;
wire n_10321;
wire n_12178;
wire n_7535;
wire n_6893;
wire n_9128;
wire n_13003;
wire n_8452;
wire n_14261;
wire n_10506;
wire n_4443;
wire n_5461;
wire n_11082;
wire n_4507;
wire n_7178;
wire n_13192;
wire n_7480;
wire n_10224;
wire n_7632;
wire n_4575;
wire n_12554;
wire n_10671;
wire n_8771;
wire n_8140;
wire n_8476;
wire n_9528;
wire n_12912;
wire n_13213;
wire n_6501;
wire n_8981;
wire n_10157;
wire n_12200;
wire n_11529;
wire n_9507;
wire n_6028;
wire n_14603;
wire n_3822;
wire n_13557;
wire n_14332;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_9533;
wire n_13890;
wire n_12611;
wire n_13767;
wire n_5362;
wire n_8137;
wire n_6709;
wire n_14285;
wire n_4355;
wire n_14443;
wire n_12322;
wire n_8469;
wire n_13270;
wire n_10808;
wire n_6798;
wire n_12303;
wire n_12507;
wire n_5702;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_7844;
wire n_3771;
wire n_5199;
wire n_11430;
wire n_11882;
wire n_12023;
wire n_14379;
wire n_13802;
wire n_14991;
wire n_9665;
wire n_4572;
wire n_12171;
wire n_8423;
wire n_13476;
wire n_12395;
wire n_12472;
wire n_12815;
wire n_5527;
wire n_6986;
wire n_11146;
wire n_8090;
wire n_5609;
wire n_12239;
wire n_5416;
wire n_10504;
wire n_4026;
wire n_11279;
wire n_4104;
wire n_10975;
wire n_4512;
wire n_13176;
wire n_4377;
wire n_5266;
wire n_7471;
wire n_13443;
wire n_13418;
wire n_9436;
wire n_5355;
wire n_9562;
wire n_6745;
wire n_11516;
wire n_11005;
wire n_8260;
wire n_4521;
wire n_8481;
wire n_13961;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_14811;
wire n_6209;
wire n_6875;
wire n_13799;
wire n_10566;
wire n_3750;
wire n_3632;
wire n_14685;
wire n_11451;
wire n_4588;
wire n_14146;
wire n_11980;
wire n_11076;
wire n_7905;
wire n_14877;
wire n_6853;
wire n_4519;
wire n_12121;
wire n_15020;
wire n_5551;
wire n_7594;
wire n_7766;
wire n_3715;
wire n_7803;
wire n_7340;
wire n_10837;
wire n_6699;
wire n_7747;
wire n_6073;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_12116;
wire n_8651;
wire n_14260;
wire n_5640;
wire n_10199;
wire n_13020;
wire n_13621;
wire n_8284;
wire n_10688;
wire n_14999;
wire n_12261;
wire n_9255;
wire n_10039;
wire n_8828;
wire n_5655;
wire n_5475;
wire n_11239;
wire n_12338;
wire n_12259;
wire n_14310;
wire n_3737;
wire n_14608;
wire n_7603;
wire n_6138;
wire n_8510;
wire n_8810;
wire n_13163;
wire n_9034;
wire n_9203;
wire n_9601;
wire n_13173;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_10443;
wire n_11623;
wire n_12825;
wire n_7494;
wire n_5921;
wire n_12222;
wire n_8024;
wire n_9946;
wire n_14383;
wire n_4400;
wire n_5168;
wire n_10887;
wire n_13253;
wire n_13119;
wire n_9967;
wire n_6477;
wire n_10735;
wire n_10274;
wire n_8739;
wire n_3734;
wire n_8373;
wire n_8133;
wire n_8919;
wire n_11740;
wire n_14469;
wire n_4778;
wire n_13525;
wire n_10482;
wire n_6159;
wire n_11012;
wire n_9647;
wire n_6283;
wire n_7396;
wire n_9912;
wire n_14237;
wire n_5322;
wire n_14774;
wire n_11698;
wire n_7116;
wire n_12779;
wire n_14782;
wire n_14694;
wire n_7519;
wire n_4352;
wire n_10485;
wire n_4441;
wire n_6943;
wire n_9329;
wire n_6827;
wire n_4761;
wire n_10652;
wire n_12465;
wire n_6173;
wire n_8318;
wire n_13042;
wire n_8542;
wire n_11059;
wire n_14592;
wire n_4347;
wire n_4095;
wire n_8543;
wire n_8846;
wire n_10791;
wire n_4593;
wire n_6312;
wire n_14803;
wire n_14895;
wire n_11236;
wire n_13514;
wire n_14183;
wire n_4727;
wire n_4568;
wire n_12852;
wire n_13994;
wire n_5371;
wire n_12334;
wire n_4043;
wire n_13162;
wire n_6997;
wire n_15044;
wire n_5418;
wire n_15095;
wire n_11196;
wire n_11629;
wire n_10411;
wire n_12847;
wire n_7770;
wire n_10286;
wire n_14679;
wire n_12511;
wire n_11643;
wire n_7664;
wire n_10913;
wire n_13199;
wire n_15068;
wire n_5316;
wire n_9890;
wire n_13969;
wire n_3831;
wire n_14736;
wire n_10273;
wire n_15005;
wire n_3801;
wire n_6300;
wire n_9609;
wire n_9883;
wire n_10172;
wire n_7815;
wire n_13209;
wire n_12014;
wire n_9046;
wire n_13407;
wire n_9361;
wire n_8163;
wire n_13980;
wire n_11609;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_10806;
wire n_6537;
wire n_13712;
wire n_5933;
wire n_13059;
wire n_12305;
wire n_4948;
wire n_4000;
wire n_13681;
wire n_14864;
wire n_9864;
wire n_13521;
wire n_4406;
wire n_12485;
wire n_7023;
wire n_8972;
wire n_9300;
wire n_12408;
wire n_13263;
wire n_12238;
wire n_7428;
wire n_5112;
wire n_10694;
wire n_5386;
wire n_11509;
wire n_6783;
wire n_11351;
wire n_9353;
wire n_4748;
wire n_9766;
wire n_7465;
wire n_13720;
wire n_3931;
wire n_4010;
wire n_11271;
wire n_8293;
wire n_5017;
wire n_9832;
wire n_14421;
wire n_10754;
wire n_14480;
wire n_4710;
wire n_14663;
wire n_12409;
wire n_13565;
wire n_11307;
wire n_13685;
wire n_5123;
wire n_4607;
wire n_9954;
wire n_4117;
wire n_8737;
wire n_3636;
wire n_13129;
wire n_14091;
wire n_7961;
wire n_10953;
wire n_11761;
wire n_7847;
wire n_9997;
wire n_10703;
wire n_14427;
wire n_11973;
wire n_4487;
wire n_5001;
wire n_9334;
wire n_7149;
wire n_8252;
wire n_15052;
wire n_6459;
wire n_9622;
wire n_10847;
wire n_11565;
wire n_14088;
wire n_13446;
wire n_11252;
wire n_8450;
wire n_4817;
wire n_7700;
wire n_9284;
wire n_5644;
wire n_14318;
wire n_13865;
wire n_9147;
wire n_8367;
wire n_12454;
wire n_10103;
wire n_8834;
wire n_6869;
wire n_8078;
wire n_10922;
wire n_10413;
wire n_11571;
wire n_4849;
wire n_10738;
wire n_12587;
wire n_4867;
wire n_13197;
wire n_5424;
wire n_7914;
wire n_13916;
wire n_10995;
wire n_7967;
wire n_9794;
wire n_11858;
wire n_4728;
wire n_14812;
wire n_13963;
wire n_7117;
wire n_14845;
wire n_9354;
wire n_8471;
wire n_11904;
wire n_12324;
wire n_13925;
wire n_4247;
wire n_4933;
wire n_12130;
wire n_6977;
wire n_4018;
wire n_8474;
wire n_12643;
wire n_3900;
wire n_7984;
wire n_13448;
wire n_10185;
wire n_11131;
wire n_4902;
wire n_11478;
wire n_4518;
wire n_10591;
wire n_11656;
wire n_14426;
wire n_12955;
wire n_4409;
wire n_4411;
wire n_11673;
wire n_11821;
wire n_8361;
wire n_6313;
wire n_3872;
wire n_11701;
wire n_10856;
wire n_14348;
wire n_13626;
wire n_4336;
wire n_6569;
wire n_4777;
wire n_9494;
wire n_6555;
wire n_9614;
wire n_11283;
wire n_13616;
wire n_12948;
wire n_14329;
wire n_9551;
wire n_3877;
wire n_13653;
wire n_6639;
wire n_7516;
wire n_5496;
wire n_13694;
wire n_3977;
wire n_9154;
wire n_13233;
wire n_10677;
wire n_7596;
wire n_13189;
wire n_4052;
wire n_13640;
wire n_5864;
wire n_6536;
wire n_14211;
wire n_4398;
wire n_8553;
wire n_6490;
wire n_8301;
wire n_15003;
wire n_10610;
wire n_6961;
wire n_13392;
wire n_4954;
wire n_12574;
wire n_12697;
wire n_9437;
wire n_5460;
wire n_7628;
wire n_9276;
wire n_4304;
wire n_6761;
wire n_14572;
wire n_9346;
wire n_11229;
wire n_3911;
wire n_5333;
wire n_6294;
wire n_14851;
wire n_11636;
wire n_6767;
wire n_8518;
wire n_7427;
wire n_4431;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_13962;
wire n_12162;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_9514;
wire n_4805;
wire n_11919;
wire n_9402;
wire n_14118;
wire n_10456;
wire n_12634;
wire n_11675;
wire n_10343;
wire n_4885;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_9580;
wire n_14134;
wire n_9005;
wire n_5804;
wire n_12236;
wire n_7979;
wire n_6376;
wire n_8621;
wire n_6167;
wire n_8993;
wire n_7926;
wire n_4701;
wire n_12632;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_12398;
wire n_14545;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_10979;
wire n_13591;
wire n_10487;
wire n_10332;
wire n_9162;
wire n_9921;
wire n_9443;
wire n_6582;
wire n_13479;
wire n_8910;
wire n_7752;
wire n_13631;
wire n_9897;
wire n_11570;
wire n_10807;
wire n_6996;
wire n_11855;
wire n_9817;
wire n_14930;
wire n_11667;
wire n_9301;
wire n_6974;
wire n_7731;
wire n_8753;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_9401;
wire n_8321;
wire n_6921;
wire n_11290;
wire n_13738;
wire n_8044;
wire n_8091;
wire n_14137;
wire n_8486;
wire n_7845;
wire n_13122;
wire n_10750;
wire n_12292;
wire n_7709;
wire n_9689;
wire n_4631;
wire n_11592;
wire n_11466;
wire n_5194;
wire n_13346;
wire n_9982;
wire n_6898;
wire n_12056;
wire n_6710;
wire n_13149;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_8508;
wire n_12679;
wire n_8261;
wire n_14179;
wire n_12811;
wire n_13100;
wire n_14821;
wire n_5886;
wire n_7080;
wire n_9886;
wire n_7744;
wire n_13232;
wire n_12897;
wire n_8034;
wire n_8841;
wire n_10970;
wire n_14401;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_12837;
wire n_4965;
wire n_10264;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_5610;
wire n_6836;
wire n_5239;
wire n_11983;
wire n_13840;
wire n_12605;
wire n_11043;
wire n_4747;
wire n_5197;
wire n_8947;
wire n_9671;
wire n_6972;
wire n_9297;
wire n_10472;
wire n_8788;
wire n_13460;
wire n_13389;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_14180;
wire n_5785;
wire n_4587;
wire n_3731;
wire n_11415;
wire n_13578;
wire n_6344;
wire n_14773;
wire n_5305;
wire n_5994;
wire n_6093;
wire n_4538;
wire n_10499;
wire n_8093;
wire n_11680;
wire n_13870;
wire n_15096;
wire n_6010;
wire n_14958;
wire n_7247;
wire n_13088;
wire n_11446;
wire n_9225;
wire n_8061;
wire n_6833;
wire n_11972;
wire n_14247;
wire n_5376;
wire n_13862;
wire n_13600;
wire n_11103;
wire n_7481;
wire n_10435;
wire n_12220;
wire n_13843;
wire n_10066;
wire n_13605;
wire n_14707;
wire n_5204;
wire n_7292;
wire n_10341;
wire n_12230;
wire n_14511;
wire n_4094;
wire n_8811;
wire n_12995;
wire n_7150;
wire n_13486;
wire n_14176;
wire n_7687;
wire n_10184;
wire n_10498;
wire n_13599;
wire n_12867;
wire n_9662;
wire n_8507;
wire n_10508;
wire n_9057;
wire n_3661;
wire n_12497;
wire n_14173;
wire n_14323;
wire n_4150;
wire n_14667;
wire n_4878;
wire n_12406;
wire n_6265;
wire n_8861;
wire n_14544;
wire n_11749;
wire n_14875;
wire n_6821;
wire n_8661;
wire n_11417;
wire n_3934;
wire n_8545;
wire n_12725;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_8755;
wire n_5788;
wire n_11490;
wire n_12401;
wire n_13404;
wire n_8573;
wire n_8191;
wire n_11704;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_10865;
wire n_11343;
wire n_14777;
wire n_15065;
wire n_9809;
wire n_13277;
wire n_12185;
wire n_13518;
wire n_14157;
wire n_8683;
wire n_10081;
wire n_8836;
wire n_6676;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_13540;
wire n_12161;
wire n_14366;
wire n_3768;
wire n_9448;
wire n_3943;
wire n_8136;
wire n_8446;
wire n_9799;
wire n_7742;
wire n_10577;
wire n_9313;
wire n_15085;
wire n_8916;
wire n_14650;
wire n_14657;
wire n_7955;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_10037;
wire n_13370;
wire n_12424;
wire n_5582;
wire n_10234;
wire n_14801;
wire n_7374;
wire n_4022;
wire n_7440;
wire n_9989;
wire n_11766;
wire n_4852;
wire n_7758;
wire n_11639;
wire n_7547;
wire n_14802;
wire n_12114;
wire n_13171;
wire n_11967;
wire n_4869;
wire n_9438;
wire n_13528;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_13419;
wire n_14087;
wire n_11457;
wire n_4426;
wire n_10832;
wire n_12490;
wire n_10036;
wire n_12571;
wire n_11932;
wire n_15053;
wire n_5746;
wire n_5292;
wire n_14656;
wire n_10853;
wire n_12508;
wire n_12582;
wire n_6648;
wire n_7880;
wire n_12052;
wire n_14757;
wire n_4601;
wire n_8075;
wire n_13937;
wire n_14298;
wire n_14623;
wire n_8857;
wire n_11275;
wire n_14253;
wire n_4220;
wire n_8587;
wire n_12337;
wire n_9675;
wire n_10030;
wire n_5630;
wire n_9667;
wire n_10676;
wire n_11819;
wire n_8071;
wire n_13159;
wire n_10815;
wire n_12928;
wire n_11589;
wire n_11309;
wire n_12927;
wire n_4066;
wire n_13347;
wire n_11803;
wire n_7513;
wire n_11067;
wire n_12321;
wire n_4515;
wire n_4351;
wire n_11274;
wire n_5264;
wire n_9537;
wire n_10833;
wire n_7413;
wire n_11174;
wire n_4403;
wire n_11795;
wire n_11770;
wire n_7540;
wire n_8646;
wire n_4858;
wire n_4509;
wire n_3700;
wire n_9866;
wire n_5504;
wire n_8630;
wire n_7622;
wire n_9602;
wire n_14392;
wire n_7005;
wire n_11266;
wire n_11151;
wire n_4223;
wire n_7353;
wire n_6219;
wire n_10071;
wire n_9885;
wire n_14115;
wire n_12592;
wire n_14992;
wire n_12698;
wire n_13343;
wire n_8315;
wire n_14282;
wire n_6965;
wire n_9260;
wire n_13938;
wire n_5025;
wire n_8314;
wire n_12048;
wire n_6720;
wire n_14615;
wire n_8149;
wire n_6032;
wire n_11413;
wire n_8581;
wire n_13932;
wire n_13094;
wire n_7174;
wire n_8565;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_14668;
wire n_14509;
wire n_4644;
wire n_7166;
wire n_5060;
wire n_4456;
wire n_7607;
wire n_8209;
wire n_9159;
wire n_5334;
wire n_4346;
wire n_7816;
wire n_13290;
wire n_9654;
wire n_8560;
wire n_7591;
wire n_5775;
wire n_8141;
wire n_14139;
wire n_7830;
wire n_7282;
wire n_6491;
wire n_13198;
wire n_8302;
wire n_10015;
wire n_9306;
wire n_11682;
wire n_7151;
wire n_11652;
wire n_12801;
wire n_6229;
wire n_11091;
wire n_11929;
wire n_9978;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_10362;
wire n_4235;
wire n_7053;
wire n_8724;
wire n_11331;
wire n_11640;
wire n_14702;
wire n_5831;
wire n_10171;
wire n_12552;
wire n_7473;
wire n_4435;
wire n_10183;
wire n_10471;
wire n_14674;
wire n_8070;
wire n_6835;
wire n_13039;
wire n_6419;
wire n_6039;
wire n_12704;
wire n_11237;
wire n_3807;
wire n_11601;
wire n_11741;
wire n_14130;
wire n_14402;
wire n_14305;
wire n_5884;
wire n_14400;
wire n_9279;
wire n_8457;
wire n_4764;
wire n_5653;
wire n_8922;
wire n_8248;
wire n_7966;
wire n_9509;
wire n_6258;
wire n_10095;
wire n_10549;
wire n_7070;
wire n_5394;
wire n_11721;
wire n_6755;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_12256;
wire n_7942;
wire n_10057;
wire n_4655;
wire n_12477;
wire n_4581;
wire n_12184;
wire n_11093;
wire n_12245;
wire n_6084;
wire n_10301;
wire n_4827;
wire n_9496;
wire n_13156;
wire n_8411;
wire n_12740;
wire n_12657;
wire n_9644;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_7666;
wire n_12089;
wire n_14051;
wire n_6472;
wire n_13957;
wire n_5421;
wire n_8527;
wire n_7211;
wire n_10394;
wire n_10154;
wire n_4399;
wire n_11097;
wire n_11681;
wire n_6531;
wire n_5309;
wire n_7901;
wire n_8689;
wire n_11522;
wire n_14724;
wire n_9750;
wire n_4782;
wire n_9980;
wire n_13164;
wire n_10818;
wire n_12145;
wire n_8988;
wire n_11105;
wire n_4363;
wire n_12647;
wire n_12377;
wire n_12721;
wire n_4864;
wire n_9251;
wire n_10141;
wire n_7368;
wire n_13624;
wire n_8549;
wire n_12541;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_12316;
wire n_11849;
wire n_6771;
wire n_11578;
wire n_13484;
wire n_10916;
wire n_10208;
wire n_6389;
wire n_13714;
wire n_10182;
wire n_13655;
wire n_9616;
wire n_15037;
wire n_12399;
wire n_8004;
wire n_10929;
wire n_8658;
wire n_9959;
wire n_8375;
wire n_10403;
wire n_5764;
wire n_10260;
wire n_6910;
wire n_5428;
wire n_9291;
wire n_9092;
wire n_10261;
wire n_6442;
wire n_12285;
wire n_13606;
wire n_6102;
wire n_8908;
wire n_5541;
wire n_4259;
wire n_15067;
wire n_13438;
wire n_10384;
wire n_6441;
wire n_5543;
wire n_10372;
wire n_9818;
wire n_10237;
wire n_9283;
wire n_5935;
wire n_5678;
wire n_4865;
wire n_11219;
wire n_4056;
wire n_13498;
wire n_14453;
wire n_4564;
wire n_3840;
wire n_7677;
wire n_5085;
wire n_8569;
wire n_3733;
wire n_13661;
wire n_8676;
wire n_10118;
wire n_5950;
wire n_12379;
wire n_13496;
wire n_7929;
wire n_10028;
wire n_12257;
wire n_3738;
wire n_10691;
wire n_8399;
wire n_5995;
wire n_12246;
wire n_11069;
wire n_6162;
wire n_5116;
wire n_4526;
wire n_6331;
wire n_13674;
wire n_6006;
wire n_14099;
wire n_8421;
wire n_6109;
wire n_4417;
wire n_11268;
wire n_6278;
wire n_9304;
wire n_12655;
wire n_13818;
wire n_14855;
wire n_6787;
wire n_10777;
wire n_11066;
wire n_6872;
wire n_4899;
wire n_6208;
wire n_14642;
wire n_6632;
wire n_13133;
wire n_9310;
wire n_5411;
wire n_7754;
wire n_14246;
wire n_4798;
wire n_9830;
wire n_9913;
wire n_11728;
wire n_7027;
wire n_8001;
wire n_5671;
wire n_8322;
wire n_12272;
wire n_6990;
wire n_12862;
wire n_8403;
wire n_6349;
wire n_14885;
wire n_13140;
wire n_11796;
wire n_13573;
wire n_7631;
wire n_6830;
wire n_8999;
wire n_12662;
wire n_8754;
wire n_5185;
wire n_7939;
wire n_8675;
wire n_7898;
wire n_10715;
wire n_12136;
wire n_14889;
wire n_6359;
wire n_9375;
wire n_8596;
wire n_10665;
wire n_10073;
wire n_10291;
wire n_13251;
wire n_14890;
wire n_8858;
wire n_8666;
wire n_11873;
wire n_8313;
wire n_7763;
wire n_10296;
wire n_13154;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3935;
wire n_7377;
wire n_11228;
wire n_8555;
wire n_5379;
wire n_3948;
wire n_4750;
wire n_12517;
wire n_13796;
wire n_6301;
wire n_12031;
wire n_11743;
wire n_14274;
wire n_10512;
wire n_8610;
wire n_13195;
wire n_13314;
wire n_14456;
wire n_13679;
wire n_12993;
wire n_10324;
wire n_13658;
wire n_12663;
wire n_7945;
wire n_5945;
wire n_14850;
wire n_11261;
wire n_13667;
wire n_9323;
wire n_6744;
wire n_4981;
wire n_10765;
wire n_9985;
wire n_12039;
wire n_11023;
wire n_8615;
wire n_11382;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_14278;
wire n_10026;
wire n_8677;
wire n_9355;
wire n_8602;
wire n_9714;
wire n_12938;
wire n_7381;
wire n_13772;
wire n_10041;
wire n_5565;
wire n_4081;
wire n_7948;
wire n_4407;
wire n_8102;
wire n_7291;
wire n_9540;
wire n_14840;
wire n_3951;
wire n_4894;
wire n_13033;
wire n_9753;
wire n_5780;
wire n_8460;
wire n_9105;
wire n_13746;
wire n_5643;
wire n_11305;
wire n_10149;
wire n_12680;
wire n_13017;
wire n_14530;
wire n_11137;
wire n_11607;
wire n_5846;
wire n_7430;
wire n_9700;
wire n_14234;
wire n_12930;
wire n_13914;
wire n_13752;
wire n_4995;
wire n_15093;
wire n_8871;
wire n_10649;
wire n_14360;
wire n_9476;
wire n_12722;
wire n_7870;
wire n_13529;
wire n_9875;
wire n_11265;
wire n_10593;
wire n_12042;
wire n_5524;
wire n_8824;
wire n_14827;
wire n_3964;
wire n_3772;
wire n_10597;
wire n_9963;
wire n_6104;
wire n_4446;
wire n_12469;
wire n_6475;
wire n_3884;
wire n_8470;
wire n_9582;
wire n_12172;
wire n_11739;
wire n_10817;
wire n_6465;
wire n_10060;
wire n_9574;
wire n_12049;
wire n_3726;
wire n_6496;
wire n_13229;
wire n_13973;
wire n_11687;
wire n_14160;
wire n_9732;
wire n_11050;
wire n_13070;
wire n_14440;
wire n_12666;
wire n_8238;
wire n_9882;
wire n_12205;
wire n_6998;
wire n_10779;
wire n_13177;
wire n_6145;
wire n_11789;
wire n_8699;
wire n_14946;
wire n_7305;
wire n_13878;
wire n_10242;
wire n_10086;
wire n_9992;
wire n_12885;
wire n_14899;
wire n_11347;
wire n_4057;
wire n_14166;
wire n_4332;
wire n_4314;
wire n_7980;
wire n_14363;
wire n_3809;
wire n_11617;
wire n_14952;
wire n_7075;
wire n_7545;
wire n_11581;
wire n_7846;
wire n_10981;
wire n_6076;
wire n_4288;
wire n_14626;
wire n_8438;
wire n_14831;
wire n_6194;
wire n_10673;
wire n_10869;
wire n_7695;
wire n_5066;
wire n_13850;
wire n_12917;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_8095;
wire n_12616;
wire n_7537;
wire n_13690;
wire n_14356;
wire n_14429;
wire n_14705;
wire n_10128;
wire n_10746;
wire n_12217;
wire n_12287;
wire n_12950;
wire n_7489;
wire n_5106;
wire n_10339;
wire n_11559;
wire n_14629;
wire n_5468;
wire n_11867;
wire n_4265;
wire n_6335;
wire n_8112;
wire n_12835;
wire n_14727;
wire n_14343;
wire n_5883;
wire n_6985;
wire n_8642;
wire n_5319;
wire n_14996;
wire n_15072;
wire n_13552;
wire n_13432;
wire n_7451;
wire n_8624;
wire n_6238;
wire n_9090;
wire n_14066;
wire n_11989;
wire n_12800;
wire n_13495;
wire n_10684;
wire n_15030;
wire n_10441;
wire n_12036;
wire n_12177;
wire n_9149;
wire n_10590;
wire n_9174;
wire n_12850;
wire n_11175;
wire n_12962;
wire n_3705;
wire n_6548;
wire n_14755;
wire n_4705;
wire n_5455;
wire n_8894;
wire n_9226;
wire n_6366;
wire n_3778;
wire n_5337;
wire n_5706;
wire n_9018;
wire n_12336;
wire n_10949;
wire n_3912;
wire n_7236;
wire n_9835;
wire n_12044;
wire n_11727;
wire n_12905;
wire n_7269;
wire n_4604;
wire n_8878;
wire n_5223;
wire n_10934;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_14018;
wire n_6620;
wire n_6502;
wire n_9702;
wire n_13409;
wire n_7560;
wire n_11725;
wire n_10279;
wire n_11291;
wire n_7326;
wire n_13548;
wire n_7060;
wire n_7572;
wire n_6885;
wire n_12495;
wire n_13139;
wire n_4217;
wire n_4395;
wire n_8807;
wire n_14207;
wire n_12565;
wire n_9968;
wire n_5074;
wire n_5364;
wire n_9924;
wire n_6529;
wire n_8732;
wire n_8169;
wire n_11958;
wire n_3728;
wire n_8803;
wire n_9515;
wire n_8017;
wire n_10527;
wire n_13506;
wire n_5895;
wire n_4639;
wire n_14756;
wire n_6951;
wire n_3713;
wire n_8801;
wire n_3663;
wire n_12584;
wire n_5649;
wire n_14258;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_12654;
wire n_13255;
wire n_6423;
wire n_9252;
wire n_15017;
wire n_14938;
wire n_10785;
wire n_7140;
wire n_7233;
wire n_10228;
wire n_11311;
wire n_12999;
wire n_14084;
wire n_13120;
wire n_5088;
wire n_6558;
wire n_8522;
wire n_5457;
wire n_7352;
wire n_7986;
wire n_9948;
wire n_7134;
wire n_5532;
wire n_12823;
wire n_11528;
wire n_12422;
wire n_6950;
wire n_7246;
wire n_12234;
wire n_6525;
wire n_7650;
wire n_9871;
wire n_11807;
wire n_14907;
wire n_6631;
wire n_6892;
wire n_11705;
wire n_8203;
wire n_14587;
wire n_7663;
wire n_13125;
wire n_9423;
wire n_11378;
wire n_11521;
wire n_11998;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_9660;
wire n_14513;
wire n_9108;
wire n_14472;
wire n_11222;
wire n_15015;
wire n_4780;
wire n_14910;
wire n_8680;
wire n_9631;
wire n_10643;
wire n_7056;
wire n_4243;
wire n_14590;
wire n_4982;
wire n_12293;
wire n_10427;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_8727;
wire n_10389;
wire n_13069;
wire n_13254;
wire n_10423;
wire n_6292;
wire n_5544;
wire n_15094;
wire n_3832;
wire n_9900;
wire n_14042;
wire n_11080;
wire n_7729;
wire n_3987;
wire n_7339;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_14409;
wire n_4991;
wire n_11533;
wire n_12572;
wire n_5538;
wire n_8138;
wire n_6658;
wire n_10863;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_6925;
wire n_8990;
wire n_5919;
wire n_10077;
wire n_12988;
wire n_8206;
wire n_9144;
wire n_12512;
wire n_7767;
wire n_11940;
wire n_13736;
wire n_8190;
wire n_6176;
wire n_13727;
wire n_9778;
wire n_8622;
wire n_13352;
wire n_5410;
wire n_11808;
wire n_13986;
wire n_7146;
wire n_15035;
wire n_8092;
wire n_13953;
wire n_3937;
wire n_10250;
wire n_6124;
wire n_7672;
wire n_14251;
wire n_8242;
wire n_4525;
wire n_12118;
wire n_12609;
wire n_14053;
wire n_14494;
wire n_3782;
wire n_7482;
wire n_12176;
wire n_9850;
wire n_14503;
wire n_14940;
wire n_6864;
wire n_9531;
wire n_13453;
wire n_7893;
wire n_4208;
wire n_8331;
wire n_7090;
wire n_3786;
wire n_11549;
wire n_7158;
wire n_14174;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_8649;
wire n_8684;
wire n_6494;
wire n_5503;
wire n_8323;
wire n_10828;
wire n_4177;
wire n_12353;
wire n_6199;
wire n_11139;
wire n_8296;
wire n_3763;
wire n_13846;
wire n_9139;
wire n_11584;
wire n_9430;
wire n_10417;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_15059;
wire n_11695;
wire n_7839;
wire n_4264;
wire n_8882;
wire n_10310;
wire n_12053;
wire n_7504;
wire n_10333;
wire n_13316;
wire n_10996;
wire n_13583;
wire n_12795;
wire n_9272;
wire n_8708;
wire n_10880;
wire n_12045;
wire n_7360;
wire n_10810;
wire n_12274;
wire n_7681;
wire n_10636;
wire n_12348;
wire n_8448;
wire n_8076;
wire n_7301;
wire n_9041;
wire n_11360;
wire n_5129;
wire n_11886;
wire n_9643;
wire n_8904;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_11920;
wire n_4276;
wire n_7794;
wire n_11479;
wire n_13388;
wire n_12006;
wire n_7366;
wire n_8184;
wire n_13344;
wire n_5219;
wire n_13336;
wire n_14516;
wire n_5605;
wire n_9944;
wire n_14103;
wire n_5170;
wire n_5654;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_13915;
wire n_14935;
wire n_10258;
wire n_6947;
wire n_11534;
wire n_8586;
wire n_5107;
wire n_9648;
wire n_5999;
wire n_4485;
wire n_8557;
wire n_9376;
wire n_10507;
wire n_8636;
wire n_7309;
wire n_13885;
wire n_4626;
wire n_6863;
wire n_9288;
wire n_10835;
wire n_6637;
wire n_6100;
wire n_13259;
wire n_7860;
wire n_6735;
wire n_14815;
wire n_9521;
wire n_9541;
wire n_13477;
wire n_8212;
wire n_6358;
wire n_4975;
wire n_9759;
wire n_14737;
wire n_12500;
wire n_12781;
wire n_13204;
wire n_7911;
wire n_13085;
wire n_11848;
wire n_8530;
wire n_9278;
wire n_9378;
wire n_11227;
wire n_8665;
wire n_5602;
wire n_9456;
wire n_13778;
wire n_9086;
wire n_7876;
wire n_6050;
wire n_11401;
wire n_14925;
wire n_9711;
wire n_8933;
wire n_14805;
wire n_13206;
wire n_7244;
wire n_7960;
wire n_5405;
wire n_13462;
wire n_12922;
wire n_14123;
wire n_3985;
wire n_5253;
wire n_9485;
wire n_4760;
wire n_11375;
wire n_4652;
wire n_4624;
wire n_9555;
wire n_10959;
wire n_7610;
wire n_12842;
wire n_9999;
wire n_11813;
wire n_14353;
wire n_9994;
wire n_10814;
wire n_5903;
wire n_6371;
wire n_8690;
wire n_8538;
wire n_7043;
wire n_12753;
wire n_10859;
wire n_6171;
wire n_7751;
wire n_8643;
wire n_6510;
wire n_4569;
wire n_6468;
wire n_9142;
wire n_9613;
wire n_11134;
wire n_4897;
wire n_9440;
wire n_5491;
wire n_8825;
wire n_11716;
wire n_12366;
wire n_3940;
wire n_7788;
wire n_14548;
wire n_5842;
wire n_6352;
wire n_8300;
wire n_13954;
wire n_10531;
wire n_14419;
wire n_5722;
wire n_7534;
wire n_9462;
wire n_5636;
wire n_7719;
wire n_11357;
wire n_9202;
wire n_5065;
wire n_7287;
wire n_10699;
wire n_12208;
wire n_7032;
wire n_8451;
wire n_11386;
wire n_13383;
wire n_3637;
wire n_14161;
wire n_4523;
wire n_5492;
wire n_9237;
wire n_10941;
wire n_11448;
wire n_5084;
wire n_10567;
wire n_6850;
wire n_8435;
wire n_5667;
wire n_12122;
wire n_14600;
wire n_10770;
wire n_5260;
wire n_11693;
wire n_7119;
wire n_8835;
wire n_4919;
wire n_13728;
wire n_15038;
wire n_10714;
wire n_9788;
wire n_13584;
wire n_4025;
wire n_13722;
wire n_5328;
wire n_14060;
wire n_14936;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_14634;
wire n_11755;
wire n_4503;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_11221;
wire n_7851;
wire n_6332;
wire n_9807;
wire n_14613;
wire n_13567;
wire n_4464;
wire n_13642;
wire n_7006;
wire n_9573;
wire n_5877;
wire n_8963;
wire n_12351;
wire n_6306;
wire n_7682;
wire n_4114;
wire n_14297;
wire n_13618;
wire n_6434;
wire n_12040;
wire n_12443;
wire n_8713;
wire n_6751;
wire n_7068;
wire n_9392;
wire n_12133;
wire n_4556;
wire n_11084;
wire n_13371;
wire n_14573;
wire n_6322;
wire n_14048;
wire n_8353;
wire n_8668;
wire n_13301;
wire n_5454;
wire n_9390;
wire n_13492;
wire n_14376;
wire n_7704;
wire n_10326;
wire n_7773;
wire n_9416;
wire n_14728;
wire n_6667;
wire n_7526;
wire n_13333;
wire n_8817;
wire n_6530;
wire n_9518;
wire n_4089;
wire n_13329;
wire n_12491;
wire n_7376;
wire n_13826;
wire n_6156;
wire n_13966;
wire n_14498;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_12452;
wire n_5621;
wire n_13788;
wire n_13437;
wire n_8213;
wire n_12233;
wire n_4327;
wire n_8591;
wire n_7973;
wire n_11885;
wire n_4218;
wire n_6429;
wire n_13423;
wire n_10966;
wire n_5165;
wire n_7239;
wire n_10047;
wire n_12633;
wire n_5573;
wire n_11253;
wire n_6405;
wire n_11551;
wire n_14761;
wire n_8532;
wire n_11380;
wire n_12936;
wire n_12035;
wire n_13928;
wire n_6613;
wire n_4353;
wire n_8043;
wire n_9196;
wire n_11172;
wire n_13947;
wire n_14420;
wire n_7969;
wire n_6248;
wire n_14059;
wire n_12915;
wire n_7821;
wire n_4990;
wire n_6088;
wire n_12275;
wire n_10784;
wire n_5529;
wire n_10248;
wire n_6894;
wire n_12947;
wire n_14678;
wire n_7267;
wire n_4959;
wire n_9589;
wire n_4161;
wire n_5800;
wire n_11539;
wire n_9898;
wire n_14520;
wire n_13257;
wire n_9373;
wire n_3992;
wire n_11976;
wire n_12308;
wire n_13063;
wire n_8606;
wire n_14669;
wire n_4103;
wire n_4466;
wire n_6204;
wire n_10351;
wire n_13834;
wire n_13951;
wire n_7915;
wire n_8121;
wire n_8868;
wire n_10408;
wire n_10921;
wire n_13340;
wire n_7387;
wire n_7431;
wire n_11731;
wire n_7654;
wire n_10551;
wire n_12760;
wire n_10656;
wire n_4844;
wire n_6296;
wire n_11531;
wire n_12318;
wire n_13379;
wire n_10313;
wire n_10639;
wire n_5257;
wire n_9983;
wire n_6290;
wire n_14983;
wire n_6288;
wire n_3655;
wire n_12700;
wire n_4688;
wire n_14517;
wire n_4765;
wire n_8276;
wire n_8718;
wire n_12364;
wire n_8182;
wire n_5645;
wire n_14512;
wire n_11392;
wire n_5180;
wire n_13490;
wire n_11204;
wire n_3640;
wire n_13025;
wire n_13672;
wire n_13754;
wire n_14785;
wire n_12985;
wire n_5779;
wire n_11627;
wire n_13697;
wire n_4388;
wire n_4206;
wire n_12340;
wire n_12478;
wire n_6140;
wire n_9039;
wire n_13744;
wire n_8359;
wire n_7441;
wire n_9849;
wire n_8597;
wire n_4738;
wire n_6211;
wire n_12788;
wire n_8562;
wire n_13470;
wire n_3909;
wire n_11485;
wire n_8211;
wire n_13998;
wire n_13943;
wire n_9962;
wire n_14814;
wire n_12826;
wire n_8430;
wire n_6307;
wire n_8007;
wire n_10871;
wire n_6164;
wire n_3944;
wire n_12752;
wire n_7394;
wire n_8600;
wire n_8311;
wire n_8943;
wire n_8441;
wire n_12194;
wire n_4434;
wire n_4837;
wire n_10747;
wire n_7022;
wire n_9829;
wire n_14772;
wire n_13637;
wire n_6860;
wire n_4219;
wire n_10459;
wire n_3659;
wire n_8978;
wire n_5012;
wire n_10121;
wire n_4620;
wire n_11387;
wire n_8198;
wire n_9988;
wire n_14417;
wire n_5697;
wire n_14652;
wire n_14002;
wire n_7188;
wire n_8526;
wire n_10705;
wire n_13099;
wire n_7573;
wire n_7879;
wire n_4438;
wire n_9848;
wire n_7087;
wire n_6147;
wire n_14911;
wire n_10334;
wire n_7985;
wire n_12689;
wire n_11691;
wire n_11358;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_15021;
wire n_9348;
wire n_6011;
wire n_8278;
wire n_7722;
wire n_7935;
wire n_8592;
wire n_6645;
wire n_11128;
wire n_12271;
wire n_13595;
wire n_14358;
wire n_14006;
wire n_8226;
wire n_6984;
wire n_4325;
wire n_12843;
wire n_13780;
wire n_10716;
wire n_12273;
wire n_10235;
wire n_13212;
wire n_13701;
wire n_10090;
wire n_13247;
wire n_10153;
wire n_14271;
wire n_11649;
wire n_10937;
wire n_13922;
wire n_7193;
wire n_10018;
wire n_13278;
wire n_8987;
wire n_13836;
wire n_4133;
wire n_3775;
wire n_11489;
wire n_6897;
wire n_7256;
wire n_12391;
wire n_4184;
wire n_5203;
wire n_12420;
wire n_14181;
wire n_9071;
wire n_10568;
wire n_9356;
wire n_9464;
wire n_4481;
wire n_12314;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_9239;
wire n_10053;
wire n_6183;
wire n_10051;
wire n_11373;
wire n_7522;
wire n_5882;
wire n_13341;
wire n_9606;
wire n_13856;
wire n_4030;
wire n_10359;
wire n_7881;
wire n_14416;
wire n_14796;
wire n_14961;
wire n_7436;
wire n_4490;
wire n_7380;
wire n_7012;
wire n_11216;
wire n_4397;
wire n_12356;
wire n_10998;
wire n_7502;
wire n_9492;
wire n_13271;
wire n_8960;
wire n_7335;
wire n_7103;
wire n_13553;
wire n_4820;
wire n_10648;
wire n_10151;
wire n_6246;
wire n_14602;
wire n_14133;
wire n_11194;
wire n_11804;
wire n_3770;
wire n_8025;
wire n_5094;
wire n_6383;
wire n_9031;
wire n_11107;
wire n_4938;
wire n_9717;
wire n_11434;
wire n_9516;
wire n_11645;
wire n_12073;
wire n_7020;
wire n_8434;
wire n_4179;
wire n_11244;
wire n_12848;
wire n_8175;
wire n_9991;
wire n_9693;
wire n_5336;
wire n_12155;
wire n_13356;
wire n_14286;
wire n_9103;
wire n_8850;
wire n_11254;
wire n_14865;
wire n_13693;
wire n_9477;
wire n_14277;
wire n_5672;
wire n_4641;
wire n_13673;
wire n_5548;
wire n_10253;
wire n_10822;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_14793;
wire n_8895;
wire n_3855;
wire n_10589;
wire n_12390;
wire n_12160;
wire n_13501;
wire n_11297;
wire n_10349;
wire n_11991;
wire n_5339;
wire n_13376;
wire n_4931;
wire n_6099;
wire n_10946;
wire n_12150;
wire n_5693;
wire n_8046;
wire n_11183;
wire n_11173;
wire n_6904;
wire n_3760;
wire n_4078;
wire n_11922;
wire n_13897;
wire n_8867;
wire n_10473;
wire n_8239;
wire n_9599;
wire n_13104;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_7825;
wire n_8183;
wire n_8924;
wire n_9001;
wire n_12840;
wire n_10893;
wire n_3828;
wire n_13215;
wire n_10218;
wire n_13482;
wire n_12964;
wire n_5514;
wire n_13075;
wire n_5091;
wire n_4404;
wire n_7533;
wire n_8578;
wire n_11548;
wire n_9777;
wire n_4787;
wire n_8848;
wire n_10903;
wire n_13445;
wire n_3667;
wire n_10458;
wire n_11868;
wire n_13562;
wire n_9222;
wire n_10148;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_9366;
wire n_6611;
wire n_10775;
wire n_11248;
wire n_10543;
wire n_9449;
wire n_3703;
wire n_4903;
wire n_15098;
wire n_11114;
wire n_11260;
wire n_11901;
wire n_12994;
wire n_5599;
wire n_14771;
wire n_6116;
wire n_7186;
wire n_10337;
wire n_4356;
wire n_8230;
wire n_9869;
wire n_10478;
wire n_12252;
wire n_11981;
wire n_6819;
wire n_8725;
wire n_4432;
wire n_13929;
wire n_5251;
wire n_7936;
wire n_13534;
wire n_13680;
wire n_6473;
wire n_12951;
wire n_13750;
wire n_9741;
wire n_13275;
wire n_4291;
wire n_11956;
wire n_10956;
wire n_10637;
wire n_13331;
wire n_13536;
wire n_11805;
wire n_15043;
wire n_5403;
wire n_4386;
wire n_12131;
wire n_12280;
wire n_4149;
wire n_8391;
wire n_6310;
wire n_7840;
wire n_10698;
wire n_11381;
wire n_14607;
wire n_9397;
wire n_8202;
wire n_11797;
wire n_11775;
wire n_12453;
wire n_10834;
wire n_7429;
wire n_6688;
wire n_12557;
wire n_7906;
wire n_8948;
wire n_8678;
wire n_9754;
wire n_4019;
wire n_10783;
wire n_9179;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7658;
wire n_7462;
wire n_7828;
wire n_8340;
wire n_8905;
wire n_12020;
wire n_13439;
wire n_4935;
wire n_8691;
wire n_13249;
wire n_12051;
wire n_6365;
wire n_10619;
wire n_14225;
wire n_4785;
wire n_3820;
wire n_13502;
wire n_13801;
wire n_5608;
wire n_13468;
wire n_3741;
wire n_11322;
wire n_12455;
wire n_10136;
wire n_7401;
wire n_13789;
wire n_8812;
wire n_12920;
wire n_14759;
wire n_13403;
wire n_9169;
wire n_6828;
wire n_12785;
wire n_14200;
wire n_11758;
wire n_5298;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_11162;
wire n_13996;
wire n_8058;
wire n_4413;
wire n_12559;
wire n_9177;
wire n_10078;
wire n_6777;
wire n_5728;
wire n_11987;
wire n_8394;
wire n_9269;
wire n_3990;
wire n_4493;
wire n_7835;
wire n_10719;
wire n_12614;
wire n_13201;
wire n_14638;
wire n_11106;
wire n_9289;
wire n_8181;
wire n_10463;
wire n_12797;
wire n_13737;
wire n_13441;
wire n_14396;
wire n_14687;
wire n_8722;
wire n_10827;
wire n_12429;
wire n_6420;
wire n_6945;
wire n_11218;
wire n_9350;
wire n_7356;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_11467;
wire n_7124;
wire n_10454;
wire n_12668;
wire n_12384;
wire n_3672;
wire n_7294;
wire n_12629;
wire n_13291;
wire n_12123;
wire n_5290;
wire n_12972;
wire n_14969;
wire n_7018;
wire n_13105;
wire n_10312;
wire n_11374;
wire n_11167;
wire n_13440;
wire n_12146;
wire n_7321;
wire n_9166;
wire n_10663;
wire n_10501;
wire n_5095;
wire n_10265;
wire n_10452;
wire n_8707;
wire n_6754;
wire n_10766;
wire n_12435;
wire n_13533;
wire n_11999;
wire n_6583;
wire n_13367;
wire n_6622;
wire n_6936;
wire n_13123;
wire n_8747;
wire n_5324;
wire n_3897;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_8742;
wire n_10470;
wire n_10563;
wire n_12921;
wire n_7108;
wire n_6882;
wire n_11455;
wire n_7585;
wire n_13930;
wire n_9125;
wire n_7386;
wire n_4570;
wire n_8552;
wire n_10288;
wire n_5101;
wire n_12581;
wire n_5019;
wire n_5911;
wire n_4296;
wire n_7362;
wire n_7888;
wire n_7417;
wire n_12029;
wire n_12548;
wire n_9641;
wire n_14460;
wire n_9960;
wire n_7187;
wire n_13111;
wire n_11884;
wire n_5589;
wire n_5841;
wire n_13060;
wire n_12727;
wire n_10776;
wire n_11611;
wire n_9785;
wire n_9923;
wire n_8224;
wire n_10771;
wire n_7544;
wire n_11087;
wire n_14556;
wire n_5712;
wire n_11960;
wire n_4606;
wire n_6166;
wire n_8628;
wire n_4774;
wire n_13108;
wire n_11422;
wire n_13948;
wire n_6966;
wire n_13563;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_9228;
wire n_14828;
wire n_7255;
wire n_4093;
wire n_12227;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_7218;
wire n_12597;
wire n_4672;
wire n_7147;
wire n_7221;
wire n_14653;
wire n_15016;
wire n_10967;
wire n_4174;
wire n_8289;
wire n_9801;
wire n_14189;
wire n_10249;
wire n_11029;
wire n_15057;
wire n_9645;
wire n_4766;
wire n_8045;
wire n_11199;
wire n_5633;
wire n_8697;
wire n_13568;
wire n_13396;
wire n_13029;
wire n_13647;
wire n_8077;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_12674;
wire n_5583;
wire n_11826;
wire n_9457;
wire n_15071;
wire n_4460;
wire n_8026;
wire n_11317;
wire n_3645;
wire n_13652;
wire n_7889;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_10742;
wire n_6237;
wire n_14538;
wire n_7196;
wire n_12913;
wire n_10390;
wire n_9330;
wire n_6341;
wire n_10012;
wire n_9365;
wire n_14861;
wire n_6590;
wire n_5501;
wire n_8444;
wire n_9178;
wire n_8654;
wire n_14021;
wire n_10035;
wire n_10753;
wire n_9181;
wire n_12112;
wire n_7923;
wire n_13965;
wire n_3938;
wire n_14465;
wire n_5377;
wire n_11033;
wire n_6697;
wire n_13168;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_13574;
wire n_14037;
wire n_7559;
wire n_11798;
wire n_12346;
wire n_4110;
wire n_11853;
wire n_7081;
wire n_9307;
wire n_10795;
wire n_10300;
wire n_10257;
wire n_6449;
wire n_7832;
wire n_7968;
wire n_9238;
wire n_12714;
wire n_11079;
wire n_11166;
wire n_13581;
wire n_6141;
wire n_10099;
wire n_8449;
wire n_11217;
wire n_12732;
wire n_13138;
wire n_14481;
wire n_3965;
wire n_10985;
wire n_4349;
wire n_14931;
wire n_8493;
wire n_7584;
wire n_9224;
wire n_3788;
wire n_10244;
wire n_12400;
wire n_4313;
wire n_6983;
wire n_12671;
wire n_7843;
wire n_13774;
wire n_10377;
wire n_6036;
wire n_11469;
wire n_10984;
wire n_12863;
wire n_12347;
wire n_8958;
wire n_10801;
wire n_11898;
wire n_8443;
wire n_4863;
wire n_12041;
wire n_9756;
wire n_7222;
wire n_9624;
wire n_6071;
wire n_8161;
wire n_13435;
wire n_11710;
wire n_6808;
wire n_8734;
wire n_9547;
wire n_11341;
wire n_8271;
wire n_9901;
wire n_9594;
wire n_11619;
wire n_11238;
wire n_9895;
wire n_10878;
wire n_13378;
wire n_6724;
wire n_3995;
wire n_9277;
wire n_11608;
wire n_14169;
wire n_4036;
wire n_14086;
wire n_12756;
wire n_6571;
wire n_15074;
wire n_5100;
wire n_7470;
wire n_9189;
wire n_5849;
wire n_8495;
wire n_6251;
wire n_7400;
wire n_14255;
wire n_9548;
wire n_14309;
wire n_12088;
wire n_12218;
wire n_14204;
wire n_6635;
wire n_10000;
wire n_3894;
wire n_9472;
wire n_13202;
wire n_14738;
wire n_13410;
wire n_11553;
wire n_4015;
wire n_14432;
wire n_3890;
wire n_5367;
wire n_13816;
wire n_8994;
wire n_8901;
wire n_8056;
wire n_10725;
wire n_12323;
wire n_14767;
wire n_9538;
wire n_7623;
wire n_12387;
wire n_14984;
wire n_10627;
wire n_8954;
wire n_13590;
wire n_5616;
wire n_13230;
wire n_7597;
wire n_11996;
wire n_5034;
wire n_6733;
wire n_7071;
wire n_15029;
wire n_8840;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_7859;
wire n_8900;
wire n_13456;
wire n_10477;
wire n_14651;
wire n_13321;
wire n_12798;
wire n_14306;
wire n_11032;
wire n_6522;
wire n_7109;
wire n_11834;
wire n_14057;
wire n_9434;
wire n_10604;
wire n_11110;
wire n_5959;
wire n_9052;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_13806;
wire n_4807;
wire n_6562;
wire n_12780;
wire n_6150;
wire n_9176;
wire n_10461;
wire n_12772;
wire n_10559;
wire n_11141;
wire n_8157;
wire n_12539;
wire n_13007;
wire n_8346;
wire n_9697;
wire n_4230;
wire n_13651;
wire n_7882;
wire n_13830;
wire n_8827;
wire n_13113;
wire n_8309;
wire n_13196;
wire n_14998;
wire n_8344;
wire n_5917;
wire n_12589;
wire n_9060;
wire n_5754;
wire n_6016;
wire n_12775;
wire n_8096;
wire n_8100;
wire n_8822;
wire n_3784;
wire n_3941;
wire n_12043;
wire n_9758;
wire n_7212;
wire n_3678;
wire n_7908;
wire n_8222;
wire n_14430;
wire n_10479;
wire n_9876;
wire n_5628;
wire n_10572;
wire n_11971;
wire n_6726;
wire n_8406;
wire n_10277;
wire n_11320;
wire n_14697;
wire n_4428;
wire n_5003;
wire n_11028;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_10139;
wire n_10230;
wire n_14294;
wire n_6689;
wire n_14245;
wire n_12476;
wire n_14858;
wire n_8866;
wire n_13724;
wire n_6143;
wire n_5614;
wire n_8693;
wire n_5134;
wire n_3953;
wire n_10207;
wire n_12536;
wire n_4122;
wire n_3976;
wire n_11368;
wire n_11144;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_7777;
wire n_8794;
wire n_6277;
wire n_9653;
wire n_7395;
wire n_4684;
wire n_5981;
wire n_11404;
wire n_14993;
wire n_12896;
wire n_13373;
wire n_6095;
wire n_7671;
wire n_10429;
wire n_8020;
wire n_14241;
wire n_12957;
wire n_13866;
wire n_6247;
wire n_4840;
wire n_10255;
wire n_9257;
wire n_13014;
wire n_9270;
wire n_6880;
wire n_10901;
wire n_3749;
wire n_10101;
wire n_5720;
wire n_3962;
wire n_14000;
wire n_13022;
wire n_13422;
wire n_5325;
wire n_13633;
wire n_5696;
wire n_12549;
wire n_5375;
wire n_4384;
wire n_8736;
wire n_6499;
wire n_12362;
wire n_6837;
wire n_13442;
wire n_14741;
wire n_14972;
wire n_15073;
wire n_4423;
wire n_10063;
wire n_13390;
wire n_4096;
wire n_12030;
wire n_7393;
wire n_8400;
wire n_6616;
wire n_9686;
wire n_13136;
wire n_13334;
wire n_13408;
wire n_13989;
wire n_14690;
wire n_7871;
wire n_14532;
wire n_14859;
wire n_12018;
wire n_10846;
wire n_6946;
wire n_4996;
wire n_8055;
wire n_8333;
wire n_10195;
wire n_11593;
wire n_11847;
wire n_9718;
wire n_11773;
wire n_4598;
wire n_14074;
wire n_14944;
wire n_5064;
wire n_9215;
wire n_5759;
wire n_12060;
wire n_4478;
wire n_5753;
wire n_10628;
wire n_8909;
wire n_5536;
wire n_15056;
wire n_7484;
wire n_5173;
wire n_11968;
wire n_6305;
wire n_13630;
wire n_14071;
wire n_14127;
wire n_6317;
wire n_3920;
wire n_9762;
wire n_9407;
wire n_10819;
wire n_12315;
wire n_12903;
wire n_4890;
wire n_13269;
wire n_14570;
wire n_5691;
wire n_13103;
wire n_5794;
wire n_13098;
wire n_11896;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_11897;
wire n_14447;
wire n_13707;
wire n_10368;
wire n_12484;
wire n_3866;
wire n_14971;
wire n_3921;
wire n_7272;
wire n_9964;
wire n_4106;
wire n_3717;
wire n_13031;
wire n_13646;
wire n_5738;
wire n_7649;
wire n_9953;
wire n_10356;
wire n_14154;
wire n_5215;
wire n_7324;
wire n_9153;
wire n_6693;
wire n_8786;
wire n_10931;
wire n_8541;
wire n_11711;
wire n_3743;
wire n_12673;
wire n_6734;
wire n_12000;
wire n_10173;
wire n_9571;
wire n_7135;
wire n_11554;
wire n_7014;
wire n_8263;
wire n_10644;
wire n_11159;
wire n_8884;
wire n_5597;
wire n_4721;
wire n_13062;
wire n_5635;
wire n_13424;
wire n_10323;
wire n_11350;
wire n_6382;
wire n_9019;
wire n_11310;
wire n_13001;
wire n_7328;
wire n_7635;
wire n_6404;
wire n_12063;
wire n_15023;
wire n_10229;
wire n_10693;
wire n_5975;
wire n_9737;
wire n_4029;
wire n_11688;
wire n_13842;
wire n_10493;
wire n_11125;
wire n_8494;
wire n_10554;
wire n_3870;
wire n_6379;
wire n_10382;
wire n_11083;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_7358;
wire n_9468;
wire n_10622;
wire n_12449;
wire n_13664;
wire n_11939;
wire n_6235;
wire n_13144;
wire n_9870;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_9026;
wire n_13900;
wire n_9710;
wire n_3952;
wire n_7265;
wire n_8638;
wire n_11126;
wire n_8710;
wire n_10019;
wire n_13512;
wire n_6789;
wire n_7184;
wire n_11090;
wire n_6440;
wire n_9725;
wire n_11953;
wire n_6417;
wire n_12845;
wire n_14557;
wire n_8177;
wire n_14013;
wire n_12062;
wire n_12636;
wire n_14784;
wire n_7491;
wire n_4495;
wire n_4762;
wire n_5942;
wire n_14436;
wire n_14524;
wire n_9084;
wire n_7728;
wire n_10488;
wire n_10767;
wire n_7690;
wire n_13084;
wire n_7219;
wire n_13375;
wire n_7479;
wire n_11040;
wire n_13852;
wire n_3998;
wire n_11751;
wire n_9419;
wire n_12793;
wire n_13203;
wire n_14378;
wire n_4141;
wire n_11158;
wire n_14488;
wire n_7270;
wire n_5940;
wire n_8170;
wire n_12367;
wire n_10579;
wire n_8893;
wire n_13473;
wire n_14923;
wire n_12317;
wire n_7390;
wire n_7805;
wire n_10474;
wire n_7807;
wire n_5121;
wire n_9973;
wire n_8589;
wire n_4107;
wire n_9820;
wire n_9479;
wire n_12724;
wire n_12954;
wire n_4667;
wire n_11094;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_12157;
wire n_14891;
wire n_11161;
wire n_11182;
wire n_10587;
wire n_7182;
wire n_12195;
wire n_4547;
wire n_11839;
wire n_11815;
wire n_5784;
wire n_4004;
wire n_10843;
wire n_12773;
wire n_6272;
wire n_8153;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_12556;
wire n_6236;
wire n_8620;
wire n_10755;
wire n_5576;
wire n_4668;
wire n_8298;
wire n_11614;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_13645;
wire n_3898;
wire n_6871;
wire n_12789;
wire n_10270;
wire n_11590;
wire n_12649;
wire n_8235;
wire n_11845;
wire n_5284;
wire n_9294;
wire n_9126;
wire n_8370;
wire n_13773;
wire n_11263;
wire n_11908;
wire n_4997;
wire n_13066;
wire n_5308;
wire n_4274;
wire n_13469;
wire n_10573;
wire n_13101;
wire n_6768;
wire n_4759;
wire n_13494;
wire n_13893;
wire n_7951;
wire n_10992;
wire n_14490;
wire n_4467;
wire n_7506;
wire n_14210;
wire n_14717;
wire n_12696;
wire n_6717;
wire n_13505;
wire n_11257;
wire n_3684;
wire n_4735;
wire n_7048;
wire n_11136;
wire n_11142;
wire n_10428;
wire n_13569;
wire n_12664;
wire n_5578;
wire n_8395;
wire n_10989;
wire n_13450;
wire n_11145;
wire n_12206;
wire n_11745;
wire n_13010;
wire n_15081;
wire n_14375;
wire n_13181;
wire n_11017;
wire n_4113;
wire n_10805;
wire n_8906;
wire n_4686;
wire n_5530;
wire n_10682;
wire n_11414;
wire n_8097;
wire n_10327;
wire n_12940;
wire n_3759;
wire n_14322;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_10528;
wire n_5741;
wire n_8570;
wire n_8902;
wire n_12404;
wire n_5991;
wire n_13815;
wire n_3933;
wire n_10365;
wire n_7330;
wire n_7928;
wire n_12201;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_15061;
wire n_9819;
wire n_8477;
wire n_5449;
wire n_10236;
wire n_5221;
wire n_6992;
wire n_10433;
wire n_13725;
wire n_13924;
wire n_4183;
wire n_12312;
wire n_4068;
wire n_4872;
wire n_10625;
wire n_6000;
wire n_10303;
wire n_9545;
wire n_4233;
wire n_7283;
wire n_7099;
wire n_3764;
wire n_11452;
wire n_10557;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_11323;
wire n_13002;
wire n_6655;
wire n_12982;
wire n_7892;
wire n_9165;
wire n_11558;
wire n_14732;
wire n_7304;
wire n_10143;
wire n_13018;
wire n_5792;
wire n_13185;
wire n_14872;
wire n_14681;
wire n_12002;
wire n_6657;
wire n_7756;
wire n_8129;
wire n_13150;
wire n_5575;
wire n_8580;
wire n_11543;
wire n_7990;
wire n_3914;
wire n_4625;
wire n_8122;
wire n_11883;
wire n_10796;
wire n_8259;
wire n_3803;
wire n_8536;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_10855;
wire n_8748;
wire n_7612;
wire n_6113;
wire n_7789;
wire n_4819;
wire n_9056;
wire n_8094;
wire n_9341;
wire n_14164;
wire n_11429;
wire n_14165;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_15027;
wire n_6519;
wire n_10357;
wire n_8572;
wire n_4900;
wire n_10681;
wire n_8120;
wire n_12598;
wire n_6842;
wire n_12942;
wire n_12750;
wire n_13575;
wire n_12729;
wire n_7588;
wire n_12033;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_11241;
wire n_9172;
wire n_14239;
wire n_3817;
wire n_12441;
wire n_9145;
wire n_13805;
wire n_6801;
wire n_8099;
wire n_9996;
wire n_11348;
wire n_10059;
wire n_10284;
wire n_4930;
wire n_7680;
wire n_8770;
wire n_5276;
wire n_6308;
wire n_14790;
wire n_7398;
wire n_6906;
wire n_14029;
wire n_5078;
wire n_11169;
wire n_4537;
wire n_11041;
wire n_7230;
wire n_8700;
wire n_11160;
wire n_9906;
wire n_6629;
wire n_5011;
wire n_10957;
wire n_14250;
wire n_12827;
wire n_4070;
wire n_11124;
wire n_6968;
wire n_9920;
wire n_4282;
wire n_9504;
wire n_6615;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_12734;
wire n_12181;
wire n_9482;
wire n_5205;
wire n_14032;
wire n_14760;
wire n_9138;
wire n_11152;
wire n_9384;
wire n_8637;
wire n_5651;
wire n_6144;
wire n_8757;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_14794;
wire n_5819;
wire n_10147;
wire n_14197;
wire n_4579;
wire n_4616;
wire n_13765;
wire n_8903;
wire n_13709;
wire n_9193;
wire n_5998;
wire n_6398;
wire n_11586;
wire n_14660;
wire n_5023;
wire n_12069;
wire n_11990;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_9527;
wire n_14554;
wire n_3791;
wire n_5351;
wire n_3905;
wire n_10889;
wire n_12363;
wire n_11019;
wire n_14028;
wire n_13170;
wire n_14368;
wire n_14699;
wire n_8585;
wire n_9064;
wire n_14056;
wire n_8982;
wire n_6415;
wire n_10816;
wire n_14374;
wire n_10032;
wire n_13385;
wire n_6857;
wire n_10489;
wire n_5476;
wire n_10200;
wire n_12442;
wire n_7842;
wire n_10898;
wire n_5856;
wire n_12499;
wire n_14588;
wire n_8709;
wire n_5446;
wire n_9383;
wire n_10825;
wire n_4895;
wire n_6722;
wire n_9735;
wire n_9943;
wire n_10290;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_12818;
wire n_15078;
wire n_6413;
wire n_7679;
wire n_11132;
wire n_4275;
wire n_13684;
wire n_6361;
wire n_3970;
wire n_9357;
wire n_11677;
wire n_13608;
wire n_10680;
wire n_12531;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_11036;
wire n_14826;
wire n_5684;
wire n_5861;
wire n_11927;
wire n_8108;
wire n_10306;
wire n_5976;
wire n_4789;
wire n_11827;
wire n_7862;
wire n_5312;
wire n_10675;
wire n_5850;
wire n_10014;
wire n_13454;
wire n_5111;
wire n_13829;
wire n_5890;
wire n_4055;
wire n_9986;
wire n_10355;
wire n_3670;
wire n_3973;
wire n_13758;
wire n_10830;
wire n_7820;
wire n_7167;
wire n_8692;
wire n_14967;
wire n_7833;
wire n_11118;
wire n_8820;
wire n_12496;
wire n_14750;
wire n_7643;
wire n_12460;
wire n_13586;
wire n_8490;
wire n_10380;
wire n_5113;
wire n_4442;
wire n_9491;
wire n_4698;
wire n_12821;
wire n_15028;
wire n_14809;
wire n_9922;
wire n_6712;
wire n_5687;
wire n_12479;
wire n_10530;
wire n_13703;
wire n_4779;
wire n_8062;
wire n_8781;
wire n_10999;
wire n_10203;
wire n_4966;
wire n_8000;
wire n_10061;
wire n_13860;
wire n_10899;
wire n_10961;
wire n_4017;
wire n_8808;
wire n_13359;
wire n_8233;
wire n_5839;
wire n_3740;
wire n_9747;
wire n_11811;
wire n_6953;
wire n_8685;
wire n_4418;
wire n_13877;
wire n_15097;
wire n_9061;
wire n_9168;
wire n_12361;
wire n_11561;
wire n_12345;
wire n_8575;
wire n_8701;
wire n_11690;
wire n_11212;
wire n_6303;
wire n_12593;
wire n_6474;
wire n_6182;
wire n_3723;
wire n_11155;
wire n_5674;
wire n_8670;
wire n_6573;
wire n_4134;
wire n_13151;
wire n_6053;
wire n_14380;
wire n_7234;
wire n_10425;
wire n_15060;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_5682;
wire n_12984;
wire n_8385;
wire n_14330;
wire n_8875;
wire n_6392;
wire n_8166;
wire n_11433;
wire n_5167;
wire n_9073;
wire n_8934;
wire n_5117;
wire n_3686;
wire n_4913;
wire n_11312;
wire n_11477;
wire n_7999;
wire n_5612;
wire n_14347;
wire n_11988;
wire n_6125;
wire n_6599;
wire n_7963;
wire n_14978;
wire n_6685;
wire n_12311;
wire n_12914;
wire n_11964;
wire n_12086;
wire n_4251;
wire n_8389;
wire n_9068;
wire n_3982;
wire n_10537;
wire n_4621;
wire n_10158;
wire n_14823;
wire n_6560;
wire n_12787;
wire n_14686;
wire n_10711;
wire n_11933;
wire n_8659;
wire n_8804;
wire n_10043;
wire n_4559;
wire n_12703;
wire n_12411;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_8439;
wire n_13337;
wire n_9544;
wire n_14108;
wire n_8814;
wire n_8369;
wire n_13867;
wire n_5301;
wire n_11574;
wire n_7800;
wire n_5007;
wire n_4077;
wire n_7615;
wire n_4642;
wire n_9286;
wire n_5898;
wire n_10930;
wire n_11313;
wire n_14700;
wire n_11206;
wire n_12263;
wire n_7298;
wire n_12959;
wire n_7581;
wire n_10131;
wire n_4049;
wire n_6641;
wire n_5214;
wire n_3862;
wire n_13057;
wire n_13551;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_3879;
wire n_6673;
wire n_10696;
wire n_12461;
wire n_12893;
wire n_13990;
wire n_8789;
wire n_7172;
wire n_7074;
wire n_10685;
wire n_5497;
wire n_8790;
wire n_11223;
wire n_8234;
wire n_11624;
wire n_4724;
wire n_5832;
wire n_13876;
wire n_13791;
wire n_14438;
wire n_7190;
wire n_11515;
wire n_7112;
wire n_14382;
wire n_13128;
wire n_13807;
wire n_13142;
wire n_7678;
wire n_10082;
wire n_9265;
wire n_11560;
wire n_13678;
wire n_9080;
wire n_13433;
wire n_5526;
wire n_8989;
wire n_10152;
wire n_15063;
wire n_13589;
wire n_3646;
wire n_12645;
wire n_6367;
wire n_4546;
wire n_6195;
wire n_6356;
wire n_8927;
wire n_11055;
wire n_14192;
wire n_3756;
wire n_11616;
wire n_9770;
wire n_14746;
wire n_9463;
wire n_7001;
wire n_12090;
wire n_13481;
wire n_13743;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_7369;
wire n_5444;
wire n_10580;
wire n_14365;
wire n_7829;
wire n_14131;
wire n_4382;
wire n_9939;
wire n_10159;
wire n_3999;
wire n_11390;
wire n_8534;
wire n_9911;
wire n_9210;
wire n_5211;
wire n_6559;
wire n_5230;
wire n_10122;
wire n_10302;
wire n_14457;
wire n_7359;
wire n_14398;
wire n_5389;
wire n_7144;
wire n_10462;
wire n_4833;
wire n_14244;
wire n_13357;
wire n_8756;
wire n_6841;
wire n_14320;
wire n_11597;
wire n_14918;
wire n_11002;
wire n_13716;
wire n_9691;
wire n_5110;
wire n_6653;
wire n_12165;
wire n_4719;
wire n_4178;
wire n_7450;
wire n_5425;
wire n_13803;
wire n_14455;
wire n_10532;
wire n_8832;
wire n_5737;
wire n_9340;
wire n_10350;
wire n_9351;
wire n_8461;
wire n_8042;
wire n_11179;
wire n_10977;
wire n_6923;
wire n_6825;
wire n_11708;
wire n_9950;
wire n_10418;
wire n_11474;
wire n_10336;
wire n_4228;
wire n_4401;
wire n_8021;
wire n_8839;
wire n_12092;
wire n_11369;
wire n_6112;
wire n_6547;
wire n_11738;
wire n_11240;
wire n_14113;
wire n_6198;
wire n_13155;
wire n_7439;
wire n_5560;
wire n_12074;
wire n_9155;
wire n_14565;
wire n_11931;
wire n_14231;
wire n_10925;
wire n_6399;
wire n_8623;
wire n_12109;
wire n_11438;
wire n_8758;
wire n_14508;
wire n_6275;
wire n_5666;
wire n_6575;
wire n_10609;
wire n_13508;
wire n_7924;
wire n_7732;
wire n_6151;
wire n_13058;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_15042;
wire n_4877;
wire n_8511;
wire n_7325;
wire n_6469;
wire n_4968;
wire n_6756;
wire n_8595;
wire n_12900;
wire n_8873;
wire n_11376;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_7459;
wire n_7191;
wire n_9201;
wire n_9823;
wire n_11051;
wire n_11812;
wire n_14304;
wire n_9688;
wire n_12330;
wire n_7096;
wire n_12519;
wire n_13872;
wire n_13597;
wire n_8455;
wire n_11838;
wire n_12717;
wire n_8280;
wire n_3903;
wire n_10102;
wire n_4834;
wire n_10908;
wire n_11333;
wire n_9595;
wire n_5272;
wire n_9530;
wire n_6826;
wire n_4158;
wire n_9227;
wire n_6015;
wire n_8372;
wire n_5361;
wire n_8598;
wire n_5683;
wire n_10939;
wire n_4171;
wire n_13503;
wire n_11178;
wire n_12595;
wire n_5847;
wire n_7551;
wire n_9400;
wire n_4045;
wire n_6678;
wire n_11188;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_9025;
wire n_5740;
wire n_13086;
wire n_8282;
wire n_7750;
wire n_10936;
wire n_11840;
wire n_5015;
wire n_12525;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_11685;
wire n_10955;
wire n_13093;
wire n_10824;
wire n_6748;
wire n_12084;
wire n_8616;
wire n_4749;
wire n_10440;
wire n_10630;
wire n_8336;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_11472;
wire n_6752;
wire n_9749;
wire n_14404;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_9285;
wire n_12997;
wire n_11295;
wire n_9972;
wire n_10058;
wire n_7652;
wire n_14533;
wire n_8847;
wire n_7808;
wire n_11171;
wire n_6500;
wire n_4270;
wire n_8135;
wire n_9214;
wire n_13299;
wire n_7051;
wire n_9859;
wire n_11030;
wire n_13394;
wire n_10295;
wire n_5152;
wire n_9003;
wire n_11443;
wire n_9271;
wire n_9258;
wire n_3680;
wire n_6628;
wire n_13849;
wire n_12661;
wire n_12693;
wire n_6297;
wire n_5905;
wire n_12203;
wire n_6975;
wire n_5409;
wire n_6329;
wire n_7536;
wire n_8979;
wire n_12080;
wire n_8529;
wire n_10658;
wire n_5688;
wire n_9763;
wire n_5128;
wire n_10894;
wire n_4566;
wire n_9597;
wire n_6293;
wire n_8417;
wire n_9965;
wire n_9076;
wire n_10912;
wire n_7952;
wire n_4576;
wire n_9393;
wire n_8498;
wire n_7991;
wire n_7676;
wire n_11769;
wire n_4061;
wire n_12486;
wire n_7553;
wire n_6905;
wire n_12623;
wire n_7425;
wire n_13698;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_14701;
wire n_5307;
wire n_12933;
wire n_12489;
wire n_8967;
wire n_8355;
wire n_9736;
wire n_4767;
wire n_13691;
wire n_7998;
wire n_14122;
wire n_4328;
wire n_5986;
wire n_8719;
wire n_6581;
wire n_10160;
wire n_10678;
wire n_14372;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_11794;
wire n_14645;
wire n_5415;
wire n_4676;
wire n_10241;
wire n_5770;
wire n_11495;
wire n_14259;
wire n_7064;
wire n_5892;
wire n_8762;
wire n_12480;
wire n_13265;
wire n_4544;
wire n_13273;
wire n_10180;
wire n_8516;
wire n_8880;
wire n_6577;
wire n_6899;
wire n_8784;
wire n_14666;
wire n_12335;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_10631;
wire n_8237;
wire n_5802;
wire n_13372;
wire n_10852;
wire n_14546;
wire n_13669;
wire n_9803;
wire n_4429;
wire n_8977;
wire n_13079;
wire n_14371;
wire n_11406;
wire n_8171;
wire n_13121;
wire n_4591;
wire n_10978;
wire n_10500;
wire n_6370;
wire n_9755;
wire n_9805;
wire n_13731;
wire n_7210;
wire n_14997;
wire n_4646;
wire n_7899;
wire n_10370;
wire n_9728;
wire n_5769;
wire n_6065;
wire n_13845;
wire n_7039;
wire n_9659;
wire n_6987;
wire n_12624;
wire n_14328;
wire n_4563;
wire n_4725;
wire n_9107;
wire n_11428;
wire n_14361;
wire n_4169;
wire n_6859;
wire n_5331;
wire n_6190;
wire n_14311;
wire n_13447;
wire n_12410;
wire n_9917;
wire n_14574;
wire n_14847;
wire n_6309;
wire n_11149;
wire n_9520;
wire n_6623;
wire n_12055;
wire n_12925;
wire n_7723;
wire n_12771;
wire n_6527;
wire n_7443;
wire n_13262;
wire n_11707;
wire n_10550;
wire n_9583;
wire n_7811;
wire n_12413;
wire n_11086;
wire n_5341;
wire n_4320;
wire n_12182;
wire n_14096;
wire n_14943;
wire n_5930;
wire n_13622;
wire n_5814;
wire n_12803;
wire n_4881;
wire n_9036;
wire n_14007;
wire n_15026;
wire n_9522;
wire n_13145;
wire n_5979;
wire n_14034;
wire n_5271;
wire n_5089;
wire n_10571;
wire n_7015;
wire n_5263;
wire n_13276;
wire n_14394;
wire n_11772;
wire n_13338;
wire n_14618;
wire n_12547;
wire n_11764;
wire n_6929;
wire n_11225;
wire n_13904;
wire n_14256;
wire n_12544;
wire n_11339;
wire n_4012;
wire n_5518;
wire n_10125;
wire n_5637;
wire n_4636;
wire n_12370;
wire n_4584;
wire n_12931;
wire n_14810;
wire n_8279;
wire n_5622;
wire n_13940;
wire n_14054;
wire n_13648;
wire n_14844;
wire n_3910;
wire n_4711;
wire n_11112;
wire n_9723;
wire n_12986;
wire n_13570;
wire n_7348;
wire n_10254;
wire n_5240;
wire n_5813;
wire n_13543;
wire n_5495;
wire n_4680;
wire n_5546;
wire n_8912;
wire n_13873;
wire n_14491;
wire n_9488;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_5224;
wire n_4191;
wire n_4293;
wire n_14267;
wire n_7155;
wire n_8227;
wire n_3688;
wire n_9231;
wire n_8938;
wire n_6865;
wire n_8787;
wire n_5393;
wire n_10017;
wire n_6535;
wire n_7213;
wire n_14987;
wire n_10866;
wire n_9047;
wire n_10348;
wire n_14846;
wire n_12991;
wire n_4671;
wire n_8270;
wire n_4209;
wire n_5966;
wire n_11072;
wire n_7456;
wire n_8335;
wire n_11359;
wire n_13459;
wire n_13449;
wire n_13781;
wire n_14974;
wire n_10657;
wire n_13899;
wire n_7420;
wire n_5041;
wire n_14223;
wire n_11605;
wire n_13395;
wire n_9798;
wire n_14463;
wire n_9681;
wire n_8054;
wire n_9414;
wire n_12419;
wire n_8607;
wire n_5431;
wire n_13760;
wire n_9979;
wire n_9093;
wire n_14151;
wire n_11959;
wire n_6482;
wire n_5026;
wire n_3863;
wire n_11318;
wire n_11830;
wire n_10842;
wire n_13012;
wire n_12865;
wire n_8150;
wire n_5059;
wire n_9379;
wire n_5505;
wire n_12009;
wire n_7715;
wire n_9486;
wire n_3732;
wire n_11881;
wire n_6605;
wire n_4250;
wire n_9134;
wire n_5329;
wire n_12481;
wire n_4699;
wire n_7007;
wire n_8358;
wire n_9410;
wire n_3906;
wire n_4127;
wire n_10045;
wire n_14672;
wire n_13594;
wire n_13991;
wire n_7909;
wire n_14751;
wire n_14307;
wire n_9151;
wire n_12278;
wire n_13102;
wire n_4292;
wire n_14407;
wire n_3641;
wire n_4577;
wire n_11863;
wire n_14715;
wire n_14563;
wire n_13558;
wire n_4854;
wire n_14428;
wire n_8281;
wire n_12562;
wire n_11494;
wire n_9182;
wire n_5908;
wire n_6018;
wire n_12744;
wire n_4202;
wire n_7168;
wire n_11850;
wire n_5212;
wire n_9976;
wire n_7736;
wire n_5000;
wire n_14107;
wire n_8396;
wire n_9591;
wire n_10322;
wire n_13952;
wire n_9838;
wire n_7177;
wire n_5939;
wire n_10033;
wire n_3766;
wire n_12615;
wire n_13027;
wire n_14478;
wire n_11258;
wire n_10886;
wire n_9568;
wire n_7780;
wire n_9701;
wire n_9261;
wire n_7379;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_11468;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_7813;
wire n_7030;
wire n_8459;
wire n_5420;
wire n_6311;
wire n_11192;
wire n_12580;
wire n_11569;
wire n_4412;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_9752;
wire n_12769;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_12540;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_3815;
wire n_6029;
wire n_13607;
wire n_13080;
wire n_8379;
wire n_11563;
wire n_15089;
wire n_6879;
wire n_13292;
wire n_5259;
wire n_5440;
wire n_5679;
wire n_5938;
wire n_3710;
wire n_9079;
wire n_6702;
wire n_4155;
wire n_11846;
wire n_3891;
wire n_5891;
wire n_14682;
wire n_10383;
wire n_13377;
wire n_4144;
wire n_5724;
wire n_10064;
wire n_10876;
wire n_5774;
wire n_8793;
wire n_11852;
wire n_6452;
wire n_4374;
wire n_12619;
wire n_8975;
wire n_14527;
wire n_14020;
wire n_6791;
wire n_9170;
wire n_11679;
wire n_8792;
wire n_5131;
wire n_7280;
wire n_8671;
wire n_8489;
wire n_7110;
wire n_6915;
wire n_7511;
wire n_10831;
wire n_6856;
wire n_7941;
wire n_7791;
wire n_9385;
wire n_11186;
wire n_11870;
wire n_12960;
wire n_13519;
wire n_8484;
wire n_3834;
wire n_8454;
wire n_11492;
wire n_13984;
wire n_10536;
wire n_10238;
wire n_7232;
wire n_8759;
wire n_12268;
wire n_11544;
wire n_7345;
wire n_4548;
wire n_5923;
wire n_8703;
wire n_11233;
wire n_12656;
wire n_5790;
wire n_12678;
wire n_14521;
wire n_10206;
wire n_14726;
wire n_4989;
wire n_14924;
wire n_4622;
wire n_4315;
wire n_12880;
wire n_9670;
wire n_12876;
wire n_6451;
wire n_6364;
wire n_13107;
wire n_12711;
wire n_13511;
wire n_6552;
wire n_14205;
wire n_10786;
wire n_8325;
wire n_13523;
wire n_5140;
wire n_6328;
wire n_9598;
wire n_4816;
wire n_8382;
wire n_7827;
wire n_8971;
wire n_6363;
wire n_11646;
wire n_10602;
wire n_10620;
wire n_13699;
wire n_14049;
wire n_13420;
wire n_7159;
wire n_8127;
wire n_11878;
wire n_10079;
wire n_10188;
wire n_3810;
wire n_8721;
wire n_9391;
wire n_12458;
wire n_6132;
wire n_6578;
wire n_8889;
wire n_6406;
wire n_10319;
wire n_5598;
wire n_13643;
wire n_13603;
wire n_11900;
wire n_9470;
wire n_12132;
wire n_14434;
wire n_5306;
wire n_6978;
wire n_12104;
wire n_12037;
wire n_9328;
wire n_12467;
wire n_4483;
wire n_12870;
wire n_5342;
wire n_9245;
wire n_10739;
wire n_12911;
wire n_8232;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_12386;
wire n_7363;
wire n_4793;
wire n_9833;
wire n_11837;
wire n_10213;
wire n_6612;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_4168;
wire n_10872;
wire n_5997;
wire n_9455;
wire n_12651;
wire n_5511;
wire n_7863;
wire n_9719;
wire n_5680;
wire n_4806;
wire n_4350;
wire n_7295;
wire n_8633;
wire n_9744;
wire n_8842;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_11871;
wire n_8956;
wire n_5280;
wire n_10969;
wire n_6375;
wire n_6479;
wire n_14507;
wire n_6866;
wire n_12563;
wire n_7831;
wire n_13825;
wire n_11674;
wire n_12621;
wire n_5235;
wire n_3836;
wire n_13798;
wire n_3963;
wire n_14564;
wire n_12331;
wire n_12304;
wire n_9698;
wire n_12339;
wire n_6170;
wire n_12270;
wire n_14599;
wire n_15049;
wire n_9124;
wire n_10669;
wire n_10718;
wire n_9695;
wire n_4187;
wire n_6447;
wire n_4166;
wire n_6263;
wire n_7093;
wire n_9497;
wire n_5206;
wire n_10895;
wire n_8641;
wire n_8479;
wire n_11610;
wire n_11187;
wire n_12210;
wire n_7466;
wire n_14525;
wire n_14058;
wire n_5419;
wire n_6130;
wire n_12858;
wire n_14153;
wire n_15101;
wire n_12382;
wire n_11280;
wire n_10757;
wire n_7651;
wire n_4937;
wire n_3980;
wire n_13324;
wire n_10513;
wire n_15018;
wire n_5103;
wire n_3755;
wire n_11148;
wire n_8179;
wire n_5803;
wire n_13286;
wire n_4258;
wire n_14272;
wire n_6014;
wire n_4498;
wire n_11396;
wire n_8973;
wire n_6935;
wire n_14953;
wire n_10194;
wire n_9775;
wire n_7530;
wire n_5285;
wire n_11426;
wire n_4064;
wire n_14980;
wire n_9038;
wire n_8308;
wire n_4936;
wire n_13406;
wire n_5387;
wire n_9630;
wire n_13071;
wire n_10692;
wire n_8378;
wire n_3841;
wire n_8733;
wire n_12107;
wire n_8809;
wire n_14337;
wire n_4770;
wire n_5985;
wire n_14439;
wire n_11723;
wire n_11009;
wire n_4907;
wire n_9652;
wire n_10021;
wire n_5058;
wire n_12381;
wire n_6907;
wire n_11706;
wire n_13284;
wire n_8500;
wire n_12653;
wire n_6158;
wire n_7661;
wire n_10782;
wire n_9709;
wire n_6541;
wire n_6119;
wire n_8447;
wire n_14202;
wire n_5018;
wire n_11949;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_13303;
wire n_15004;
wire n_10457;
wire n_9324;
wire n_13311;
wire n_3690;
wire n_9934;
wire n_13364;
wire n_13813;
wire n_11957;
wire n_5192;
wire n_8548;
wire n_11538;
wire n_5141;
wire n_14743;
wire n_3716;
wire n_5133;
wire n_8412;
wire n_6226;
wire n_4712;
wire n_11264;
wire n_3837;
wire n_11211;
wire n_12774;
wire n_11880;
wire n_9668;
wire n_14340;
wire n_7145;
wire n_10385;
wire n_11377;
wire n_12064;
wire n_9877;
wire n_4310;
wire n_12503;
wire n_9657;
wire n_10111;
wire n_11302;
wire n_6338;
wire n_12425;
wire n_14319;
wire n_14922;
wire n_11921;
wire n_13358;
wire n_5159;
wire n_9352;
wire n_3954;
wire n_9395;
wire n_12807;
wire n_14621;
wire n_8425;
wire n_10809;
wire n_9349;
wire n_4674;
wire n_4908;
wire n_14734;
wire n_8241;
wire n_7823;
wire n_9209;
wire n_7467;
wire n_5097;
wire n_14555;
wire n_10113;
wire n_15010;
wire n_11267;
wire n_10990;
wire n_7932;
wire n_11626;
wire n_14957;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_11694;
wire n_13811;
wire n_14014;
wire n_4159;
wire n_3714;
wire n_11618;
wire n_9969;
wire n_3739;
wire n_9937;
wire n_5816;
wire n_4069;
wire n_7541;
wire n_3718;
wire n_10545;
wire n_12715;
wire n_4862;
wire n_7241;
wire n_7717;
wire n_14945;
wire n_5300;
wire n_10595;
wire n_10973;
wire n_13883;
wire n_11011;
wire n_13814;
wire n_12015;
wire n_12968;
wire n_9618;
wire n_10732;
wire n_14257;
wire n_10009;
wire n_11776;
wire n_6625;
wire n_4850;
wire n_11165;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_12135;
wire n_7464;
wire n_9082;
wire n_11366;
wire n_6302;
wire n_14279;
wire n_9424;
wire n_8274;
wire n_9453;
wire n_5748;
wire n_13757;
wire n_6759;
wire n_5525;
wire n_9637;
wire n_8152;
wire n_6706;
wire n_10526;
wire n_8550;
wire n_3889;
wire n_6139;
wire n_14190;
wire n_4256;
wire n_14185;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_6999;
wire n_7054;
wire n_12817;
wire n_13832;
wire n_4224;
wire n_6403;
wire n_6483;
wire n_8829;
wire n_9183;
wire n_9205;
wire n_14630;
wire n_13935;
wire n_12869;
wire n_9009;
wire n_13325;
wire n_4024;
wire n_13841;
wire n_6228;
wire n_11315;
wire n_5650;
wire n_14104;
wire n_10044;
wire n_14344;
wire n_13207;
wire n_12059;
wire n_14188;
wire n_11098;
wire n_12586;
wire n_5400;
wire n_13043;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_10221;
wire n_4702;
wire n_13281;
wire n_6888;
wire n_8266;
wire n_13960;
wire n_15086;
wire n_14069;
wire n_8515;
wire n_10109;
wire n_10169;
wire n_4252;
wire n_13556;
wire n_4457;
wire n_8648;
wire n_6063;
wire n_10329;
wire n_10928;
wire n_9030;
wire n_9024;
wire n_9523;
wire n_9377;
wire n_10891;
wire n_8946;
wire n_15099;
wire n_10839;
wire n_11875;
wire n_6800;
wire n_5139;
wire n_13260;
wire n_9716;
wire n_6922;
wire n_9380;
wire n_14543;
wire n_5481;
wire n_6890;
wire n_14474;
wire n_8744;
wire n_9000;
wire n_9679;
wire n_9116;
wire n_9742;
wire n_9016;
wire n_7503;
wire n_6070;
wire n_13979;
wire n_13308;
wire n_9006;
wire n_12514;
wire n_13381;
wire n_11524;
wire n_10091;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7296;
wire n_6647;
wire n_7273;
wire n_5733;
wire n_14704;
wire n_10029;
wire n_9690;
wire n_8765;
wire n_4132;
wire n_13483;
wire n_14675;
wire n_5871;
wire n_9852;
wire n_7543;
wire n_4261;
wire n_13400;
wire n_10600;
wire n_9914;
wire n_11056;
wire n_11514;
wire n_12438;
wire n_6184;
wire n_14268;
wire n_4886;
wire n_11774;
wire n_8627;
wire n_4090;
wire n_7507;
wire n_9451;
wire n_10849;
wire n_5043;
wire n_11108;
wire n_9760;
wire n_7555;
wire n_13910;
wire n_5707;
wire n_13907;
wire n_10947;
wire n_4001;
wire n_13369;
wire n_10272;
wire n_12099;
wire n_9035;
wire n_15077;
wire n_12806;
wire n_4371;
wire n_5836;
wire n_9211;
wire n_5281;
wire n_14873;
wire n_6716;
wire n_6422;
wire n_12887;
wire n_12776;
wire n_4473;
wire n_4007;
wire n_12898;
wire n_4268;
wire n_9677;
wire n_13464;
wire n_5048;
wire n_11954;
wire n_14965;
wire n_5521;
wire n_12191;
wire n_7578;
wire n_5028;
wire n_13611;
wire n_4480;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_8195;
wire n_9070;
wire n_5585;
wire n_6397;
wire n_12578;
wire n_4824;
wire n_4120;
wire n_14012;
wire n_4427;
wire n_11864;
wire n_3745;
wire n_14221;
wire n_14232;
wire n_7033;
wire n_9881;
wire n_6121;
wire n_9669;
wire n_7531;
wire n_4142;
wire n_9958;
wire n_4082;
wire n_9858;
wire n_8462;
wire n_5561;
wire n_9981;
wire n_4085;
wire n_10391;
wire n_4073;
wire n_4260;
wire n_8377;
wire n_11157;
wire n_14390;
wire n_4163;
wire n_4439;
wire n_12509;
wire n_13345;
wire n_12235;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_14932;
wire n_9588;
wire n_6954;
wire n_11733;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_12471;
wire n_13632;
wire n_13756;
wire n_12365;
wire n_5875;
wire n_8428;
wire n_8103;
wire n_13417;
wire n_4262;
wire n_14350;
wire n_9021;
wire n_13130;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_8362;
wire n_12083;
wire n_9682;
wire n_10137;
wire n_10344;
wire n_7131;
wire n_4720;
wire n_7769;
wire n_10882;
wire n_11540;
wire n_11861;
wire n_6903;
wire n_9050;
wire n_11724;
wire n_9303;
wire n_14775;
wire n_12065;
wire n_9495;
wire n_13970;
wire n_12167;
wire n_11220;
wire n_14220;
wire n_4685;
wire n_6101;
wire n_9415;
wire n_5968;
wire n_14451;
wire n_10196;
wire n_8491;
wire n_9058;
wire n_4334;
wire n_6941;
wire n_9845;
wire n_8831;
wire n_4511;
wire n_5812;
wire n_14100;
wire n_6148;
wire n_5515;
wire n_8324;
wire n_11459;
wire n_11355;
wire n_6106;
wire n_9822;
wire n_12087;
wire n_6604;
wire n_14510;
wire n_12243;
wire n_4014;
wire n_7418;
wire n_12267;
wire n_5250;
wire n_12569;
wire n_4757;
wire n_7688;
wire n_10518;
wire n_11101;
wire n_9640;
wire n_11899;
wire n_8348;
wire n_5607;
wire n_14313;
wire n_4175;
wire n_8288;
wire n_10613;
wire n_10583;
wire n_14719;
wire n_4648;
wire n_14452;
wire n_11481;
wire n_14308;
wire n_11712;
wire n_11612;
wire n_8269;
wire n_5006;
wire n_14288;
wire n_7806;
wire n_10335;
wire n_10085;
wire n_10840;
wire n_6566;
wire n_14833;
wire n_13152;
wire n_12599;
wire n_8625;
wire n_5734;
wire n_6081;
wire n_8458;
wire n_4892;
wire n_8806;
wire n_13857;
wire n_7204;
wire n_10560;
wire n_3823;
wire n_8180;
wire n_4173;
wire n_8601;
wire n_8499;
wire n_4970;
wire n_9062;
wire n_3816;
wire n_13315;
wire n_14606;
wire n_13180;
wire n_14097;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_8306;
wire n_12513;
wire n_12091;
wire n_9722;
wire n_12375;
wire n_6047;
wire n_14788;
wire n_8167;
wire n_5438;
wire n_10486;
wire n_9791;
wire n_12307;
wire n_9229;
wire n_11603;
wire n_11890;
wire n_4627;
wire n_8613;
wire n_9603;
wire n_11790;
wire n_8913;
wire n_11060;
wire n_7354;
wire n_7448;
wire n_8800;
wire n_6244;
wire n_13474;
wire n_13224;
wire n_12684;
wire n_8768;
wire n_6861;
wire n_13702;
wire n_9099;
wire n_3783;
wire n_10919;
wire n_13797;
wire n_3843;
wire n_14388;
wire n_12288;
wire n_9309;
wire n_12418;
wire n_13853;
wire n_7852;
wire n_13762;
wire n_10952;
wire n_5725;
wire n_12566;
wire n_7925;
wire n_12415;
wire n_13037;
wire n_9432;
wire n_9454;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_11744;
wire n_13919;
wire n_14466;
wire n_9065;
wire n_11650;
wire n_5163;
wire n_11518;
wire n_7748;
wire n_5768;
wire n_12949;
wire n_4961;
wire n_7556;
wire n_14061;
wire n_3753;
wire n_7640;
wire n_8187;
wire n_10352;
wire n_14962;
wire n_8881;
wire n_9704;
wire n_4718;
wire n_11663;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_9837;
wire n_10991;
wire n_4317;
wire n_4855;
wire n_9431;
wire n_10167;
wire n_3969;
wire n_12681;
wire n_12859;
wire n_14413;
wire n_9160;
wire n_10911;
wire n_4154;
wire n_9433;
wire n_14050;
wire n_6588;
wire n_9256;
wire n_10442;
wire n_12829;
wire n_13593;
wire n_11282;
wire n_14912;
wire n_9706;
wire n_12448;
wire n_13044;
wire n_7900;
wire n_7050;
wire n_4023;
wire n_9808;
wire n_9915;
wire n_13723;
wire n_10534;
wire n_14156;
wire n_5685;
wire n_4420;
wire n_11726;
wire n_13188;
wire n_5773;
wire n_7136;
wire n_10465;
wire n_10406;
wire n_12188;
wire n_12943;
wire n_8316;
wire n_7318;
wire n_13923;
wire n_12149;
wire n_6055;
wire n_5138;
wire n_12783;
wire n_8397;
wire n_9184;
wire n_5374;
wire n_10373;
wire n_13472;
wire n_9133;
wire n_6108;
wire n_8115;
wire n_12129;
wire n_12631;
wire n_6165;
wire n_14387;
wire n_10965;
wire n_6621;
wire n_13148;
wire n_7175;
wire n_5349;
wire n_4973;
wire n_7810;
wire n_9109;
wire n_4640;
wire n_13964;
wire n_6323;
wire n_10517;
wire n_12588;
wire n_12652;
wire n_8523;
wire n_9207;
wire n_11458;
wire n_4396;
wire n_13485;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_13531;
wire n_13355;
wire n_13368;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_13160;
wire n_10484;
wire n_5766;
wire n_11255;
wire n_5216;
wire n_6597;
wire n_13676;
wire n_10561;
wire n_13183;
wire n_9673;
wire n_13601;
wire n_8891;
wire n_12523;
wire n_7817;
wire n_3818;
wire n_8294;
wire n_11856;
wire n_14312;
wire n_6933;
wire n_4387;
wire n_7878;
wire n_8338;
wire n_4951;
wire n_12579;
wire n_9010;
wire n_14904;
wire n_8915;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_11442;
wire n_13052;
wire n_7289;
wire n_14754;
wire n_5805;
wire n_7665;
wire n_8131;
wire n_11747;
wire n_9552;
wire n_3719;
wire n_7855;
wire n_11008;
wire n_10371;
wire n_3681;
wire n_11243;
wire n_9841;
wire n_12675;
wire n_13006;
wire n_9230;
wire n_12174;
wire n_14947;
wire n_14659;
wire n_7764;
wire n_4308;
wire n_12113;
wire n_12831;
wire n_10198;
wire n_8027;
wire n_6216;
wire n_10096;
wire n_3830;
wire n_10582;
wire n_11425;
wire n_10638;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_9132;
wire n_11992;
wire n_6949;
wire n_6509;
wire n_14198;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_8855;
wire n_10483;
wire n_11657;
wire n_4152;
wire n_13820;
wire n_12470;
wire n_14039;
wire n_8546;
wire n_9878;
wire n_11536;
wire n_11717;
wire n_9069;
wire n_8966;
wire n_12154;
wire n_8487;
wire n_7263;
wire n_8844;
wire n_14995;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_5611;
wire n_10662;
wire n_13471;
wire n_6911;
wire n_9674;
wire n_11512;
wire n_11327;
wire n_8533;
wire n_4281;
wire n_4661;
wire n_12799;
wire n_4200;
wire n_13114;
wire n_15002;
wire n_8869;
wire n_5900;
wire n_4962;
wire n_14956;
wire n_9786;
wire n_13976;
wire n_6327;
wire n_8584;
wire n_13200;
wire n_11140;
wire n_8932;
wire n_14862;
wire n_9063;
wire n_8998;
wire n_6607;
wire n_9188;
wire n_9467;
wire n_9372;
wire n_10960;
wire n_11078;
wire n_4958;
wire n_9743;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_11620;
wire n_7209;
wire n_5171;
wire n_12617;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_12919;
wire n_8480;
wire n_9926;
wire n_7240;
wire n_10094;
wire n_12095;
wire n_14620;
wire n_10749;
wire n_11907;
wire n_4071;
wire n_14291;
wire n_4921;
wire n_14092;
wire n_12432;
wire n_12796;
wire n_8911;
wire n_11352;
wire n_5427;
wire n_5639;
wire n_14293;
wire n_7725;
wire n_8398;
wire n_4361;
wire n_10585;
wire n_15039;
wire n_5417;
wire n_8772;
wire n_12008;
wire n_4614;
wire n_12279;
wire n_9480;
wire n_8307;
wire n_14005;
wire n_14884;
wire n_10896;
wire n_8767;
wire n_9113;
wire n_13764;
wire n_9158;
wire n_12156;
wire n_11851;
wire n_4945;
wire n_14441;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_14688;
wire n_13264;
wire n_8010;
wire n_7278;
wire n_11986;
wire n_12637;
wire n_12301;
wire n_9263;
wire n_8347;
wire n_11734;
wire n_7630;
wire n_11517;
wire n_11022;
wire n_14468;
wire n_11831;
wire n_10162;
wire n_12302;
wire n_14766;
wire n_8466;
wire n_6416;
wire n_5488;
wire n_4693;
wire n_12190;
wire n_14222;
wire n_15054;
wire n_9632;
wire n_10353;
wire n_8813;
wire n_8354;
wire n_4326;
wire n_6695;
wire n_8204;
wire n_14067;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_14598;
wire n_6127;
wire n_7565;
wire n_11259;
wire n_14446;
wire n_11197;
wire n_9282;
wire n_4305;
wire n_14747;
wire n_14909;
wire n_5781;
wire n_7883;
wire n_6600;
wire n_10933;
wire n_14046;
wire n_12192;
wire n_7410;
wire n_12010;
wire n_12977;
wire n_4213;
wire n_10546;
wire n_7097;
wire n_12864;
wire n_3692;
wire n_13227;
wire n_13869;
wire n_9503;
wire n_6421;
wire n_10724;
wire n_5747;
wire n_7414;
wire n_11427;
wire n_10660;
wire n_13348;
wire n_13166;
wire n_7495;
wire n_9782;
wire n_5969;
wire n_13350;
wire n_9114;
wire n_8312;
wire n_9855;
wire n_4929;
wire n_8040;
wire n_14242;
wire n_11153;
wire n_9347;
wire n_4964;
wire n_13615;
wire n_9469;
wire n_9746;
wire n_9680;
wire n_10923;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_9633;
wire n_12746;
wire n_10836;
wire n_13266;
wire n_6458;
wire n_10884;
wire n_4139;
wire n_13319;
wire n_13623;
wire n_15062;
wire n_8132;
wire n_6746;
wire n_12436;
wire n_4031;
wire n_7586;
wire n_10780;
wire n_9501;
wire n_12528;
wire n_7720;
wire n_6719;
wire n_13544;
wire n_12792;
wire n_14586;
wire n_5437;
wire n_9148;
wire n_13530;
wire n_11475;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_12973;
wire n_14095;
wire n_11385;
wire n_14191;
wire n_6506;
wire n_14289;
wire n_6287;
wire n_4583;
wire n_13092;
wire n_6662;
wire n_8650;
wire n_12923;
wire n_10870;
wire n_12916;
wire n_9585;
wire n_10267;
wire n_13888;
wire n_8974;
wire n_10379;
wire n_4210;
wire n_5245;
wire n_14561;
wire n_7189;
wire n_8688;
wire n_4666;
wire n_3751;
wire n_10821;
wire n_10740;
wire n_8983;
wire n_10558;
wire n_6851;
wire n_8116;
wire n_12144;
wire n_9338;
wire n_12716;
wire n_6687;
wire n_10297;
wire n_6884;
wire n_8356;
wire n_8013;
wire n_9075;
wire n_13981;
wire n_14614;
wire n_3698;
wire n_3927;
wire n_4540;
wire n_3961;
wire n_6780;
wire n_6513;
wire n_12463;
wire n_12524;
wire n_4891;
wire n_8519;
wire n_14484;
wire n_7841;
wire n_10497;
wire n_6619;
wire n_10354;
wire n_11456;
wire n_8193;
wire n_14536;
wire n_5603;
wire n_10888;
wire n_6804;
wire n_9370;
wire n_11647;
wire n_12392;
wire n_13205;
wire n_13421;
wire n_12173;
wire n_9409;
wire n_14140;
wire n_5716;
wire n_3993;
wire n_10138;
wire n_4940;
wire n_6516;
wire n_10358;
wire n_5208;
wire n_7490;
wire n_7792;
wire n_10578;
wire n_6924;
wire n_4590;
wire n_13745;
wire n_7492;
wire n_12168;
wire n_12349;
wire n_13349;
wire n_10948;
wire n_5606;
wire n_13730;
wire n_15087;
wire n_4830;
wire n_12665;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_11736;
wire n_14339;
wire n_14804;
wire n_4664;
wire n_9626;
wire n_14501;
wire n_3860;
wire n_8154;
wire n_15007;
wire n_12067;
wire n_5456;
wire n_12546;
wire n_7073;
wire n_13489;
wire n_14825;
wire n_11393;
wire n_10007;
wire n_5093;
wire n_10904;
wire n_10386;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_9961;
wire n_13488;
wire n_14718;
wire n_5727;
wire n_4906;
wire n_9098;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_11325;
wire n_14612;
wire n_9861;
wire n_6788;
wire n_13638;
wire n_14869;
wire n_4883;
wire n_11660;
wire n_4162;
wire n_10448;
wire n_3665;
wire n_14985;
wire n_5115;
wire n_12963;
wire n_14110;
wire n_6393;
wire n_9536;
wire n_8566;
wire n_12282;
wire n_8086;
wire n_14316;
wire n_12620;
wire n_8746;
wire n_11411;
wire n_6249;
wire n_14506;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_13268;
wire n_12431;
wire n_3800;
wire n_9593;
wire n_9017;
wire n_5407;
wire n_14595;
wire n_11281;
wire n_11841;
wire n_4608;
wire n_11658;
wire n_5232;
wire n_14765;
wire n_9703;
wire n_14215;
wire n_7271;
wire n_3991;
wire n_12830;
wire n_11025;
wire n_6572;
wire n_12213;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_11372;
wire n_4536;
wire n_10450;
wire n_13117;
wire n_13510;
wire n_12397;
wire n_14781;
wire n_14920;
wire n_13665;
wire n_5149;
wire n_5967;
wire n_7569;
wire n_5151;
wire n_7003;
wire n_9565;
wire n_7897;
wire n_4773;
wire n_14954;
wire n_7962;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_13179;
wire n_13429;
wire n_10320;
wire n_4611;
wire n_14835;
wire n_8113;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_4960;
wire n_10308;
wire n_14216;
wire n_8652;
wire n_3864;
wire n_13993;
wire n_4658;
wire n_5135;
wire n_7419;
wire n_15025;
wire n_11545;
wire n_12974;
wire n_14078;
wire n_13717;
wire n_5827;
wire n_11465;
wire n_9337;
wire n_5494;
wire n_4362;
wire n_14314;
wire n_4306;
wire n_6200;
wire n_11437;
wire n_10304;
wire n_11436;
wire n_7784;
wire n_13804;
wire n_4422;
wire n_10902;
wire n_8714;
wire n_6123;
wire n_10607;
wire n_6934;
wire n_7094;
wire n_7500;
wire n_11463;
wire n_14152;
wire n_10605;
wire n_11394;
wire n_6082;
wire n_10668;
wire n_8944;
wire n_12487;
wire n_13660;
wire n_13861;
wire n_9232;
wire n_12385;
wire n_9320;
wire n_10713;
wire n_4555;
wire n_11191;
wire n_14937;
wire n_9167;
wire n_10464;
wire n_5136;
wire n_7864;
wire n_5228;
wire n_14580;
wire n_10596;
wire n_14654;
wire n_10034;
wire n_11068;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_13081;
wire n_7790;
wire n_14249;
wire n_4215;
wire n_6952;
wire n_7062;
wire n_4280;
wire n_10875;
wire n_4047;
wire n_12735;
wire n_9526;
wire n_5471;
wire n_8107;
wire n_7642;
wire n_5434;
wire n_12475;
wire n_14300;
wire n_9077;
wire n_5941;
wire n_7045;
wire n_12646;
wire n_5879;
wire n_11277;
wire n_11665;
wire n_5558;
wire n_11061;
wire n_13777;
wire n_9692;
wire n_13444;
wire n_13800;
wire n_14022;
wire n_5350;
wire n_13267;
wire n_13959;
wire n_9141;
wire n_11483;
wire n_5338;
wire n_7238;
wire n_12733;
wire n_7126;
wire n_9745;
wire n_5669;
wire n_9787;
wire n_3854;
wire n_8674;
wire n_11073;
wire n_14105;
wire n_12944;
wire n_13362;
wire n_14637;
wire n_7931;
wire n_10309;
wire n_12061;
wire n_12265;
wire n_13190;
wire n_12380;
wire n_8482;
wire n_11462;
wire n_8992;
wire n_14703;
wire n_13032;
wire n_6979;
wire n_11224;
wire n_10024;
wire n_9892;
wire n_6203;
wire n_7405;
wire n_10762;
wire n_7739;
wire n_13790;
wire n_10490;
wire n_14357;
wire n_8761;
wire n_7207;
wire n_9078;
wire n_8899;
wire n_11127;
wire n_4027;
wire n_7934;
wire n_9015;
wire n_7454;
wire n_14283;
wire n_9012;
wire n_4599;
wire n_12794;
wire n_5830;
wire n_6796;
wire n_4812;
wire n_9233;
wire n_12890;
wire n_14492;
wire n_9217;
wire n_13576;
wire n_14644;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_4628;
wire n_11632;
wire n_10974;
wire n_9435;
wire n_5668;
wire n_5878;
wire n_4873;
wire n_8926;
wire n_5588;
wire n_4657;
wire n_11692;
wire n_11762;
wire n_14662;
wire n_5765;
wire n_11843;
wire n_14341;
wire n_14470;
wire n_3950;
wire n_9389;
wire n_11344;
wire n_4458;
wire n_11403;
wire n_6596;
wire n_12926;
wire n_4121;
wire n_5090;
wire n_14159;
wire n_6870;
wire n_10520;
wire n_7639;
wire n_13666;
wire n_12247;
wire n_12881;
wire n_5613;
wire n_4476;
wire n_10914;
wire n_10129;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_13710;
wire n_11510;
wire n_10084;
wire n_14082;
wire n_7251;
wire n_10519;
wire n_7776;
wire n_12966;
wire n_6080;
wire n_10318;
wire n_13785;
wire n_7059;
wire n_13287;
wire n_14665;
wire n_8561;
wire n_10877;
wire n_8255;
wire n_7035;
wire n_10468;
wire n_14752;
wire n_5571;
wire n_11854;
wire n_12894;
wire n_8029;
wire n_10906;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_14632;
wire n_5513;
wire n_6747;
wire n_12276;
wire n_6281;
wire n_13588;
wire n_4803;
wire n_5972;
wire n_10289;
wire n_14496;
wire n_9381;
wire n_4079;
wire n_13261;
wire n_4091;
wire n_13634;
wire n_9873;
wire n_11925;
wire n_12594;
wire n_10905;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_13030;
wire n_14043;
wire n_9575;
wire n_5145;
wire n_12529;
wire n_14636;
wire n_11817;
wire n_3712;
wire n_6094;
wire n_15036;
wire n_6444;
wire n_11961;
wire n_12001;
wire n_5132;
wire n_5191;
wire n_10298;
wire n_12433;
wire n_6333;
wire n_10940;
wire n_6262;
wire n_12765;
wire n_13704;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_9023;
wire n_12097;
wire n_6240;
wire n_10723;
wire n_5359;
wire n_13627;
wire n_6412;
wire n_9412;
wire n_5293;
wire n_7782;
wire n_7220;
wire n_10293;
wire n_11824;
wire n_4316;
wire n_3697;
wire n_10361;
wire n_7438;
wire n_11269;
wire n_11270;
wire n_9955;
wire n_10161;
wire n_10432;
wire n_7515;
wire n_11532;
wire n_7574;
wire n_12402;
wire n_4044;
wire n_12728;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_8921;
wire n_3971;
wire n_13191;
wire n_13784;
wire n_13766;
wire n_10640;
wire n_11546;
wire n_7065;
wire n_10271;
wire n_11314;
wire n_5510;
wire n_6046;
wire n_7894;
wire n_9418;
wire n_7868;
wire n_6973;
wire n_9733;
wire n_14963;
wire n_5363;
wire n_7285;
wire n_8286;
wire n_5200;
wire n_9502;
wire n_5659;
wire n_5618;
wire n_15045;
wire n_6325;
wire n_13374;
wire n_9765;
wire n_9029;
wire n_11130;
wire n_10163;
wire n_13824;
wire n_6737;
wire n_12262;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_8178;
wire n_14175;
wire n_5369;
wire n_11935;
wire n_13452;
wire n_5258;
wire n_12708;
wire n_5255;
wire n_14423;
wire n_13656;
wire n_10576;
wire n_9623;
wire n_11822;
wire n_10424;
wire n_12805;
wire n_7008;
wire n_11035;
wire n_8925;
wire n_10404;
wire n_14138;
wire n_8432;
wire n_6111;
wire n_10130;
wire n_12901;
wire n_7505;
wire n_3758;
wire n_8047;
wire n_6260;
wire n_7501;
wire n_10214;
wire n_12971;
wire n_5080;
wire n_11389;
wire n_6665;
wire n_9783;
wire n_7566;
wire n_7937;
wire n_12658;
wire n_7055;
wire n_14568;
wire n_14562;
wire n_12372;
wire n_8268;
wire n_11501;
wire n_12564;
wire n_8053;
wire n_13141;
wire n_11015;
wire n_5858;
wire n_5817;
wire n_10317;
wire n_6690;
wire n_9840;
wire n_5723;
wire n_10491;
wire n_5295;
wire n_6137;
wire n_10712;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_9909;
wire n_10192;
wire n_7113;
wire n_12204;
wire n_14684;
wire n_4998;
wire n_15055;
wire n_10453;
wire n_11034;
wire n_8735;
wire n_11895;
wire n_7872;
wire n_12543;
wire n_13895;
wire n_10219;
wire n_5627;
wire n_12888;
wire n_13854;
wire n_4167;
wire n_14062;
wire n_8845;
wire n_7242;
wire n_5155;
wire n_14467;
wire n_3835;
wire n_6461;
wire n_8830;
wire n_12013;
wire n_11662;
wire n_3967;
wire n_5016;
wire n_14706;
wire n_7954;
wire n_6212;
wire n_6908;
wire n_7819;
wire n_6570;
wire n_14362;
wire n_12741;
wire n_8022;
wire n_9532;
wire n_8415;
wire n_9112;
wire n_6498;
wire n_3902;
wire n_10062;
wire n_4730;
wire n_7228;
wire n_9561;
wire n_6692;
wire n_8547;
wire n_14553;
wire n_10788;
wire n_11500;
wire n_15092;
wire n_6074;
wire n_10910;
wire n_7561;
wire n_6380;
wire n_3654;
wire n_10892;
wire n_10216;
wire n_9091;
wire n_14377;
wire n_5996;
wire n_8386;
wire n_8426;
wire n_9326;
wire n_8672;
wire n_11977;
wire n_10049;
wire n_5327;
wire n_7994;
wire n_9180;
wire n_10431;
wire n_11215;
wire n_8540;
wire n_6045;
wire n_9932;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_13705;
wire n_14535;
wire n_14776;
wire n_9220;
wire n_9834;
wire n_7415;
wire n_13726;
wire n_9474;
wire n_14770;
wire n_14551;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_9542;
wire n_11530;
wire n_7598;
wire n_14406;
wire n_15001;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_15000;
wire n_14449;
wire n_12889;
wire n_14290;
wire n_8192;
wire n_14919;
wire n_5791;
wire n_8791;
wire n_9458;
wire n_10608;
wire n_4204;
wire n_9642;
wire n_14768;
wire n_5098;
wire n_6772;
wire n_6877;
wire n_9020;
wire n_6823;
wire n_9910;
wire n_6806;
wire n_7426;
wire n_11014;
wire n_5906;
wire n_8350;
wire n_11439;
wire n_14744;
wire n_12526;
wire n_9100;
wire n_11119;
wire n_11752;
wire n_14081;
wire n_14410;
wire n_4743;
wire n_8816;
wire n_3805;
wire n_7957;
wire n_3825;
wire n_8712;
wire n_14549;
wire n_8048;
wire n_6831;
wire n_15058;
wire n_3657;
wire n_10395;
wire n_4924;
wire n_3928;
wire n_12255;
wire n_9781;
wire n_13881;
wire n_8663;
wire n_4859;
wire n_7217;
wire n_9940;
wire n_12068;
wire n_10802;
wire n_6284;
wire n_7058;
wire n_6157;
wire n_4654;
wire n_5423;
wire n_7497;
wire n_8503;
wire n_6785;
wire n_8254;
wire n_6374;
wire n_8959;
wire n_13280;
wire n_9117;
wire n_6930;
wire n_12784;
wire n_9198;
wire n_6017;
wire n_3792;
wire n_4733;
wire n_11729;
wire n_8506;
wire n_4272;
wire n_11289;
wire n_3974;
wire n_3871;
wire n_11699;
wire n_7735;
wire n_8265;
wire n_8465;
wire n_8049;
wire n_12277;
wire n_4269;
wire n_4695;
wire n_6838;
wire n_11902;
wire n_12212;
wire n_12126;
wire n_5736;
wire n_6937;
wire n_12686;
wire n_6443;
wire n_6105;
wire n_13328;
wire n_10080;
wire n_7558;
wire n_13554;
wire n_12344;
wire n_12250;
wire n_8937;
wire n_12961;
wire n_14142;
wire n_5069;
wire n_7442;
wire n_10574;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_9249;
wire n_11628;
wire n_10594;
wire n_11784;
wire n_12193;
wire n_3968;
wire n_9398;
wire n_5099;
wire n_11622;
wire n_14033;
wire n_4704;
wire n_14269;
wire n_4551;
wire n_11763;
wire n_13393;
wire n_5052;
wire n_6091;
wire n_11606;
wire n_12749;
wire n_6674;
wire n_4957;
wire n_10155;
wire n_14585;
wire n_6034;
wire n_15032;
wire n_7499;
wire n_4072;
wire n_9751;
wire n_14866;
wire n_13134;
wire n_5579;
wire n_8381;
wire n_13399;
wire n_7085;
wire n_13413;
wire n_12079;
wire n_4781;
wire n_9579;
wire n_11006;
wire n_10879;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_6762;
wire n_15090;
wire n_7341;
wire n_7895;
wire n_13602;
wire n_4424;
wire n_11321;
wire n_13250;
wire n_8366;
wire n_10792;
wire n_8101;
wire n_7611;
wire n_9925;
wire n_10655;
wire n_14065;
wire n_7391;
wire n_14713;
wire n_3711;
wire n_10890;
wire n_12187;
wire n_12093;
wire n_5837;
wire n_14539;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_8384;
wire n_13035;
wire n_9889;
wire n_5642;
wire n_14299;
wire n_12705;
wire n_7224;
wire n_5880;
wire n_8728;
wire n_6169;
wire n_11133;
wire n_4746;
wire n_12241;
wire n_14114;
wire n_12211;
wire n_15082;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_15100;
wire n_10212;
wire n_8023;
wire n_13770;
wire n_13975;
wire n_8052;
wire n_11001;
wire n_7627;
wire n_9998;
wire n_11143;
wire n_10654;
wire n_9729;
wire n_5118;
wire n_5105;
wire n_14112;
wire n_3850;
wire n_13833;
wire n_13886;
wire n_4459;
wire n_11757;
wire n_13169;
wire n_8614;
wire n_5793;
wire n_5591;
wire n_13237;
wire n_7856;
wire n_4050;
wire n_9081;
wire n_7496;
wire n_12446;
wire n_12640;
wire n_12699;
wire n_9784;
wire n_13354;
wire n_13696;
wire n_5623;
wire n_12856;
wire n_14834;
wire n_10005;
wire n_10544;
wire n_10217;
wire n_12231;
wire n_5681;
wire n_4853;
wire n_11421;
wire n_11780;
wire n_12745;
wire n_14798;
wire n_9856;
wire n_9101;
wire n_7399;
wire n_12841;
wire n_6213;
wire n_8656;
wire n_10393;
wire n_6118;
wire n_5256;
wire n_11793;
wire n_12527;
wire n_7605;
wire n_14386;
wire n_11400;
wire n_5220;
wire n_12814;
wire n_5732;
wire n_8897;
wire n_3852;
wire n_9696;
wire n_12545;
wire n_5178;
wire n_11621;
wire n_6814;
wire n_4520;
wire n_13913;
wire n_7342;
wire n_12354;
wire n_4008;
wire n_8014;
wire n_9825;
wire n_13783;
wire n_5507;
wire n_10093;
wire n_8564;
wire n_11969;
wire n_14926;
wire n_7472;
wire n_7214;
wire n_12685;
wire n_5077;
wire n_10850;
wire n_12886;
wire n_13297;
wire n_8371;
wire n_10945;
wire n_5872;
wire n_13564;
wire n_14601;
wire n_11791;
wire n_7408;
wire n_3858;
wire n_8231;
wire n_9250;
wire n_6115;
wire n_4502;
wire n_9572;
wire n_10541;
wire n_6858;
wire n_12196;
wire n_10375;
wire n_11948;
wire n_11910;
wire n_8558;
wire n_4851;
wire n_5735;
wire n_12119;
wire n_9483;
wire n_10275;
wire n_9816;
wire n_9253;
wire n_15080;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_9136;
wire n_14280;
wire n_7837;
wire n_8357;
wire n_10726;
wire n_9426;
wire n_3924;
wire n_8870;
wire n_9831;
wire n_4571;
wire n_13434;
wire n_14017;
wire n_14395;
wire n_8143;
wire n_11064;
wire n_14187;
wire n_6430;
wire n_14027;
wire n_6193;
wire n_10614;
wire n_5314;
wire n_6462;
wire n_8422;
wire n_12094;
wire n_12096;
wire n_9896;
wire n_9650;
wire n_13657;
wire n_12730;
wire n_10002;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_14639;
wire n_4205;
wire n_5953;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_11974;
wire n_12202;
wire n_6779;
wire n_6518;
wire n_9767;
wire n_6797;
wire n_11367;
wire n_14094;
wire n_4454;
wire n_7938;
wire n_8253;
wire n_4229;
wire n_14730;
wire n_5952;
wire n_4739;
wire n_12534;
wire n_13692;
wire n_5820;
wire n_5483;
wire n_12120;
wire n_9028;
wire n_9055;
wire n_5718;
wire n_10251;
wire n_14722;
wire n_11562;
wire n_11866;
wire n_13585;
wire n_6916;
wire n_3904;
wire n_5150;
wire n_11383;
wire n_12854;
wire n_8563;
wire n_9949;
wire n_4838;
wire n_5075;
wire n_11655;
wire n_12553;
wire n_7812;
wire n_12816;
wire n_14906;
wire n_4879;
wire n_5051;
wire n_14486;
wire n_11552;
wire n_14807;
wire n_9684;
wire n_3926;
wire n_6152;
wire n_10010;
wire n_9724;
wire n_13430;
wire n_3996;
wire n_4221;
wire n_8243;
wire n_10226;
wire n_11117;
wire n_8236;
wire n_14964;
wire n_11046;
wire n_8292;
wire n_14640;
wire n_14901;
wire n_11547;
wire n_12676;
wire n_13327;
wire n_4181;
wire n_14412;
wire n_14391;
wire n_5777;
wire n_7949;
wire n_8611;
wire n_7046;
wire n_12720;
wire n_4225;
wire n_10475;
wire n_13365;
wire n_10020;
wire n_9826;
wire n_5142;
wire n_14195;
wire n_10467;
wire n_4153;
wire n_5156;
wire n_13118;
wire n_5926;
wire n_8011;
wire n_9839;
wire n_14431;
wire n_4300;
wire n_9399;
wire n_4783;
wire n_12535;
wire n_14254;
wire n_13279;
wire n_3769;
wire n_12283;
wire n_12506;
wire n_14044;
wire n_6589;
wire n_7579;
wire n_4530;
wire n_4267;
wire n_8139;
wire n_12046;
wire n_8123;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_10720;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_10907;
wire n_6197;
wire n_6971;
wire n_9938;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_13844;
wire n_14462;
wire n_11256;
wire n_7460;
wire n_9658;
wire n_11914;
wire n_9605;
wire n_12124;
wire n_11934;
wire n_14731;
wire n_10868;
wire n_11047;
wire n_9013;
wire n_14004;
wire n_8730;
wire n_9417;
wire n_13945;
wire n_14841;
wire n_8156;
wire n_9290;
wire n_9212;
wire n_13431;
wire n_13342;
wire n_9721;
wire n_14913;
wire n_14789;
wire n_12189;
wire n_10615;
wire n_7698;
wire n_12884;
wire n_13187;
wire n_7886;
wire n_6154;
wire n_7344;
wire n_14504;
wire n_6020;
wire n_13082;
wire n_9586;
wire n_7904;
wire n_12310;
wire n_11004;
wire n_4182;
wire n_10751;
wire n_12683;
wire n_13821;
wire n_11287;
wire n_5701;
wire n_4825;
wire n_10706;
wire n_4440;
wire n_10774;
wire n_11208;
wire n_4549;
wire n_12108;
wire n_12502;
wire n_3955;
wire n_9104;
wire n_7079;
wire n_10225;
wire n_11963;
wire n_10570;
wire n_9293;
wire n_11860;
wire n_13298;
wire n_5120;
wire n_8645;
wire n_10744;
wire n_11625;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_10416;
wire n_4303;
wire n_4574;
wire n_14933;
wire n_7774;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_8618;
wire n_6696;
wire n_11181;
wire n_11787;
wire n_14024;
wire n_5222;
wire n_4839;
wire n_13810;
wire n_8285;
wire n_5743;
wire n_4016;
wire n_9919;
wire n_10396;
wire n_8826;
wire n_6210;
wire n_10123;
wire n_5772;
wire n_12899;
wire n_14252;
wire n_8715;
wire n_12761;
wire n_14522;
wire n_8782;
wire n_6964;
wire n_14399;
wire n_10083;
wire n_5801;
wire n_6117;
wire n_14331;
wire n_4231;
wire n_8117;
wire n_12918;
wire n_11825;
wire n_6202;
wire n_7279;
wire n_7670;
wire n_11364;
wire n_4923;
wire n_12713;
wire n_3652;
wire n_14126;
wire n_12522;
wire n_12822;
wire n_9445;
wire n_14148;
wire n_4097;
wire n_14031;
wire n_6681;
wire n_13539;
wire n_5971;
wire n_4083;
wire n_11420;
wire n_12223;
wire n_13532;
wire n_11470;
wire n_4461;
wire n_13089;
wire n_5392;
wire n_8497;
wire n_12082;
wire n_9930;
wire n_6661;
wire n_8018;
wire n_6640;
wire n_12151;
wire n_3916;
wire n_13335;
wire n_7940;
wire n_14493;
wire n_11230;
wire n_12757;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_10731;
wire n_11063;
wire n_10347;
wire n_11074;
wire n_13411;
wire n_6455;
wire n_7721;
wire n_9727;
wire n_4273;
wire n_15034;
wire n_7606;
wire n_5443;
wire n_12025;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_10926;
wire n_6644;
wire n_13879;
wire n_13848;
wire n_14534;
wire n_4389;
wire n_6896;
wire n_14475;
wire n_3930;
wire n_12183;
wire n_14633;
wire n_4448;
wire n_11669;
wire n_10734;
wire n_6832;
wire n_8798;
wire n_7836;
wire n_12143;
wire n_6160;
wire n_14473;
wire n_7564;
wire n_11493;
wire n_12158;
wire n_7884;
wire n_8673;
wire n_10281;
wire n_6718;
wire n_9685;
wire n_11486;
wire n_8502;
wire n_6542;
wire n_10126;
wire n_10759;
wire n_13293;
wire n_11786;
wire n_10650;
wire n_14083;
wire n_11777;
wire n_6031;
wire n_5568;
wire n_5502;
wire n_9421;
wire n_8577;
wire n_11722;
wire n_14487;
wire n_7653;
wire n_10092;
wire n_10445;
wire n_5656;
wire n_8531;
wire n_8635;
wire n_6763;
wire n_4831;
wire n_5974;
wire n_9567;
wire n_6280;
wire n_9298;
wire n_11941;
wire n_10116;
wire n_6438;
wire n_13614;
wire n_10048;
wire n_9059;
wire n_12937;
wire n_8485;
wire n_3662;
wire n_13285;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_13596;
wire n_8872;
wire n_8752;
wire n_13609;
wire n_9396;
wire n_5413;
wire n_6758;
wire n_4596;
wire n_12459;
wire n_13715;
wire n_13398;
wire n_7976;
wire n_9234;
wire n_9425;
wire n_12648;
wire n_10364;
wire n_5412;
wire n_9620;
wire n_3694;
wire n_6069;
wire n_10963;
wire n_5752;
wire n_10191;
wire n_6874;
wire n_13330;
wire n_4726;
wire n_13235;
wire n_4751;
wire n_4222;
wire n_8341;
wire n_13412;
wire n_13995;
wire n_14867;
wire n_12638;
wire n_8521;
wire n_6030;
wire n_11209;
wire n_8199;
wire n_12976;
wire n_13091;
wire n_13306;
wire n_13561;
wire n_6077;
wire n_8005;
wire n_11718;
wire n_4119;
wire n_3799;
wire n_7743;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_9517;
wire n_4474;
wire n_6386;
wire n_9639;
wire n_9192;
wire n_14128;
wire n_12762;
wire n_9102;
wire n_5217;
wire n_10003;
wire n_10025;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_5957;
wire n_12066;
wire n_11234;
wire n_12021;
wire n_14822;
wire n_8283;
wire n_13016;
wire n_13048;
wire n_10502;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_8291;
wire n_4214;
wire n_8176;
wire n_10674;
wire n_5158;
wire n_4884;
wire n_14942;
wire n_6708;
wire n_7737;
wire n_10179;
wire n_14076;
wire n_7433;
wire n_11000;
wire n_12447;
wire n_13939;
wire n_11702;
wire n_4366;
wire n_10466;
wire n_12667;
wire n_4009;
wire n_12221;
wire n_7347;
wire n_8145;
wire n_9487;
wire n_10268;
wire n_4580;
wire n_13560;
wire n_6792;
wire n_14389;
wire n_12906;
wire n_7633;
wire n_12851;
wire n_6177;
wire n_5912;
wire n_11431;
wire n_10679;
wire n_12691;
wire n_7798;
wire n_10492;
wire n_11177;
wire n_12980;
wire n_4129;
wire n_4871;
wire n_12416;
wire n_13436;
wire n_4999;
wire n_13023;
wire n_13985;
wire n_11454;
wire n_6033;
wire n_9221;
wire n_12989;
wire n_11418;
wire n_5557;
wire n_7397;
wire n_12739;
wire n_7389;
wire n_13074;
wire n_12791;
wire n_5472;
wire n_7602;
wire n_13920;
wire n_13795;
wire n_14483;
wire n_4112;
wire n_8069;
wire n_6002;
wire n_14696;
wire n_14571;
wire n_14753;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_14903;
wire n_5396;
wire n_7693;
wire n_14052;
wire n_5335;
wire n_8888;
wire n_12650;
wire n_12319;
wire n_6557;
wire n_7300;
wire n_9566;
wire n_12692;
wire n_12403;
wire n_14908;
wire n_9578;
wire n_8483;
wire n_14820;
wire n_8797;
wire n_5960;
wire n_8605;
wire n_8041;
wire n_4236;
wire n_9868;
wire n_13451;
wire n_14778;
wire n_5002;
wire n_11750;
wire n_14124;
wire n_14442;
wire n_11572;
wire n_7532;
wire n_11038;
wire n_11049;
wire n_9292;
wire n_10460;
wire n_13363;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_12669;
wire n_11491;
wire n_14838;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_11109;
wire n_5859;
wire n_10968;
wire n_8760;
wire n_4734;
wire n_8928;
wire n_10004;
wire n_11894;
wire n_10729;
wire n_13689;
wire n_8374;
wire n_14276;
wire n_8917;
wire n_6163;
wire n_4635;
wire n_10811;
wire n_7118;
wire n_14540;
wire n_8006;
wire n_11806;
wire n_4013;
wire n_9884;
wire n_11504;
wire n_6778;
wire n_6285;
wire n_7946;
wire n_8723;
wire n_9857;
wire n_11737;
wire n_12127;
wire n_11637;
wire n_6025;
wire n_14622;
wire n_13769;
wire n_8957;
wire n_12058;
wire n_7257;
wire n_4242;
wire n_11799;
wire n_10944;
wire n_11788;
wire n_13537;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_13143;
wire n_13808;
wire n_10140;
wire n_12868;
wire n_14226;
wire n_12642;
wire n_10013;
wire n_14106;
wire n_12600;
wire n_7933;
wire n_5283;
wire n_8409;
wire n_9815;
wire n_9110;
wire n_7669;
wire n_5268;
wire n_10110;
wire n_13909;
wire n_6318;
wire n_10133;
wire n_14531;
wire n_14720;
wire n_8215;
wire n_11453;
wire n_11184;
wire n_8220;
wire n_9471;
wire n_9048;
wire n_4561;
wire n_7927;
wire n_11356;
wire n_6089;
wire n_4021;
wire n_8629;
wire n_3880;
wire n_13045;
wire n_5122;
wire n_7910;
wire n_11955;
wire n_12005;
wire n_13426;
wire n_14596;
wire n_6315;
wire n_10592;
wire n_14887;
wire n_7970;
wire n_14172;
wire n_4955;
wire n_10476;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_14147;
wire n_12953;
wire n_14593;
wire n_13507;
wire n_11488;
wire n_13040;
wire n_12369;
wire n_9394;
wire n_3650;
wire n_8991;
wire n_12300;
wire n_5840;
wire n_13015;
wire n_14934;
wire n_6343;
wire n_10186;
wire n_11938;
wire n_14988;
wire n_11946;
wire n_9191;
wire n_11918;
wire n_9004;
wire n_12832;
wire n_13839;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_7865;
wire n_6052;
wire n_11412;
wire n_13522;
wire n_10700;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_12290;
wire n_13208;
wire n_6886;
wire n_13761;
wire n_14219;
wire n_12169;
wire n_8783;
wire n_6912;
wire n_8326;
wire n_10496;
wire n_11249;
wire n_13538;
wire n_10521;
wire n_12838;
wire n_5914;
wire n_14523;
wire n_11464;
wire n_12325;
wire n_8504;
wire n_10695;
wire n_14763;
wire n_8445;
wire n_11950;
wire n_13847;
wire n_11648;
wire n_8250;
wire n_10994;
wire n_11576;
wire n_4715;
wire n_5039;
wire n_9118;
wire n_13950;
wire n_6061;
wire n_4369;
wire n_14025;
wire n_15006;
wire n_12969;
wire n_13214;
wire n_5378;
wire n_10758;
wire n_13559;
wire n_8408;
wire n_4543;
wire n_10120;
wire n_11410;
wire n_4941;
wire n_11251;
wire n_7252;
wire n_5542;
wire n_4394;
wire n_9051;
wire n_7133;
wire n_6883;
wire n_10345;
wire n_13065;
wire n_5519;
wire n_12809;
wire n_9908;
wire n_12748;
wire n_13639;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_8155;
wire n_5278;
wire n_8818;
wire n_11641;
wire n_12264;
wire n_11633;
wire n_7518;
wire n_9123;
wire n_12352;
wire n_5586;
wire n_13221;
wire n_10232;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_8660;
wire n_5187;
wire n_4944;
wire n_13619;
wire n_12054;
wire n_5675;
wire n_14055;
wire n_4135;
wire n_8275;
wire n_9327;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_11555;
wire n_9687;
wire n_14552;
wire n_8297;
wire n_9828;
wire n_6749;
wire n_13921;
wire n_11984;
wire n_14355;
wire n_6839;
wire n_10533;
wire n_13053;
wire n_14448;
wire n_9519;
wire n_10611;
wire n_7711;
wire n_13635;
wire n_12368;
wire n_10089;
wire n_12137;
wire n_3744;
wire n_4263;
wire n_11651;
wire n_14038;
wire n_7705;
wire n_10455;
wire n_8590;
wire n_6051;
wire n_4716;
wire n_12538;
wire n_4942;
wire n_6217;
wire n_13671;
wire n_6680;
wire n_5844;
wire n_12016;
wire n_7972;
wire n_15075;
wire n_6532;
wire n_13517;
wire n_6155;
wire n_4745;
wire n_6446;
wire n_8072;
wire n_12644;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_7854;
wire n_7707;
wire n_10632;
wire n_12017;
wire n_13428;
wire n_11672;
wire n_11696;
wire n_3907;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_6526;
wire n_8142;
wire n_10820;
wire n_14914;
wire n_10601;
wire n_13455;
wire n_6339;
wire n_4629;
wire n_14594;
wire n_12197;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_12892;
wire n_5662;
wire n_4857;
wire n_14213;
wire n_9802;
wire n_9315;
wire n_9296;
wire n_8599;
wire n_10447;
wire n_4080;
wire n_12373;
wire n_12660;
wire n_14393;
wire n_4226;
wire n_4741;
wire n_10022;
wire n_14526;
wire n_5265;
wire n_4752;
wire n_14184;
wire n_11567;
wire n_10305;
wire n_14769;
wire n_12855;
wire n_14795;
wire n_3986;
wire n_4376;
wire n_10031;
wire n_12877;
wire n_5705;
wire n_4753;
wire n_12350;
wire n_14691;
wire n_14576;
wire n_13137;
wire n_10798;
wire n_12388;
wire n_4552;
wire n_7656;
wire n_10760;
wire n_11202;
wire n_6845;
wire n_3885;
wire n_9405;
wire n_14647;
wire n_12891;
wire n_9302;
wire n_7105;
wire n_5196;
wire n_12836;
wire n_13892;
wire n_5181;
wire n_13636;
wire n_11779;
wire n_11888;
wire n_10166;
wire n_14317;
wire n_15024;
wire n_3709;
wire n_6829;
wire n_11684;
wire n_11879;
wire n_5574;
wire n_11054;
wire n_5126;
wire n_6508;
wire n_9842;
wire n_9977;
wire n_9887;
wire n_14893;
wire n_4067;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_7570;
wire n_8246;
wire n_11116;
wire n_9524;
wire n_11129;
wire n_7771;
wire n_4385;
wire n_13742;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_5368;
wire n_9322;
wire n_11937;
wire n_10098;
wire n_15079;
wire n_10510;
wire n_13905;
wire n_13934;
wire n_10848;
wire n_10042;
wire n_8057;
wire n_9122;
wire n_8349;
wire n_5626;
wire n_9333;
wire n_13240;
wire n_8743;
wire n_6603;
wire n_6114;
wire n_14073;
wire n_9590;
wire n_13515;
wire n_6576;
wire n_3651;
wire n_7943;
wire n_4333;
wire n_7364;
wire n_8473;
wire n_10993;
wire n_13838;
wire n_10342;
wire n_7208;
wire n_12286;
wire n_6245;
wire n_12992;
wire n_14132;
wire n_10439;
wire n_11923;
wire n_12844;
wire n_14284;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_13868;
wire n_9676;
wire n_3789;
wire n_10444;
wire n_7714;
wire n_9902;
wire n_10054;
wire n_12759;
wire n_8535;
wire n_10728;
wire n_4815;
wire n_9621;
wire n_13175;
wire n_7202;
wire n_9140;
wire n_4246;
wire n_9604;
wire n_7011;
wire n_4609;
wire n_13759;
wire n_7621;
wire n_5291;
wire n_8068;
wire n_10565;
wire n_10540;
wire n_14444;
wire n_12935;
wire n_9821;
wire n_11943;
wire n_14158;
wire n_10748;
wire n_5876;
wire n_10178;
wire n_11995;
wire n_11058;
wire n_6970;
wire n_11842;
wire n_12076;
wire n_12790;
wire n_12979;
wire n_5114;
wire n_6409;
wire n_6704;
wire n_6876;
wire n_4088;
wire n_12659;
wire n_7778;
wire n_3682;
wire n_4357;
wire n_9343;
wire n_7028;
wire n_12532;
wire n_4472;
wire n_4462;
wire n_7313;
wire n_7320;
wire n_6255;
wire n_14437;
wire n_7343;
wire n_5288;
wire n_5540;
wire n_5699;
wire n_11473;
wire n_7525;
wire n_13735;
wire n_7875;
wire n_5810;
wire n_11568;
wire n_14384;
wire n_13258;
wire n_4148;
wire n_4151;
wire n_13617;
wire n_12702;
wire n_6938;
wire n_12050;
wire n_4373;
wire n_12138;
wire n_5762;
wire n_13713;
wire n_4934;
wire n_5218;
wire n_8785;
wire n_9952;
wire n_12473;
wire n_13013;
wire n_14577;
wire n_10686;
wire n_8327;
wire n_12606;
wire n_9219;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_13625;
wire n_4630;
wire n_5408;
wire n_10971;
wire n_6427;
wire n_4331;
wire n_4643;
wire n_13051;
wire n_13054;
wire n_4475;
wire n_3989;
wire n_7753;
wire n_10076;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_11924;
wire n_12374;
wire n_8168;
wire n_14837;
wire n_14266;
wire n_14064;
wire n_8392;
wire n_7038;
wire n_12967;
wire n_14745;
wire n_4683;
wire n_5366;
wire n_10132;
wire n_10282;
wire n_13649;
wire n_9872;
wire n_12956;
wire n_6360;
wire n_11203;
wire n_13026;
wire n_9553;
wire n_10900;
wire n_6146;
wire n_10616;
wire n_9447;
wire n_6270;
wire n_11585;
wire n_9150;
wire n_3706;
wire n_5477;
wire n_9592;
wire n_5451;
wire n_9984;
wire n_12695;
wire n_3923;
wire n_14111;
wire n_11416;
wire n_4696;
wire n_11526;
wire n_11742;
wire n_13855;
wire n_12179;
wire n_8419;
wire n_11809;
wire n_5086;
wire n_9814;
wire n_10858;
wire n_12038;
wire n_5901;
wire n_6353;
wire n_14359;
wire n_4011;
wire n_10769;
wire n_9446;
wire n_4905;
wire n_14689;
wire n_15088;
wire n_10211;
wire n_10023;
wire n_11877;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_12105;
wire n_9461;
wire n_10772;
wire n_9793;
wire n_6691;
wire n_3748;
wire n_8997;
wire n_14324;
wire n_4278;
wire n_13184;
wire n_4623;
wire n_4910;
wire n_12360;
wire n_12297;
wire n_4410;
wire n_12952;
wire n_9874;
wire n_13332;
wire n_7392;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_14567;
wire n_6239;
wire n_4553;
wire n_6803;
wire n_10446;
wire n_11735;
wire n_14981;
wire n_7919;
wire n_15050;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_14281;
wire n_4809;
wire n_14876;
wire n_8109;
wire n_5226;
wire n_7657;
wire n_3660;
wire n_14129;
wire n_7995;
wire n_11405;
wire n_5867;
wire n_6048;
wire n_8985;
wire n_13318;
wire n_14733;
wire n_5079;
wire n_5590;
wire n_10331;
wire n_12103;
wire n_6773;
wire n_9403;
wire n_3833;
wire n_5632;
wire n_14515;
wire n_8390;
wire n_11480;
wire n_11874;
wire n_4841;
wire n_12115;
wire n_6336;
wire n_3814;
wire n_8463;
wire n_14120;
wire n_7041;
wire n_7802;
wire n_4842;
wire n_4911;
wire n_14243;
wire n_4340;
wire n_7370;
wire n_13366;
wire n_10181;
wire n_10074;
wire n_9731;
wire n_5660;
wire n_11104;
wire n_13677;
wire n_4645;
wire n_7557;
wire n_11862;
wire n_11952;
wire n_14529;
wire n_6174;
wire n_3725;
wire n_4920;
wire n_12828;
wire n_4972;
wire n_13322;
wire n_6023;
wire n_6776;
wire n_14894;
wire n_13078;
wire n_5426;
wire n_9947;
wire n_6463;
wire n_13387;
wire n_14370;
wire n_7896;
wire n_13226;
wire n_9699;
wire n_6372;
wire n_10962;
wire n_11037;
wire n_9305;
wire n_10481;
wire n_14624;
wire n_7176;
wire n_12003;
wire n_14194;
wire n_14868;
wire n_10220;
wire n_13917;
wire n_10381;
wire n_8517;
wire n_12332;
wire n_5778;
wire n_5625;
wire n_6396;
wire n_10642;
wire n_9218;
wire n_13317;
wire n_11556;
wire n_3917;
wire n_6669;
wire n_9096;
wire n_10634;
wire n_3942;
wire n_13480;
wire n_10170;
wire n_10142;
wire n_10569;
wire n_12326;
wire n_3765;
wire n_14489;
wire n_5531;
wire n_9534;
wire n_7826;
wire n_5429;
wire n_11044;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_11042;
wire n_12141;
wire n_4451;
wire n_6394;
wire n_9164;
wire n_9546;
wire n_3844;
wire n_12622;
wire n_11226;
wire n_4054;
wire n_5448;
wire n_7590;
wire n_5432;
wire n_14977;
wire n_13732;
wire n_9358;
wire n_11985;
wire n_5160;
wire n_11328;
wire n_13545;
wire n_8208;
wire n_6995;
wire n_7185;
wire n_10127;
wire n_14214;
wire n_11525;
wire n_3988;
wire n_9730;
wire n_6254;
wire n_6161;
wire n_13246;
wire n_9066;
wire n_10800;
wire n_11020;
wire n_9185;
wire n_9318;
wire n_10374;
wire n_8134;
wire n_7987;
wire n_14367;
wire n_4324;
wire n_4821;
wire n_10328;
wire n_8631;
wire n_14542;
wire n_5445;
wire n_8694;
wire n_11892;
wire n_8965;
wire n_8647;
wire n_13288;
wire n_11013;
wire n_12343;
wire n_7332;
wire n_6660;
wire n_5719;
wire n_4771;
wire n_7225;
wire n_10529;
wire n_12396;
wire n_13823;
wire n_6128;
wire n_4086;
wire n_7037;
wire n_11820;
wire n_14900;
wire n_11587;
wire n_14863;
wire n_4814;
wire n_12081;
wire n_13157;
wire n_10314;
wire n_14966;
wire n_3648;
wire n_5749;
wire n_11697;
wire n_12296;
wire n_8427;
wire n_9339;
wire n_5332;
wire n_13038;
wire n_9596;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_10006;
wire n_10667;
wire n_7258;
wire n_7432;
wire n_9156;
wire n_11441;
wire n_11242;
wire n_3701;
wire n_11916;
wire n_14591;
wire n_11435;
wire n_12804;
wire n_13999;
wire n_11471;
wire n_6334;
wire n_10346;
wire n_13236;
wire n_8984;
wire n_6848;
wire n_14502;
wire n_10539;
wire n_8345;
wire n_10414;
wire n_6321;
wire n_7765;
wire n_4708;
wire n_9708;
wire n_9268;
wire n_8764;
wire n_6794;
wire n_10340;
wire n_4826;
wire n_13310;
wire n_10245;
wire n_14479;
wire n_11644;
wire n_7761;
wire n_7197;
wire n_12466;
wire n_12701;
wire n_5489;
wire n_12106;
wire n_6400;
wire n_3767;
wire n_12560;
wire n_4589;
wire n_9097;
wire n_5057;
wire n_10280;
wire n_12895;
wire n_11432;
wire n_4578;
wire n_12342;
wire n_6705;
wire n_7775;
wire n_9636;
wire n_10256;
wire n_14559;
wire n_14676;
wire n_7619;
wire n_12125;
wire n_5436;
wire n_5907;
wire n_11120;
wire n_5072;
wire n_11391;
wire n_6044;
wire n_11164;
wire n_11527;
wire n_3674;
wire n_5286;
wire n_8083;
wire n_8853;
wire n_11371;
wire n_6495;
wire n_5013;
wire n_10917;
wire n_7403;
wire n_13933;
wire n_6902;
wire n_6470;
wire n_14619;
wire n_9473;
wire n_10727;
wire n_11591;
wire n_10145;
wire n_12341;
wire n_9560;
wire n_5569;
wire n_8038;
wire n_10938;
wire n_9175;
wire n_8711;
wire n_10976;
wire n_5439;
wire n_8229;
wire n_8949;
wire n_14248;
wire n_14928;
wire n_10612;
wire n_5619;
wire n_4147;
wire n_6481;
wire n_9810;
wire n_14079;
wire n_7548;
wire n_4925;
wire n_9244;
wire n_14878;
wire n_9584;
wire n_12047;
wire n_6534;
wire n_11460;
wire n_13289;
wire n_4974;
wire n_8567;
wire n_10797;
wire n_13320;
wire n_9439;
wire n_11915;
wire n_14224;
wire n_13210;
wire n_14015;
wire n_4932;
wire n_4510;
wire n_8655;
wire n_9235;
wire n_6181;
wire n_6728;
wire n_8705;
wire n_11642;
wire n_9043;
wire n_9768;
wire n_11306;
wire n_3787;
wire n_14566;
wire n_13549;
wire n_5119;
wire n_9037;
wire n_5715;
wire n_9085;
wire n_12434;
wire n_8085;
wire n_14874;
wire n_8777;
wire n_6133;
wire n_11891;
wire n_14951;
wire n_8852;
wire n_9264;
wire n_6528;
wire n_10114;
wire n_7604;
wire n_7407;
wire n_14499;
wire n_8185;
wire n_3827;
wire n_12998;
wire n_13427;
wire n_10845;
wire n_4447;
wire n_8513;
wire n_6670;
wire n_12248;
wire n_14155;
wire n_6774;
wire n_8365;
wire n_11007;
wire n_14229;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_11557;
wire n_12405;
wire n_6038;
wire n_4818;
wire n_7727;
wire n_4514;
wire n_4800;
wire n_10599;
wire n_11231;
wire n_3960;
wire n_9550;
wire n_9836;
wire n_13228;
wire n_6282;
wire n_13244;
wire n_9929;
wire n_12134;
wire n_8035;
wire n_8505;
wire n_11399;
wire n_11092;
wire n_4433;
wire n_11163;
wire n_8874;
wire n_11542;
wire n_10008;
wire n_6700;
wire n_7334;
wire n_7684;
wire n_7755;
wire n_8098;
wire n_4341;
wire n_10623;
wire n_9187;
wire n_13880;
wire n_11276;
wire n_4312;
wire n_10511;
wire n_5932;
wire n_12770;
wire n_13011;
wire n_14418;
wire n_6178;
wire n_11575;
wire n_10503;
wire n_6234;
wire n_14880;
wire n_11732;
wire n_6012;
wire n_4633;
wire n_14518;
wire n_9406;
wire n_3838;
wire n_10857;
wire n_9342;
wire n_13323;
wire n_4277;
wire n_13222;
wire n_13604;
wire n_14119;
wire n_14321;
wire n_7787;
wire n_14808;
wire n_4140;
wire n_8067;
wire n_3675;
wire n_12421;
wire n_5092;
wire n_10708;
wire n_14136;
wire n_13106;
wire n_14950;
wire n_7849;
wire n_5186;
wire n_12550;
wire n_13126;
wire n_11045;
wire n_7367;
wire n_8619;
wire n_9851;
wire n_9559;
wire n_11993;
wire n_14818;
wire n_11508;
wire n_12755;
wire n_8679;
wire n_9806;
wire n_8644;
wire n_12306;
wire n_12965;
wire n_11982;
wire n_10516;
wire n_4662;
wire n_3779;
wire n_6715;
wire n_11395;
wire n_5828;
wire n_11634;
wire n_7200;
wire n_13068;
wire n_9860;
wire n_4882;
wire n_4993;
wire n_11887;
wire n_11301;
wire n_15031;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_13402;
wire n_6337;
wire n_13997;
wire n_4868;
wire n_8923;
wire n_8970;
wire n_8332;
wire n_10119;
wire n_14302;
wire n_10548;
wire n_11010;
wire n_11408;
wire n_8632;
wire n_14829;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_8876;
wire n_3925;
wire n_10733;
wire n_10547;
wire n_11670;
wire n_13218;
wire n_14011;
wire n_5238;
wire n_10067;
wire n_14646;
wire n_13958;
wire n_13239;
wire n_4059;
wire n_8856;
wire n_12603;
wire n_14230;
wire n_11604;
wire n_9240;
wire n_4595;
wire n_7877;
wire n_11506;
wire n_11666;
wire n_8945;
wire n_11503;
wire n_8918;
wire n_14433;
wire n_7799;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_11857;
wire n_5631;
wire n_8028;
wire n_6539;
wire n_7243;
wire n_7179;
wire n_9345;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_10222;
wire n_11193;
wire n_13983;
wire n_11293;
wire n_12439;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_8774;
wire n_5326;
wire n_12072;
wire n_14199;
wire n_8779;
wire n_13949;
wire n_8968;
wire n_13941;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_8404;
wire n_4669;
wire n_13090;
wire n_6595;
wire n_4339;
wire n_12558;
wire n_12244;
wire n_12199;
wire n_11214;
wire n_4041;
wire n_5459;
wire n_7738;
wire n_13851;
wire n_14209;
wire n_14986;
wire n_4060;
wire n_9223;
wire n_9499;
wire n_10647;
wire n_14177;
wire n_14495;
wire n_11362;
wire n_11288;
wire n_11409;
wire n_15091;
wire n_5528;
wire n_13036;
wire n_11027;
wire n_12996;
wire n_5391;
wire n_12873;
wire n_8073;
wire n_4541;
wire n_5422;
wire n_3824;
wire n_7785;
wire n_13225;
wire n_6385;
wire n_14485;
wire n_6289;
wire n_12591;
wire n_5267;
wire n_4494;
wire n_10581;
wire n_13587;
wire n_5523;
wire n_4796;
wire n_7373;
wire n_9576;
wire n_9120;
wire n_14832;
wire n_14917;
wire n_10097;
wire n_10405;
wire n_15009;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_12726;
wire n_9651;
wire n_12833;
wire n_14206;
wire n_6257;
wire n_14240;
wire n_12690;
wire n_11031;
wire n_14080;
wire n_13076;
wire n_9386;
wire n_11285;
wire n_10813;
wire n_6852;
wire n_6346;
wire n_11346;
wire n_12618;
wire n_4775;
wire n_9779;
wire n_5044;
wire n_5809;
wire n_12414;
wire n_11513;
wire n_5365;
wire n_14888;
wire n_7587;
wire n_13729;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_11250;
wire n_7874;
wire n_3886;
wire n_11340;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_14381;
wire n_14739;
wire n_7372;
wire n_7760;
wire n_10588;
wire n_4248;
wire n_9635;
wire n_5915;
wire n_6818;
wire n_9444;
wire n_10943;
wire n_11190;
wire n_5452;
wire n_7226;
wire n_8930;
wire n_4754;
wire n_13992;
wire n_7057;
wire n_12736;
wire n_7685;
wire n_8031;
wire n_11818;
wire n_8750;
wire n_14193;
wire n_14649;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_6815;
wire n_6753;
wire n_4845;
wire n_9364;
wire n_9581;
wire n_9512;
wire n_9317;
wire n_3893;
wire n_14625;
wire n_14661;
wire n_14968;
wire n_8593;
wire n_14047;
wire n_13592;
wire n_4585;
wire n_7730;
wire n_14262;
wire n_14723;
wire n_13165;
wire n_8509;
wire n_9314;
wire n_9459;
wire n_8405;
wire n_13659;
wire n_14558;
wire n_9549;
wire n_11564;
wire n_10641;
wire n_7913;
wire n_4383;
wire n_11719;
wire n_8492;
wire n_6764;
wire n_14569;
wire n_5535;
wire n_9275;
wire n_3875;
wire n_13670;
wire n_15102;
wire n_10210;
wire n_5370;
wire n_11944;
wire n_13967;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_4003;
wire n_13248;
wire n_11785;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_5594;
wire n_4301;
wire n_11754;
wire n_4586;
wire n_14369;
wire n_4048;
wire n_14301;
wire n_9865;
wire n_6471;
wire n_11075;
wire n_11511;
wire n_12981;
wire n_13061;
wire n_13546;
wire n_3777;
wire n_6627;
wire n_10027;
wire n_5761;
wire n_10263;
wire n_10722;
wire n_14422;
wire n_13005;
wire n_13978;
wire n_11771;
wire n_4784;
wire n_7203;
wire n_8429;
wire n_8854;
wire n_9757;
wire n_7512;
wire n_5550;
wire n_12333;
wire n_11912;
wire n_5082;
wire n_4046;
wire n_9656;
wire n_10426;
wire n_11284;
wire n_5209;
wire n_7215;
wire n_10246;
wire n_13500;
wire n_6636;
wire n_15033;
wire n_4199;
wire n_13004;
wire n_10617;
wire n_5929;
wire n_10909;
wire n_5559;
wire n_12694;
wire n_13972;
wire n_14295;
wire n_5478;
wire n_11298;
wire n_7388;
wire n_7694;
wire n_6243;
wire n_6488;
wire n_4286;
wire n_9629;
wire n_13864;
wire n_11185;
wire n_5102;
wire n_11498;
wire n_6022;
wire n_8686;
wire n_6457;
wire n_10299;
wire n_4470;
wire n_12904;
wire n_7982;
wire n_13874;
wire n_11384;
wire n_10763;
wire n_10494;
wire n_4058;
wire n_13520;
wire n_3664;
wire n_8773;
wire n_10743;
wire n_8225;
wire n_8583;
wire n_4188;
wire n_3913;
wire n_6867;
wire n_8887;
wire n_9556;
wire n_5868;
wire n_6538;
wire n_6230;
wire n_4034;
wire n_12810;
wire n_9259;
wire n_9995;
wire n_14680;
wire n_12820;
wire n_6633;
wire n_9371;
wire n_8080;
wire n_11496;
wire n_6187;
wire n_6172;
wire n_13274;
wire n_10050;
wire n_13827;
wire n_5275;
wire n_14927;
wire n_10702;
wire n_4689;
wire n_13572;
wire n_14236;
wire n_5071;
wire n_7311;
wire n_5989;
wire n_8964;
wire n_11768;
wire n_15051;
wire n_12085;
wire n_14748;
wire n_9008;
wire n_6574;
wire n_11388;
wire n_11683;
wire n_13786;
wire n_8929;
wire n_8539;
wire n_6395;
wire n_4402;
wire n_9484;
wire n_8745;
wire n_4239;
wire n_6854;
wire n_7996;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_8776;
wire n_8588;
wire n_8554;
wire n_9319;
wire n_11748;
wire n_7488;
wire n_5227;
wire n_13463;
wire n_9442;
wire n_14351;
wire n_10165;
wire n_14385;
wire n_7198;
wire n_4201;
wire n_10366;
wire n_12207;
wire n_8802;
wire n_13242;
wire n_13194;
wire n_9587;
wire n_6784;
wire n_14915;
wire n_6168;
wire n_13871;
wire n_14168;
wire n_9904;
wire n_9157;
wire n_8431;
wire n_8453;
wire n_6766;
wire n_5242;
wire n_8955;
wire n_3704;
wire n_12510;
wire n_8634;
wire n_14575;
wire n_4123;
wire n_6330;
wire n_5520;
wire n_8896;
wire n_14695;
wire n_3633;
wire n_4479;
wire n_7950;
wire n_7249;
wire n_13741;
wire n_9713;
wire n_11210;
wire n_9452;
wire n_10104;
wire n_14186;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_8837;
wire n_7031;
wire n_4539;
wire n_8907;
wire n_6799;
wire n_10115;
wire n_14514;
wire n_14853;
wire n_13654;
wire n_8015;
wire n_14149;
wire n_10397;
wire n_14454;
wire n_9974;
wire n_13245;
wire n_10398;
wire n_5920;
wire n_6672;
wire n_13193;
wire n_6149;
wire n_8256;
wire n_13739;
wire n_14578;
wire n_10065;
wire n_11156;
wire n_10243;
wire n_10087;
wire n_12628;
wire n_7142;
wire n_11598;
wire n_13977;
wire n_5808;
wire n_14003;
wire n_6054;
wire n_7089;
wire n_11176;
wire n_12687;
wire n_4682;
wire n_7916;
wire n_12260;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_6450;
wire n_12445;
wire n_13776;
wire n_3729;
wire n_8074;
wire n_12878;
wire n_14023;
wire n_4978;
wire n_4690;
wire n_10174;
wire n_12281;
wire n_10266;
wire n_12879;
wire n_10509;
wire n_12355;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_7042;
wire n_4736;
wire n_3780;
wire n_8778;
wire n_8039;
wire n_10415;
wire n_5244;
wire n_6523;
wire n_13127;
wire n_5382;
wire n_14581;
wire n_8065;
wire n_6107;
wire n_9634;
wire n_3957;
wire n_12601;
wire n_11893;
wire n_12004;
wire n_11828;
wire n_6775;
wire n_5274;
wire n_10873;
wire n_3848;
wire n_8194;
wire n_12291;
wire n_4284;
wire n_14125;
wire n_11582;
wire n_8207;
wire n_13109;
wire n_3919;
wire n_10106;
wire n_12474;
wire n_13414;
wire n_9241;
wire n_6232;
wire n_13688;
wire n_6445;
wire n_10422;
wire n_10736;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_9903;
wire n_8582;
wire n_10378;
wire n_6056;
wire n_8537;
wire n_6932;
wire n_13425;
wire n_7036;
wire n_4513;
wire n_3829;
wire n_9615;
wire n_4053;
wire n_8951;
wire n_7759;
wire n_9600;
wire n_11095;
wire n_7818;
wire n_11180;
wire n_9748;
wire n_9945;
wire n_5125;
wire n_12024;
wire n_4040;
wire n_9927;
wire n_5587;
wire n_6855;
wire n_14072;
wire n_11876;
wire n_5789;
wire n_8217;
wire n_10046;
wire n_13182;
wire n_14787;
wire n_13911;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_10954;
wire n_10388;
wire n_14883;
wire n_8437;
wire n_5249;
wire n_8849;
wire n_7447;
wire n_10659;
wire n_13124;
wire n_13956;
wire n_14617;
wire n_7944;
wire n_5198;
wire n_11709;
wire n_5360;
wire n_10804;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_9295;
wire n_5269;
wire n_13819;
wire n_11602;
wire n_11304;
wire n_6252;
wire n_12934;
wire n_5866;
wire n_6493;
wire n_14843;
wire n_8568;
wire n_10239;
wire n_12723;
wire n_7947;
wire n_12428;
wire n_4005;
wire n_10841;
wire n_12857;
wire n_13566;
wire n_14315;
wire n_9916;
wire n_4904;
wire n_8980;
wire n_13682;
wire n_5899;
wire n_11630;
wire n_13339;
wire n_7629;
wire n_13478;
wire n_8051;
wire n_7104;
wire n_4792;
wire n_8716;
wire n_11461;
wire n_3812;
wire n_9844;
wire n_7601;
wire n_4980;
wire n_11135;
wire n_12520;
wire n_14303;
wire n_11994;
wire n_12457;
wire n_12743;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_7757;
wire n_8030;
wire n_9316;
wire n_9663;
wire n_13918;
wire n_10168;
wire n_13526;
wire n_5865;
wire n_13019;
wire n_14335;
wire n_10075;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_14848;
wire n_3774;
wire n_14989;
wire n_10068;
wire n_11596;
wire n_10276;
wire n_12533;
wire n_8749;
wire n_11024;
wire n_7138;
wire n_7290;
wire n_14424;
wire n_8544;
wire n_13077;
wire n_13524;
wire n_8249;
wire n_12555;
wire n_9628;
wire n_14560;
wire n_6679;
wire n_8496;
wire n_9789;
wire n_14273;
wire n_13296;
wire n_13891;
wire n_4956;
wire n_14090;
wire n_5380;
wire n_5924;
wire n_12839;
wire n_7625;
wire n_5822;
wire n_10495;
wire n_9299;
wire n_12251;
wire n_6259;
wire n_7284;
wire n_4947;
wire n_11246;
wire n_14693;
wire n_11715;
wire n_4656;
wire n_12766;
wire n_12983;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_12573;
wire n_12945;
wire n_11970;
wire n_15047;
wire n_4729;
wire n_14839;
wire n_5786;
wire n_4987;
wire n_13466;
wire n_5182;
wire n_4971;
wire n_11113;
wire n_12451;
wire n_7971;
wire n_12542;
wire n_12376;
wire n_9022;
wire n_10927;
wire n_6630;
wire n_13116;
wire n_12585;
wire n_10704;
wire n_5658;
wire n_11613;
wire n_5388;
wire n_13256;
wire n_13968;
wire n_4823;
wire n_13942;
wire n_9427;
wire n_4875;
wire n_13231;
wire n_6279;
wire n_8698;
wire n_8695;
wire n_9344;
wire n_14461;
wire n_12530;
wire n_13718;
wire n_8751;
wire n_10603;
wire n_12875;
wire n_11085;
wire n_3762;
wire n_6813;
wire n_9764;
wire n_12808;
wire n_5564;
wire n_11294;
wire n_13024;
wire n_8273;
wire n_14897;
wire n_11021;
wire n_14041;
wire n_14817;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_14799;
wire n_7106;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_7644;
wire n_12494;
wire n_10011;
wire n_6057;
wire n_4137;
wire n_7529;
wire n_8986;
wire n_11905;
wire n_6675;
wire n_12488;
wire n_4529;
wire n_4323;
wire n_12229;
wire n_6476;
wire n_13740;
wire n_8200;
wire n_14397;
wire n_3972;
wire n_10055;
wire n_7907;
wire n_13064;
wire n_10982;
wire n_8188;
wire n_11926;
wire n_11951;
wire n_8528;
wire n_12219;
wire n_13041;
wire n_14879;
wire n_6207;
wire n_5539;
wire n_10764;
wire n_14333;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_9088;
wire n_12630;
wire n_6524;
wire n_10787;
wire n_5036;
wire n_12910;
wire n_5547;
wire n_4772;
wire n_6225;
wire n_4322;
wire n_8920;
wire n_8267;
wire n_12758;
wire n_13302;
wire n_10972;
wire n_7297;
wire n_6291;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_12883;
wire n_9734;
wire n_9505;
wire n_9664;
wire n_12672;
wire n_7199;
wire n_14167;
wire n_5273;
wire n_10262;
wire n_10826;
wire n_8360;
wire n_13828;
wire n_4677;
wire n_3901;
wire n_8036;
wire n_9510;
wire n_5261;
wire n_11423;
wire n_6520;
wire n_14162;
wire n_7853;
wire n_7648;
wire n_9413;
wire n_9888;
wire n_14085;
wire n_3757;
wire n_8393;
wire n_11484;
wire n_8821;
wire n_11760;
wire n_9863;
wire n_12946;
wire n_13397;
wire n_10881;
wire n_8160;
wire n_9199;
wire n_11370;
wire n_5193;
wire n_10707;
wire n_9014;
wire n_10204;
wire n_9411;
wire n_12394;
wire n_12706;
wire n_12613;
wire n_4909;
wire n_11909;
wire n_13882;
wire n_9336;
wire n_9360;
wire n_10556;
wire n_9543;
wire n_3635;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_13252;
wire n_14783;
wire n_5005;
wire n_13174;
wire n_3882;
wire n_7487;
wire n_10717;
wire n_6425;
wire n_13931;
wire n_5993;
wire n_3826;
wire n_13541;
wire n_12978;
wire n_14201;
wire n_12253;
wire n_14710;
wire n_7638;
wire n_8833;
wire n_14296;
wire n_5703;
wire n_8240;
wire n_12450;
wire n_14857;
wire n_7988;
wire n_4634;
wire n_13579;
wire n_9404;
wire n_14643;
wire n_8579;
wire n_6432;
wire n_5534;
wire n_14354;
wire n_9678;
wire n_12444;
wire n_8258;
wire n_9854;
wire n_7259;
wire n_11071;
wire n_11979;
wire n_13050;
wire n_8626;
wire n_13384;
wire n_12289;
wire n_6540;
wire n_6955;
wire n_9481;
wire n_5174;
wire n_10862;
wire n_4952;
wire n_12583;
wire n_5157;
wire n_13936;
wire n_4380;
wire n_9672;
wire n_14009;
wire n_9893;
wire n_4126;
wire n_7237;
wire n_8935;
wire n_11928;
wire n_5087;
wire n_12590;
wire n_3802;
wire n_6388;
wire n_4506;
wire n_12596;
wire n_10240;
wire n_5904;
wire n_9478;
wire n_13465;
wire n_4880;
wire n_11792;
wire n_9266;
wire n_9813;
wire n_12551;
wire n_14026;
wire n_6760;
wire n_13817;
wire n_8009;
wire n_11329;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_10205;
wire n_10338;
wire n_12034;
wire n_14275;
wire n_11573;
wire n_11703;
wire n_9042;
wire n_4943;
wire n_11671;
wire n_8012;
wire n_11445;
wire n_14692;
wire n_7576;
wire n_9506;
wire n_8608;
wire n_13946;
wire n_8008;
wire n_12498;
wire n_10285;
wire n_14040;
wire n_6795;
wire n_14464;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_12228;
wire n_5815;
wire n_12378;
wire n_11832;
wire n_6261;
wire n_5873;
wire n_4193;
wire n_4075;
wire n_13926;
wire n_9666;
wire n_10112;
wire n_14163;
wire n_6487;
wire n_9146;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_15046;
wire n_3647;
wire n_10056;
wire n_9862;
wire n_5755;
wire n_10283;
wire n_9274;
wire n_8702;
wire n_5949;
wire n_10469;
wire n_13944;
wire n_5195;
wire n_7483;
wire n_4136;
wire n_6608;
wire n_14145;
wire n_7858;
wire n_9619;
wire n_12742;
wire n_4393;
wire n_7385;
wire n_11088;
wire n_12423;
wire n_10618;
wire n_13902;
wire n_3720;
wire n_8576;
wire n_9508;
wire n_4535;
wire n_10105;
wire n_7668;
wire n_13008;
wire n_8662;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_13504;
wire n_5955;
wire n_7476;
wire n_15022;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_8436;
wire n_11154;
wire n_13491;
wire n_9987;
wire n_8124;
wire n_8148;
wire n_14135;
wire n_12518;
wire n_8033;
wire n_6843;
wire n_12764;
wire n_7953;
wire n_8343;
wire n_5246;
wire n_5964;
wire n_11065;
wire n_13812;
wire n_12417;
wire n_3724;
wire n_8118;
wire n_14182;
wire n_13751;
wire n_12209;
wire n_12882;
wire n_7266;
wire n_5164;
wire n_11449;
wire n_4196;
wire n_6969;
wire n_11447;
wire n_8741;
wire n_12427;
wire n_13894;
wire n_14217;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_14882;
wire n_5498;
wire n_7100;
wire n_15012;
wire n_4370;
wire n_14541;
wire n_5783;
wire n_11123;
wire n_8478;
wire n_5183;
wire n_11319;
wire n_11676;
wire n_6075;
wire n_7082;
wire n_9569;
wire n_6120;
wire n_6659;
wire n_13513;
wire n_6750;
wire n_11018;
wire n_5549;
wire n_9935;
wire n_14477;
wire n_9707;
wire n_13663;
wire n_14664;
wire n_8376;
wire n_3761;
wire n_9827;
wire n_7689;
wire n_13858;
wire n_4889;
wire n_7132;
wire n_11537;
wire n_8763;
wire n_13361;
wire n_5442;
wire n_13792;
wire n_5739;
wire n_7824;
wire n_8996;
wire n_12707;
wire n_13161;
wire n_9007;
wire n_4828;
wire n_9797;
wire n_13132;
wire n_6003;
wire n_5385;
wire n_8726;
wire n_13662;
wire n_8799;
wire n_4558;
wire n_7796;
wire n_10670;
wire n_9053;
wire n_6478;
wire n_6066;
wire n_9450;
wire n_13272;
wire n_12437;
wire n_7034;
wire n_6086;
wire n_9121;
wire n_6650;
wire n_4722;
wire n_6224;
wire n_10789;
wire n_14725;
wire n_10387;
wire n_8303;
wire n_8796;
wire n_4768;
wire n_12941;
wire n_10661;
wire n_13859;
wire n_11638;
wire n_14476;
wire n_4100;
wire n_10088;
wire n_12026;
wire n_10629;
wire n_14208;
wire n_13898;
wire n_7084;
wire n_5845;
wire n_9617;
wire n_9089;
wire n_8883;
wire n_7293;
wire n_10505;
wire n_8251;
wire n_10247;
wire n_9236;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_10860;
wire n_6060;
wire n_7253;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_12537;
wire n_14547;
wire n_9493;
wire n_8860;
wire n_14364;
wire n_8003;
wire n_6410;
wire n_12607;
wire n_5973;
wire n_4465;
wire n_12958;
wire n_12849;
wire n_14849;
wire n_5537;
wire n_5304;
wire n_8524;
wire n_13863;
wire n_13835;
wire n_6059;
wire n_5130;
wire n_12329;
wire n_13650;
wire n_8914;
wire n_10524;
wire n_7520;
wire n_12032;
wire n_12159;
wire n_5162;
wire n_4808;
wire n_8520;
wire n_9490;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_10376;
wire n_12737;
wire n_4482;
wire n_11213;
wire n_10986;
wire n_12504;
wire n_12987;
wire n_14780;
wire n_6267;
wire n_8165;
wire n_11523;
wire n_9525;
wire n_9127;
wire n_9119;
wire n_12521;
wire n_5855;
wire n_11903;
wire n_9002;
wire n_10069;
wire n_10697;
wire n_11100;
wire n_13695;
wire n_12866;
wire n_14030;
wire n_8330;
wire n_12226;
wire n_8682;
wire n_5757;
wire n_6437;
wire n_7331;
wire n_6610;
wire n_7918;
wire n_12170;
wire n_11440;
wire n_10259;
wire n_8467;
wire n_13216;
wire n_8775;
wire n_8886;
wire n_10844;
wire n_12482;
wire n_4926;
wire n_11476;
wire n_8696;
wire n_4116;
wire n_14742;
wire n_6957;
wire n_14658;
wire n_5704;
wire n_7514;
wire n_11966;
wire n_10330;
wire n_7163;
wire n_7620;
wire n_11115;
wire n_9867;
wire n_14089;
wire n_5473;
wire n_11765;
wire n_3754;
wire n_4612;
wire n_5946;
wire n_10197;
wire n_6711;
wire n_14648;
wire n_8464;
wire n_12440;
wire n_4287;
wire n_13313;
wire n_7445;
wire n_10584;
wire n_6847;
wire n_9131;
wire n_9790;
wire n_10522;
wire n_5177;
wire n_11200;
wire n_15011;
wire n_10752;
wire n_11332;
wire n_7123;
wire n_6384;
wire n_10854;
wire n_4516;
wire n_11189;
wire n_12834;
wire n_3794;
wire n_10768;
wire n_14791;
wire n_8720;
wire n_4505;
wire n_14779;
wire n_7959;
wire n_10542;
wire n_9611;
wire n_7563;
wire n_6298;
wire n_11170;
wire n_11337;
wire n_13987;
wire n_9032;
wire n_14218;
wire n_14982;
wire n_9428;
wire n_9990;
wire n_7361;
wire n_12929;
wire n_11278;
wire n_5172;
wire n_4602;
wire n_8186;
wire n_4449;
wire n_9705;
wire n_8890;
wire n_13497;
wire n_7322;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_9774;
wire n_5070;
wire n_14941;
wire n_12022;
wire n_6377;
wire n_12358;
wire n_13793;
wire n_12242;
wire n_4445;
wire n_14010;
wire n_5566;
wire n_10419;
wire n_5414;
wire n_8738;
wire n_13186;
wire n_4870;
wire n_10645;
wire n_11713;
wire n_12214;
wire n_13282;
wire n_13988;
wire n_6348;
wire n_7713;
wire n_10412;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_5450;
wire n_11195;
wire n_6834;
wire n_10124;
wire n_11975;
wire n_5313;
wire n_12254;
wire n_13073;
wire n_13580;
wire n_14178;
wire n_14816;
wire n_12320;
wire n_9374;
wire n_14960;
wire n_4914;
wire n_10737;
wire n_9792;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_14008;
wire n_8066;
wire n_5874;
wire n_14459;
wire n_7977;
wire n_14582;
wire n_14970;
wire n_10294;
wire n_14063;
wire n_10687;
wire n_12763;
wire n_11402;
wire n_14597;
wire n_14976;
wire n_8342;
wire n_13527;
wire n_7508;
wire n_9771;
wire n_10480;
wire n_9712;
wire n_7021;
wire n_13831;
wire n_12627;
wire n_5270;
wire n_11345;
wire n_5956;
wire n_7834;
wire n_14670;
wire n_4345;
wire n_14349;
wire n_5188;
wire n_9905;
wire n_6078;
wire n_7000;
wire n_8571;
wire n_9163;
wire n_9308;
wire n_4318;
wire n_10038;
wire n_10721;
wire n_7921;
wire n_8877;
wire n_4185;
wire n_8862;
wire n_10144;
wire n_8402;
wire n_10410;
wire n_4797;
wire n_7130;
wire n_10823;
wire n_15070;
wire n_10176;
wire n_11714;
wire n_5823;
wire n_3997;
wire n_13687;
wire n_5465;
wire n_4032;
wire n_9387;
wire n_7538;
wire n_11778;
wire n_12492;
wire n_13794;
wire n_7517;
wire n_14948;
wire n_5853;
wire n_14758;
wire n_10799;
wire n_10315;
wire n_7077;
wire n_11300;
wire n_12561;
wire n_14497;
wire n_4343;
wire n_13382;
wire n_11338;
wire n_4212;
wire n_12359;
wire n_6642;
wire n_4124;
wire n_11577;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_10525;
wire n_11930;
wire n_5148;
wire n_4994;
wire n_13353;
wire n_15076;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_11334;
wire n_4378;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_9847;
wire n_12688;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_10932;
wire n_10227;
wire n_11096;
wire n_9577;
wire n_10951;
wire n_4309;
wire n_9111;
wire n_8805;
wire n_10646;
wire n_6511;
wire n_3721;
wire n_12635;
wire n_6507;
wire n_12677;
wire n_14338;
wire n_9513;
wire n_12568;
wire n_11482;
wire n_14819;
wire n_9853;
wire n_11759;
wire n_10710;
wire n_7319;
wire n_7997;
wire n_12610;
wire n_6497;
wire n_12639;
wire n_6001;
wire n_6007;
wire n_9130;
wire n_10409;
wire n_9941;
wire n_9135;
wire n_14414;
wire n_6606;
wire n_4560;
wire n_10709;
wire n_10633;
wire n_5318;
wire n_11829;
wire n_5395;
wire n_14327;
wire n_13901;
wire n_7078;
wire n_7047;
wire n_8144;
wire n_5067;
wire n_3699;
wire n_7107;
wire n_10606;
wire n_13047;
wire n_14077;
wire n_13049;
wire n_3873;
wire n_11936;
wire n_3693;
wire n_10325;
wire n_7469;
wire n_3857;
wire n_13055;
wire n_14786;
wire n_8111;
wire n_11308;

CKINVDCx5p33_ASAP7_75t_R g3632 ( 
.A(n_3237),
.Y(n_3632)
);

BUFx10_ASAP7_75t_L g3633 ( 
.A(n_2243),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_1275),
.Y(n_3634)
);

CKINVDCx5p33_ASAP7_75t_R g3635 ( 
.A(n_3571),
.Y(n_3635)
);

CKINVDCx5p33_ASAP7_75t_R g3636 ( 
.A(n_2970),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3401),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_85),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_625),
.Y(n_3639)
);

CKINVDCx5p33_ASAP7_75t_R g3640 ( 
.A(n_3176),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_2871),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_3195),
.Y(n_3642)
);

CKINVDCx5p33_ASAP7_75t_R g3643 ( 
.A(n_1051),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_132),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_2101),
.Y(n_3645)
);

CKINVDCx5p33_ASAP7_75t_R g3646 ( 
.A(n_789),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_682),
.Y(n_3647)
);

CKINVDCx5p33_ASAP7_75t_R g3648 ( 
.A(n_2559),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_940),
.Y(n_3649)
);

CKINVDCx16_ASAP7_75t_R g3650 ( 
.A(n_3240),
.Y(n_3650)
);

CKINVDCx5p33_ASAP7_75t_R g3651 ( 
.A(n_3120),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_526),
.Y(n_3652)
);

CKINVDCx5p33_ASAP7_75t_R g3653 ( 
.A(n_570),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_380),
.Y(n_3654)
);

CKINVDCx5p33_ASAP7_75t_R g3655 ( 
.A(n_3007),
.Y(n_3655)
);

CKINVDCx5p33_ASAP7_75t_R g3656 ( 
.A(n_3175),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_2518),
.Y(n_3657)
);

BUFx3_ASAP7_75t_L g3658 ( 
.A(n_1276),
.Y(n_3658)
);

CKINVDCx20_ASAP7_75t_R g3659 ( 
.A(n_908),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_2536),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_43),
.Y(n_3661)
);

INVxp67_ASAP7_75t_SL g3662 ( 
.A(n_720),
.Y(n_3662)
);

CKINVDCx5p33_ASAP7_75t_R g3663 ( 
.A(n_2652),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_3192),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3282),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3336),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_1389),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_1089),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_3538),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_1441),
.Y(n_3670)
);

CKINVDCx20_ASAP7_75t_R g3671 ( 
.A(n_62),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_174),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3217),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2851),
.Y(n_3674)
);

CKINVDCx20_ASAP7_75t_R g3675 ( 
.A(n_3261),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_251),
.Y(n_3676)
);

CKINVDCx5p33_ASAP7_75t_R g3677 ( 
.A(n_34),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_1958),
.Y(n_3678)
);

BUFx8_ASAP7_75t_SL g3679 ( 
.A(n_2661),
.Y(n_3679)
);

INVx1_ASAP7_75t_SL g3680 ( 
.A(n_3241),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_1851),
.Y(n_3681)
);

BUFx5_ASAP7_75t_L g3682 ( 
.A(n_3166),
.Y(n_3682)
);

CKINVDCx5p33_ASAP7_75t_R g3683 ( 
.A(n_732),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_66),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3050),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_1289),
.Y(n_3686)
);

INVx1_ASAP7_75t_SL g3687 ( 
.A(n_3450),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_2687),
.Y(n_3688)
);

CKINVDCx5p33_ASAP7_75t_R g3689 ( 
.A(n_3185),
.Y(n_3689)
);

CKINVDCx5p33_ASAP7_75t_R g3690 ( 
.A(n_2764),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_533),
.Y(n_3691)
);

CKINVDCx5p33_ASAP7_75t_R g3692 ( 
.A(n_1133),
.Y(n_3692)
);

CKINVDCx20_ASAP7_75t_R g3693 ( 
.A(n_1303),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3389),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_3179),
.Y(n_3695)
);

CKINVDCx5p33_ASAP7_75t_R g3696 ( 
.A(n_954),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_1344),
.Y(n_3697)
);

BUFx3_ASAP7_75t_L g3698 ( 
.A(n_3533),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_564),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_1887),
.Y(n_3700)
);

CKINVDCx5p33_ASAP7_75t_R g3701 ( 
.A(n_591),
.Y(n_3701)
);

CKINVDCx5p33_ASAP7_75t_R g3702 ( 
.A(n_3272),
.Y(n_3702)
);

CKINVDCx5p33_ASAP7_75t_R g3703 ( 
.A(n_3590),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_2567),
.Y(n_3704)
);

CKINVDCx5p33_ASAP7_75t_R g3705 ( 
.A(n_43),
.Y(n_3705)
);

CKINVDCx5p33_ASAP7_75t_R g3706 ( 
.A(n_83),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_154),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_2914),
.Y(n_3708)
);

CKINVDCx5p33_ASAP7_75t_R g3709 ( 
.A(n_2870),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3549),
.Y(n_3710)
);

INVx3_ASAP7_75t_L g3711 ( 
.A(n_27),
.Y(n_3711)
);

INVx2_ASAP7_75t_SL g3712 ( 
.A(n_1817),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_447),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_2223),
.Y(n_3714)
);

INVx1_ASAP7_75t_SL g3715 ( 
.A(n_2899),
.Y(n_3715)
);

CKINVDCx20_ASAP7_75t_R g3716 ( 
.A(n_652),
.Y(n_3716)
);

CKINVDCx5p33_ASAP7_75t_R g3717 ( 
.A(n_2602),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_801),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_3592),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_1675),
.Y(n_3720)
);

CKINVDCx5p33_ASAP7_75t_R g3721 ( 
.A(n_251),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_1268),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_864),
.Y(n_3723)
);

INVx2_ASAP7_75t_SL g3724 ( 
.A(n_47),
.Y(n_3724)
);

CKINVDCx5p33_ASAP7_75t_R g3725 ( 
.A(n_3034),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3552),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_974),
.Y(n_3727)
);

INVx1_ASAP7_75t_SL g3728 ( 
.A(n_852),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_214),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_505),
.Y(n_3730)
);

CKINVDCx5p33_ASAP7_75t_R g3731 ( 
.A(n_221),
.Y(n_3731)
);

CKINVDCx5p33_ASAP7_75t_R g3732 ( 
.A(n_1772),
.Y(n_3732)
);

INVx1_ASAP7_75t_SL g3733 ( 
.A(n_1715),
.Y(n_3733)
);

CKINVDCx5p33_ASAP7_75t_R g3734 ( 
.A(n_2386),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_597),
.Y(n_3735)
);

CKINVDCx5p33_ASAP7_75t_R g3736 ( 
.A(n_2356),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_2091),
.Y(n_3737)
);

BUFx10_ASAP7_75t_L g3738 ( 
.A(n_1110),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_777),
.Y(n_3739)
);

CKINVDCx16_ASAP7_75t_R g3740 ( 
.A(n_2033),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3329),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_1715),
.Y(n_3742)
);

CKINVDCx5p33_ASAP7_75t_R g3743 ( 
.A(n_1808),
.Y(n_3743)
);

BUFx6f_ASAP7_75t_L g3744 ( 
.A(n_2740),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_482),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3188),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_3245),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_1300),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_3254),
.Y(n_3749)
);

INVx1_ASAP7_75t_SL g3750 ( 
.A(n_3036),
.Y(n_3750)
);

CKINVDCx5p33_ASAP7_75t_R g3751 ( 
.A(n_838),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3224),
.Y(n_3752)
);

CKINVDCx20_ASAP7_75t_R g3753 ( 
.A(n_3200),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_2218),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_3189),
.Y(n_3755)
);

CKINVDCx5p33_ASAP7_75t_R g3756 ( 
.A(n_2838),
.Y(n_3756)
);

CKINVDCx5p33_ASAP7_75t_R g3757 ( 
.A(n_3294),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_1072),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3340),
.Y(n_3759)
);

CKINVDCx20_ASAP7_75t_R g3760 ( 
.A(n_3534),
.Y(n_3760)
);

BUFx2_ASAP7_75t_L g3761 ( 
.A(n_401),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3326),
.Y(n_3762)
);

INVx2_ASAP7_75t_SL g3763 ( 
.A(n_3071),
.Y(n_3763)
);

CKINVDCx5p33_ASAP7_75t_R g3764 ( 
.A(n_51),
.Y(n_3764)
);

CKINVDCx5p33_ASAP7_75t_R g3765 ( 
.A(n_3268),
.Y(n_3765)
);

CKINVDCx5p33_ASAP7_75t_R g3766 ( 
.A(n_3233),
.Y(n_3766)
);

CKINVDCx14_ASAP7_75t_R g3767 ( 
.A(n_284),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_762),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_1377),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_2483),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_3504),
.Y(n_3771)
);

INVx1_ASAP7_75t_SL g3772 ( 
.A(n_2474),
.Y(n_3772)
);

CKINVDCx5p33_ASAP7_75t_R g3773 ( 
.A(n_387),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_843),
.Y(n_3774)
);

CKINVDCx5p33_ASAP7_75t_R g3775 ( 
.A(n_3161),
.Y(n_3775)
);

CKINVDCx5p33_ASAP7_75t_R g3776 ( 
.A(n_3253),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_2819),
.Y(n_3777)
);

CKINVDCx5p33_ASAP7_75t_R g3778 ( 
.A(n_3153),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_2086),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_1155),
.Y(n_3780)
);

CKINVDCx5p33_ASAP7_75t_R g3781 ( 
.A(n_3192),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_3168),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_2502),
.Y(n_3783)
);

CKINVDCx5p33_ASAP7_75t_R g3784 ( 
.A(n_6),
.Y(n_3784)
);

CKINVDCx5p33_ASAP7_75t_R g3785 ( 
.A(n_1237),
.Y(n_3785)
);

CKINVDCx5p33_ASAP7_75t_R g3786 ( 
.A(n_1130),
.Y(n_3786)
);

CKINVDCx5p33_ASAP7_75t_R g3787 ( 
.A(n_1320),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_1163),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_1429),
.Y(n_3789)
);

CKINVDCx5p33_ASAP7_75t_R g3790 ( 
.A(n_21),
.Y(n_3790)
);

CKINVDCx5p33_ASAP7_75t_R g3791 ( 
.A(n_676),
.Y(n_3791)
);

CKINVDCx5p33_ASAP7_75t_R g3792 ( 
.A(n_999),
.Y(n_3792)
);

BUFx3_ASAP7_75t_L g3793 ( 
.A(n_39),
.Y(n_3793)
);

BUFx6f_ASAP7_75t_L g3794 ( 
.A(n_1802),
.Y(n_3794)
);

BUFx10_ASAP7_75t_L g3795 ( 
.A(n_1532),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_1910),
.Y(n_3796)
);

CKINVDCx5p33_ASAP7_75t_R g3797 ( 
.A(n_547),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_2211),
.Y(n_3798)
);

CKINVDCx5p33_ASAP7_75t_R g3799 ( 
.A(n_1095),
.Y(n_3799)
);

CKINVDCx5p33_ASAP7_75t_R g3800 ( 
.A(n_902),
.Y(n_3800)
);

CKINVDCx20_ASAP7_75t_R g3801 ( 
.A(n_1599),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_656),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_1456),
.Y(n_3803)
);

CKINVDCx5p33_ASAP7_75t_R g3804 ( 
.A(n_2892),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3180),
.Y(n_3805)
);

CKINVDCx5p33_ASAP7_75t_R g3806 ( 
.A(n_3480),
.Y(n_3806)
);

CKINVDCx5p33_ASAP7_75t_R g3807 ( 
.A(n_3513),
.Y(n_3807)
);

CKINVDCx5p33_ASAP7_75t_R g3808 ( 
.A(n_3163),
.Y(n_3808)
);

CKINVDCx20_ASAP7_75t_R g3809 ( 
.A(n_2158),
.Y(n_3809)
);

HB1xp67_ASAP7_75t_L g3810 ( 
.A(n_3299),
.Y(n_3810)
);

CKINVDCx5p33_ASAP7_75t_R g3811 ( 
.A(n_1664),
.Y(n_3811)
);

CKINVDCx5p33_ASAP7_75t_R g3812 ( 
.A(n_3382),
.Y(n_3812)
);

CKINVDCx5p33_ASAP7_75t_R g3813 ( 
.A(n_1447),
.Y(n_3813)
);

BUFx6f_ASAP7_75t_L g3814 ( 
.A(n_1618),
.Y(n_3814)
);

BUFx6f_ASAP7_75t_L g3815 ( 
.A(n_2947),
.Y(n_3815)
);

BUFx10_ASAP7_75t_L g3816 ( 
.A(n_3302),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3332),
.Y(n_3817)
);

CKINVDCx20_ASAP7_75t_R g3818 ( 
.A(n_1760),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_396),
.Y(n_3819)
);

CKINVDCx5p33_ASAP7_75t_R g3820 ( 
.A(n_229),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_205),
.Y(n_3821)
);

CKINVDCx5p33_ASAP7_75t_R g3822 ( 
.A(n_1867),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_2173),
.Y(n_3823)
);

CKINVDCx5p33_ASAP7_75t_R g3824 ( 
.A(n_3205),
.Y(n_3824)
);

CKINVDCx16_ASAP7_75t_R g3825 ( 
.A(n_464),
.Y(n_3825)
);

CKINVDCx20_ASAP7_75t_R g3826 ( 
.A(n_656),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_1539),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_956),
.Y(n_3828)
);

CKINVDCx20_ASAP7_75t_R g3829 ( 
.A(n_3346),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_2931),
.Y(n_3830)
);

CKINVDCx5p33_ASAP7_75t_R g3831 ( 
.A(n_195),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3222),
.Y(n_3832)
);

CKINVDCx5p33_ASAP7_75t_R g3833 ( 
.A(n_2419),
.Y(n_3833)
);

CKINVDCx5p33_ASAP7_75t_R g3834 ( 
.A(n_2124),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_2331),
.Y(n_3835)
);

CKINVDCx5p33_ASAP7_75t_R g3836 ( 
.A(n_3221),
.Y(n_3836)
);

CKINVDCx5p33_ASAP7_75t_R g3837 ( 
.A(n_363),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_2852),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3174),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_863),
.Y(n_3840)
);

CKINVDCx5p33_ASAP7_75t_R g3841 ( 
.A(n_3224),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_896),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_296),
.Y(n_3843)
);

BUFx10_ASAP7_75t_L g3844 ( 
.A(n_790),
.Y(n_3844)
);

CKINVDCx5p33_ASAP7_75t_R g3845 ( 
.A(n_2826),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_126),
.Y(n_3846)
);

CKINVDCx5p33_ASAP7_75t_R g3847 ( 
.A(n_2148),
.Y(n_3847)
);

CKINVDCx5p33_ASAP7_75t_R g3848 ( 
.A(n_1742),
.Y(n_3848)
);

CKINVDCx5p33_ASAP7_75t_R g3849 ( 
.A(n_1992),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_2393),
.Y(n_3850)
);

CKINVDCx5p33_ASAP7_75t_R g3851 ( 
.A(n_796),
.Y(n_3851)
);

BUFx6f_ASAP7_75t_L g3852 ( 
.A(n_3186),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_2304),
.Y(n_3853)
);

CKINVDCx20_ASAP7_75t_R g3854 ( 
.A(n_1968),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_1252),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_1003),
.Y(n_3856)
);

CKINVDCx5p33_ASAP7_75t_R g3857 ( 
.A(n_367),
.Y(n_3857)
);

BUFx5_ASAP7_75t_L g3858 ( 
.A(n_343),
.Y(n_3858)
);

INVx1_ASAP7_75t_SL g3859 ( 
.A(n_235),
.Y(n_3859)
);

CKINVDCx20_ASAP7_75t_R g3860 ( 
.A(n_57),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_3196),
.Y(n_3861)
);

CKINVDCx5p33_ASAP7_75t_R g3862 ( 
.A(n_733),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_1102),
.Y(n_3863)
);

CKINVDCx5p33_ASAP7_75t_R g3864 ( 
.A(n_3407),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_1543),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_2480),
.Y(n_3866)
);

CKINVDCx5p33_ASAP7_75t_R g3867 ( 
.A(n_3525),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_2785),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_1127),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_1875),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3596),
.Y(n_3871)
);

CKINVDCx5p33_ASAP7_75t_R g3872 ( 
.A(n_2458),
.Y(n_3872)
);

CKINVDCx5p33_ASAP7_75t_R g3873 ( 
.A(n_2829),
.Y(n_3873)
);

CKINVDCx5p33_ASAP7_75t_R g3874 ( 
.A(n_3227),
.Y(n_3874)
);

CKINVDCx5p33_ASAP7_75t_R g3875 ( 
.A(n_77),
.Y(n_3875)
);

CKINVDCx5p33_ASAP7_75t_R g3876 ( 
.A(n_3220),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_2517),
.Y(n_3877)
);

CKINVDCx5p33_ASAP7_75t_R g3878 ( 
.A(n_203),
.Y(n_3878)
);

CKINVDCx5p33_ASAP7_75t_R g3879 ( 
.A(n_777),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_1117),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3443),
.Y(n_3881)
);

CKINVDCx5p33_ASAP7_75t_R g3882 ( 
.A(n_1458),
.Y(n_3882)
);

CKINVDCx20_ASAP7_75t_R g3883 ( 
.A(n_1290),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_2871),
.Y(n_3884)
);

CKINVDCx5p33_ASAP7_75t_R g3885 ( 
.A(n_93),
.Y(n_3885)
);

CKINVDCx5p33_ASAP7_75t_R g3886 ( 
.A(n_3609),
.Y(n_3886)
);

CKINVDCx5p33_ASAP7_75t_R g3887 ( 
.A(n_2021),
.Y(n_3887)
);

CKINVDCx16_ASAP7_75t_R g3888 ( 
.A(n_330),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_2788),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_441),
.Y(n_3890)
);

CKINVDCx16_ASAP7_75t_R g3891 ( 
.A(n_3629),
.Y(n_3891)
);

CKINVDCx5p33_ASAP7_75t_R g3892 ( 
.A(n_1786),
.Y(n_3892)
);

CKINVDCx5p33_ASAP7_75t_R g3893 ( 
.A(n_2108),
.Y(n_3893)
);

CKINVDCx5p33_ASAP7_75t_R g3894 ( 
.A(n_1667),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3582),
.Y(n_3895)
);

CKINVDCx5p33_ASAP7_75t_R g3896 ( 
.A(n_2956),
.Y(n_3896)
);

CKINVDCx5p33_ASAP7_75t_R g3897 ( 
.A(n_93),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_1662),
.Y(n_3898)
);

CKINVDCx5p33_ASAP7_75t_R g3899 ( 
.A(n_1756),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3088),
.Y(n_3900)
);

CKINVDCx5p33_ASAP7_75t_R g3901 ( 
.A(n_3128),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_141),
.Y(n_3902)
);

BUFx3_ASAP7_75t_L g3903 ( 
.A(n_984),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_1634),
.Y(n_3904)
);

CKINVDCx5p33_ASAP7_75t_R g3905 ( 
.A(n_1383),
.Y(n_3905)
);

CKINVDCx5p33_ASAP7_75t_R g3906 ( 
.A(n_3275),
.Y(n_3906)
);

CKINVDCx5p33_ASAP7_75t_R g3907 ( 
.A(n_2634),
.Y(n_3907)
);

BUFx2_ASAP7_75t_L g3908 ( 
.A(n_2698),
.Y(n_3908)
);

CKINVDCx5p33_ASAP7_75t_R g3909 ( 
.A(n_2840),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3403),
.Y(n_3910)
);

CKINVDCx5p33_ASAP7_75t_R g3911 ( 
.A(n_3243),
.Y(n_3911)
);

BUFx10_ASAP7_75t_L g3912 ( 
.A(n_2743),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3259),
.Y(n_3913)
);

BUFx10_ASAP7_75t_L g3914 ( 
.A(n_2309),
.Y(n_3914)
);

CKINVDCx20_ASAP7_75t_R g3915 ( 
.A(n_2335),
.Y(n_3915)
);

CKINVDCx5p33_ASAP7_75t_R g3916 ( 
.A(n_3385),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_2340),
.Y(n_3917)
);

CKINVDCx5p33_ASAP7_75t_R g3918 ( 
.A(n_2979),
.Y(n_3918)
);

BUFx6f_ASAP7_75t_L g3919 ( 
.A(n_2741),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_2439),
.Y(n_3920)
);

CKINVDCx5p33_ASAP7_75t_R g3921 ( 
.A(n_3215),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_178),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_151),
.Y(n_3923)
);

INVx2_ASAP7_75t_SL g3924 ( 
.A(n_2140),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_287),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_2955),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3208),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_1038),
.Y(n_3928)
);

INVx1_ASAP7_75t_SL g3929 ( 
.A(n_710),
.Y(n_3929)
);

CKINVDCx5p33_ASAP7_75t_R g3930 ( 
.A(n_2547),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_2091),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_1678),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3541),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_762),
.Y(n_3934)
);

CKINVDCx16_ASAP7_75t_R g3935 ( 
.A(n_225),
.Y(n_3935)
);

BUFx6f_ASAP7_75t_L g3936 ( 
.A(n_408),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_1788),
.Y(n_3937)
);

HB1xp67_ASAP7_75t_L g3938 ( 
.A(n_1883),
.Y(n_3938)
);

CKINVDCx5p33_ASAP7_75t_R g3939 ( 
.A(n_3476),
.Y(n_3939)
);

BUFx3_ASAP7_75t_L g3940 ( 
.A(n_2018),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3457),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_2025),
.Y(n_3942)
);

CKINVDCx5p33_ASAP7_75t_R g3943 ( 
.A(n_1107),
.Y(n_3943)
);

CKINVDCx5p33_ASAP7_75t_R g3944 ( 
.A(n_1181),
.Y(n_3944)
);

CKINVDCx5p33_ASAP7_75t_R g3945 ( 
.A(n_1362),
.Y(n_3945)
);

INVx1_ASAP7_75t_SL g3946 ( 
.A(n_3194),
.Y(n_3946)
);

CKINVDCx5p33_ASAP7_75t_R g3947 ( 
.A(n_331),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_2087),
.Y(n_3948)
);

CKINVDCx20_ASAP7_75t_R g3949 ( 
.A(n_1862),
.Y(n_3949)
);

CKINVDCx16_ASAP7_75t_R g3950 ( 
.A(n_2213),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_816),
.Y(n_3951)
);

CKINVDCx14_ASAP7_75t_R g3952 ( 
.A(n_692),
.Y(n_3952)
);

CKINVDCx5p33_ASAP7_75t_R g3953 ( 
.A(n_2200),
.Y(n_3953)
);

BUFx10_ASAP7_75t_L g3954 ( 
.A(n_2703),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_1423),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_314),
.Y(n_3956)
);

CKINVDCx20_ASAP7_75t_R g3957 ( 
.A(n_3467),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3246),
.Y(n_3958)
);

CKINVDCx5p33_ASAP7_75t_R g3959 ( 
.A(n_119),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_1141),
.Y(n_3960)
);

CKINVDCx5p33_ASAP7_75t_R g3961 ( 
.A(n_1187),
.Y(n_3961)
);

BUFx6f_ASAP7_75t_L g3962 ( 
.A(n_3133),
.Y(n_3962)
);

CKINVDCx5p33_ASAP7_75t_R g3963 ( 
.A(n_182),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_1253),
.Y(n_3964)
);

INVx2_ASAP7_75t_SL g3965 ( 
.A(n_2666),
.Y(n_3965)
);

HB1xp67_ASAP7_75t_L g3966 ( 
.A(n_2367),
.Y(n_3966)
);

BUFx6f_ASAP7_75t_L g3967 ( 
.A(n_482),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_2135),
.Y(n_3968)
);

CKINVDCx20_ASAP7_75t_R g3969 ( 
.A(n_514),
.Y(n_3969)
);

CKINVDCx5p33_ASAP7_75t_R g3970 ( 
.A(n_485),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_1290),
.Y(n_3971)
);

BUFx3_ASAP7_75t_L g3972 ( 
.A(n_2770),
.Y(n_3972)
);

CKINVDCx5p33_ASAP7_75t_R g3973 ( 
.A(n_185),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3041),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3102),
.Y(n_3975)
);

CKINVDCx5p33_ASAP7_75t_R g3976 ( 
.A(n_867),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3232),
.Y(n_3977)
);

CKINVDCx20_ASAP7_75t_R g3978 ( 
.A(n_2400),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_3349),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_2388),
.Y(n_3980)
);

CKINVDCx5p33_ASAP7_75t_R g3981 ( 
.A(n_1628),
.Y(n_3981)
);

CKINVDCx5p33_ASAP7_75t_R g3982 ( 
.A(n_1575),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_1251),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3324),
.Y(n_3984)
);

CKINVDCx20_ASAP7_75t_R g3985 ( 
.A(n_2714),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3307),
.Y(n_3986)
);

BUFx10_ASAP7_75t_L g3987 ( 
.A(n_118),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_1434),
.Y(n_3988)
);

CKINVDCx5p33_ASAP7_75t_R g3989 ( 
.A(n_1351),
.Y(n_3989)
);

INVx2_ASAP7_75t_SL g3990 ( 
.A(n_3296),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_1368),
.Y(n_3991)
);

INVx1_ASAP7_75t_SL g3992 ( 
.A(n_1947),
.Y(n_3992)
);

INVx1_ASAP7_75t_SL g3993 ( 
.A(n_2966),
.Y(n_3993)
);

CKINVDCx20_ASAP7_75t_R g3994 ( 
.A(n_347),
.Y(n_3994)
);

CKINVDCx5p33_ASAP7_75t_R g3995 ( 
.A(n_3021),
.Y(n_3995)
);

CKINVDCx5p33_ASAP7_75t_R g3996 ( 
.A(n_609),
.Y(n_3996)
);

CKINVDCx20_ASAP7_75t_R g3997 ( 
.A(n_1852),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_1210),
.Y(n_3998)
);

CKINVDCx5p33_ASAP7_75t_R g3999 ( 
.A(n_2680),
.Y(n_3999)
);

CKINVDCx5p33_ASAP7_75t_R g4000 ( 
.A(n_1291),
.Y(n_4000)
);

BUFx10_ASAP7_75t_L g4001 ( 
.A(n_2570),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_1771),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_2747),
.Y(n_4003)
);

CKINVDCx5p33_ASAP7_75t_R g4004 ( 
.A(n_2823),
.Y(n_4004)
);

CKINVDCx5p33_ASAP7_75t_R g4005 ( 
.A(n_2890),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_2368),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_3308),
.Y(n_4007)
);

CKINVDCx5p33_ASAP7_75t_R g4008 ( 
.A(n_1448),
.Y(n_4008)
);

BUFx6f_ASAP7_75t_L g4009 ( 
.A(n_2982),
.Y(n_4009)
);

CKINVDCx5p33_ASAP7_75t_R g4010 ( 
.A(n_3190),
.Y(n_4010)
);

CKINVDCx14_ASAP7_75t_R g4011 ( 
.A(n_1831),
.Y(n_4011)
);

CKINVDCx5p33_ASAP7_75t_R g4012 ( 
.A(n_3583),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_1179),
.Y(n_4013)
);

CKINVDCx5p33_ASAP7_75t_R g4014 ( 
.A(n_3512),
.Y(n_4014)
);

CKINVDCx5p33_ASAP7_75t_R g4015 ( 
.A(n_2487),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_906),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_1247),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_717),
.Y(n_4018)
);

BUFx5_ASAP7_75t_L g4019 ( 
.A(n_1344),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_198),
.Y(n_4020)
);

CKINVDCx5p33_ASAP7_75t_R g4021 ( 
.A(n_2509),
.Y(n_4021)
);

CKINVDCx5p33_ASAP7_75t_R g4022 ( 
.A(n_2471),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3070),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_201),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_2516),
.Y(n_4025)
);

CKINVDCx20_ASAP7_75t_R g4026 ( 
.A(n_12),
.Y(n_4026)
);

INVx2_ASAP7_75t_SL g4027 ( 
.A(n_934),
.Y(n_4027)
);

BUFx2_ASAP7_75t_L g4028 ( 
.A(n_2514),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_2743),
.Y(n_4029)
);

CKINVDCx5p33_ASAP7_75t_R g4030 ( 
.A(n_3198),
.Y(n_4030)
);

BUFx2_ASAP7_75t_L g4031 ( 
.A(n_1080),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3074),
.Y(n_4032)
);

CKINVDCx5p33_ASAP7_75t_R g4033 ( 
.A(n_2976),
.Y(n_4033)
);

CKINVDCx5p33_ASAP7_75t_R g4034 ( 
.A(n_2250),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_926),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_340),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_421),
.Y(n_4037)
);

INVxp67_ASAP7_75t_L g4038 ( 
.A(n_1826),
.Y(n_4038)
);

CKINVDCx5p33_ASAP7_75t_R g4039 ( 
.A(n_3134),
.Y(n_4039)
);

CKINVDCx5p33_ASAP7_75t_R g4040 ( 
.A(n_1130),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_3561),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_1759),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_740),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_469),
.Y(n_4044)
);

CKINVDCx5p33_ASAP7_75t_R g4045 ( 
.A(n_1528),
.Y(n_4045)
);

CKINVDCx5p33_ASAP7_75t_R g4046 ( 
.A(n_763),
.Y(n_4046)
);

CKINVDCx5p33_ASAP7_75t_R g4047 ( 
.A(n_3238),
.Y(n_4047)
);

CKINVDCx5p33_ASAP7_75t_R g4048 ( 
.A(n_1858),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_1998),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_1291),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_2810),
.Y(n_4051)
);

CKINVDCx5p33_ASAP7_75t_R g4052 ( 
.A(n_1490),
.Y(n_4052)
);

BUFx6f_ASAP7_75t_L g4053 ( 
.A(n_791),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_1493),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_2778),
.Y(n_4055)
);

CKINVDCx5p33_ASAP7_75t_R g4056 ( 
.A(n_167),
.Y(n_4056)
);

CKINVDCx20_ASAP7_75t_R g4057 ( 
.A(n_1984),
.Y(n_4057)
);

CKINVDCx5p33_ASAP7_75t_R g4058 ( 
.A(n_3164),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_1265),
.Y(n_4059)
);

INVx1_ASAP7_75t_SL g4060 ( 
.A(n_1840),
.Y(n_4060)
);

CKINVDCx5p33_ASAP7_75t_R g4061 ( 
.A(n_3390),
.Y(n_4061)
);

CKINVDCx20_ASAP7_75t_R g4062 ( 
.A(n_3319),
.Y(n_4062)
);

CKINVDCx5p33_ASAP7_75t_R g4063 ( 
.A(n_3328),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_1337),
.Y(n_4064)
);

INVx1_ASAP7_75t_SL g4065 ( 
.A(n_3286),
.Y(n_4065)
);

INVxp33_ASAP7_75t_L g4066 ( 
.A(n_3140),
.Y(n_4066)
);

CKINVDCx5p33_ASAP7_75t_R g4067 ( 
.A(n_382),
.Y(n_4067)
);

CKINVDCx5p33_ASAP7_75t_R g4068 ( 
.A(n_3153),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_782),
.Y(n_4069)
);

CKINVDCx5p33_ASAP7_75t_R g4070 ( 
.A(n_2111),
.Y(n_4070)
);

CKINVDCx5p33_ASAP7_75t_R g4071 ( 
.A(n_3271),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_2737),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_2586),
.Y(n_4073)
);

CKINVDCx5p33_ASAP7_75t_R g4074 ( 
.A(n_1662),
.Y(n_4074)
);

CKINVDCx5p33_ASAP7_75t_R g4075 ( 
.A(n_2270),
.Y(n_4075)
);

CKINVDCx5p33_ASAP7_75t_R g4076 ( 
.A(n_1120),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_702),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_3242),
.Y(n_4078)
);

CKINVDCx16_ASAP7_75t_R g4079 ( 
.A(n_96),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_162),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_452),
.Y(n_4081)
);

BUFx3_ASAP7_75t_L g4082 ( 
.A(n_1644),
.Y(n_4082)
);

CKINVDCx5p33_ASAP7_75t_R g4083 ( 
.A(n_1726),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3262),
.Y(n_4084)
);

CKINVDCx5p33_ASAP7_75t_R g4085 ( 
.A(n_3444),
.Y(n_4085)
);

CKINVDCx5p33_ASAP7_75t_R g4086 ( 
.A(n_907),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_188),
.Y(n_4087)
);

CKINVDCx5p33_ASAP7_75t_R g4088 ( 
.A(n_2293),
.Y(n_4088)
);

CKINVDCx5p33_ASAP7_75t_R g4089 ( 
.A(n_381),
.Y(n_4089)
);

INVx2_ASAP7_75t_SL g4090 ( 
.A(n_908),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_3199),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_1617),
.Y(n_4092)
);

CKINVDCx5p33_ASAP7_75t_R g4093 ( 
.A(n_70),
.Y(n_4093)
);

CKINVDCx5p33_ASAP7_75t_R g4094 ( 
.A(n_1798),
.Y(n_4094)
);

CKINVDCx5p33_ASAP7_75t_R g4095 ( 
.A(n_2780),
.Y(n_4095)
);

CKINVDCx5p33_ASAP7_75t_R g4096 ( 
.A(n_805),
.Y(n_4096)
);

CKINVDCx5p33_ASAP7_75t_R g4097 ( 
.A(n_3472),
.Y(n_4097)
);

CKINVDCx5p33_ASAP7_75t_R g4098 ( 
.A(n_785),
.Y(n_4098)
);

CKINVDCx5p33_ASAP7_75t_R g4099 ( 
.A(n_1678),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3258),
.Y(n_4100)
);

HB1xp67_ASAP7_75t_L g4101 ( 
.A(n_496),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3234),
.Y(n_4102)
);

CKINVDCx5p33_ASAP7_75t_R g4103 ( 
.A(n_1813),
.Y(n_4103)
);

CKINVDCx5p33_ASAP7_75t_R g4104 ( 
.A(n_127),
.Y(n_4104)
);

CKINVDCx5p33_ASAP7_75t_R g4105 ( 
.A(n_2394),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_1655),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3091),
.Y(n_4107)
);

CKINVDCx5p33_ASAP7_75t_R g4108 ( 
.A(n_3263),
.Y(n_4108)
);

BUFx2_ASAP7_75t_L g4109 ( 
.A(n_2762),
.Y(n_4109)
);

BUFx3_ASAP7_75t_L g4110 ( 
.A(n_1197),
.Y(n_4110)
);

CKINVDCx5p33_ASAP7_75t_R g4111 ( 
.A(n_3523),
.Y(n_4111)
);

CKINVDCx5p33_ASAP7_75t_R g4112 ( 
.A(n_2628),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_331),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_1270),
.Y(n_4114)
);

CKINVDCx20_ASAP7_75t_R g4115 ( 
.A(n_3316),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_585),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_1365),
.Y(n_4117)
);

CKINVDCx5p33_ASAP7_75t_R g4118 ( 
.A(n_3558),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_1537),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_531),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3438),
.Y(n_4121)
);

CKINVDCx5p33_ASAP7_75t_R g4122 ( 
.A(n_593),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3344),
.Y(n_4123)
);

CKINVDCx5p33_ASAP7_75t_R g4124 ( 
.A(n_1967),
.Y(n_4124)
);

CKINVDCx5p33_ASAP7_75t_R g4125 ( 
.A(n_2411),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_1302),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_3286),
.Y(n_4127)
);

CKINVDCx5p33_ASAP7_75t_R g4128 ( 
.A(n_1555),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_395),
.Y(n_4129)
);

CKINVDCx16_ASAP7_75t_R g4130 ( 
.A(n_2682),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_192),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_232),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3442),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_67),
.Y(n_4134)
);

INVx2_ASAP7_75t_SL g4135 ( 
.A(n_310),
.Y(n_4135)
);

INVx2_ASAP7_75t_R g4136 ( 
.A(n_3249),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_629),
.Y(n_4137)
);

CKINVDCx5p33_ASAP7_75t_R g4138 ( 
.A(n_502),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_58),
.Y(n_4139)
);

BUFx6f_ASAP7_75t_L g4140 ( 
.A(n_2810),
.Y(n_4140)
);

INVx2_ASAP7_75t_SL g4141 ( 
.A(n_3317),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_2208),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_1029),
.Y(n_4143)
);

CKINVDCx5p33_ASAP7_75t_R g4144 ( 
.A(n_1508),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_3267),
.Y(n_4145)
);

CKINVDCx5p33_ASAP7_75t_R g4146 ( 
.A(n_1956),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_2833),
.Y(n_4147)
);

CKINVDCx5p33_ASAP7_75t_R g4148 ( 
.A(n_3312),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_1245),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_1020),
.Y(n_4150)
);

CKINVDCx5p33_ASAP7_75t_R g4151 ( 
.A(n_3372),
.Y(n_4151)
);

CKINVDCx5p33_ASAP7_75t_R g4152 ( 
.A(n_3445),
.Y(n_4152)
);

BUFx6f_ASAP7_75t_L g4153 ( 
.A(n_2917),
.Y(n_4153)
);

HB1xp67_ASAP7_75t_L g4154 ( 
.A(n_3231),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_214),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_3234),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_1985),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_206),
.Y(n_4158)
);

CKINVDCx5p33_ASAP7_75t_R g4159 ( 
.A(n_1289),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3330),
.Y(n_4160)
);

CKINVDCx5p33_ASAP7_75t_R g4161 ( 
.A(n_3201),
.Y(n_4161)
);

CKINVDCx5p33_ASAP7_75t_R g4162 ( 
.A(n_516),
.Y(n_4162)
);

BUFx3_ASAP7_75t_L g4163 ( 
.A(n_798),
.Y(n_4163)
);

INVx1_ASAP7_75t_SL g4164 ( 
.A(n_2233),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_1893),
.Y(n_4165)
);

CKINVDCx5p33_ASAP7_75t_R g4166 ( 
.A(n_3200),
.Y(n_4166)
);

INVxp67_ASAP7_75t_L g4167 ( 
.A(n_262),
.Y(n_4167)
);

CKINVDCx5p33_ASAP7_75t_R g4168 ( 
.A(n_284),
.Y(n_4168)
);

BUFx3_ASAP7_75t_L g4169 ( 
.A(n_3335),
.Y(n_4169)
);

CKINVDCx20_ASAP7_75t_R g4170 ( 
.A(n_3515),
.Y(n_4170)
);

CKINVDCx5p33_ASAP7_75t_R g4171 ( 
.A(n_92),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3247),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_2486),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_2934),
.Y(n_4174)
);

CKINVDCx5p33_ASAP7_75t_R g4175 ( 
.A(n_2227),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_1593),
.Y(n_4176)
);

CKINVDCx5p33_ASAP7_75t_R g4177 ( 
.A(n_3197),
.Y(n_4177)
);

CKINVDCx5p33_ASAP7_75t_R g4178 ( 
.A(n_2275),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_3271),
.Y(n_4179)
);

CKINVDCx5p33_ASAP7_75t_R g4180 ( 
.A(n_1418),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_2476),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3278),
.Y(n_4182)
);

BUFx6f_ASAP7_75t_L g4183 ( 
.A(n_118),
.Y(n_4183)
);

CKINVDCx5p33_ASAP7_75t_R g4184 ( 
.A(n_1972),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3581),
.Y(n_4185)
);

CKINVDCx5p33_ASAP7_75t_R g4186 ( 
.A(n_434),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_184),
.Y(n_4187)
);

CKINVDCx5p33_ASAP7_75t_R g4188 ( 
.A(n_3279),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_2218),
.Y(n_4189)
);

INVx1_ASAP7_75t_SL g4190 ( 
.A(n_27),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_253),
.Y(n_4191)
);

BUFx5_ASAP7_75t_L g4192 ( 
.A(n_456),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_1696),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_3280),
.Y(n_4194)
);

CKINVDCx20_ASAP7_75t_R g4195 ( 
.A(n_2650),
.Y(n_4195)
);

CKINVDCx5p33_ASAP7_75t_R g4196 ( 
.A(n_3102),
.Y(n_4196)
);

BUFx8_ASAP7_75t_SL g4197 ( 
.A(n_2907),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_359),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_413),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3434),
.Y(n_4200)
);

CKINVDCx5p33_ASAP7_75t_R g4201 ( 
.A(n_3284),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_265),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_1869),
.Y(n_4203)
);

CKINVDCx5p33_ASAP7_75t_R g4204 ( 
.A(n_2566),
.Y(n_4204)
);

INVxp67_ASAP7_75t_L g4205 ( 
.A(n_584),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_1362),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3171),
.Y(n_4207)
);

CKINVDCx5p33_ASAP7_75t_R g4208 ( 
.A(n_502),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_1443),
.Y(n_4209)
);

BUFx6f_ASAP7_75t_L g4210 ( 
.A(n_2894),
.Y(n_4210)
);

CKINVDCx5p33_ASAP7_75t_R g4211 ( 
.A(n_1041),
.Y(n_4211)
);

BUFx10_ASAP7_75t_L g4212 ( 
.A(n_2309),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_2440),
.Y(n_4213)
);

CKINVDCx5p33_ASAP7_75t_R g4214 ( 
.A(n_891),
.Y(n_4214)
);

CKINVDCx20_ASAP7_75t_R g4215 ( 
.A(n_2316),
.Y(n_4215)
);

CKINVDCx16_ASAP7_75t_R g4216 ( 
.A(n_783),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_2434),
.Y(n_4217)
);

CKINVDCx20_ASAP7_75t_R g4218 ( 
.A(n_3388),
.Y(n_4218)
);

CKINVDCx5p33_ASAP7_75t_R g4219 ( 
.A(n_589),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3243),
.Y(n_4220)
);

INVxp67_ASAP7_75t_L g4221 ( 
.A(n_3554),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_2527),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_1538),
.Y(n_4223)
);

CKINVDCx5p33_ASAP7_75t_R g4224 ( 
.A(n_3398),
.Y(n_4224)
);

CKINVDCx5p33_ASAP7_75t_R g4225 ( 
.A(n_1992),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_2688),
.Y(n_4226)
);

CKINVDCx5p33_ASAP7_75t_R g4227 ( 
.A(n_3187),
.Y(n_4227)
);

CKINVDCx14_ASAP7_75t_R g4228 ( 
.A(n_1028),
.Y(n_4228)
);

CKINVDCx5p33_ASAP7_75t_R g4229 ( 
.A(n_3236),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_1443),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_2012),
.Y(n_4231)
);

CKINVDCx5p33_ASAP7_75t_R g4232 ( 
.A(n_2163),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_551),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_3430),
.Y(n_4234)
);

CKINVDCx16_ASAP7_75t_R g4235 ( 
.A(n_1396),
.Y(n_4235)
);

CKINVDCx20_ASAP7_75t_R g4236 ( 
.A(n_2114),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_370),
.Y(n_4237)
);

CKINVDCx5p33_ASAP7_75t_R g4238 ( 
.A(n_3257),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_878),
.Y(n_4239)
);

CKINVDCx5p33_ASAP7_75t_R g4240 ( 
.A(n_1071),
.Y(n_4240)
);

CKINVDCx5p33_ASAP7_75t_R g4241 ( 
.A(n_2306),
.Y(n_4241)
);

BUFx10_ASAP7_75t_L g4242 ( 
.A(n_1684),
.Y(n_4242)
);

CKINVDCx20_ASAP7_75t_R g4243 ( 
.A(n_2713),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_3313),
.Y(n_4244)
);

CKINVDCx5p33_ASAP7_75t_R g4245 ( 
.A(n_869),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_26),
.Y(n_4246)
);

HB1xp67_ASAP7_75t_L g4247 ( 
.A(n_3155),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_2998),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_1088),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_488),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_2834),
.Y(n_4251)
);

CKINVDCx5p33_ASAP7_75t_R g4252 ( 
.A(n_2954),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_3551),
.Y(n_4253)
);

CKINVDCx16_ASAP7_75t_R g4254 ( 
.A(n_2183),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3613),
.Y(n_4255)
);

CKINVDCx5p33_ASAP7_75t_R g4256 ( 
.A(n_3165),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_1949),
.Y(n_4257)
);

CKINVDCx5p33_ASAP7_75t_R g4258 ( 
.A(n_2147),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_1852),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_1814),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_2114),
.Y(n_4261)
);

CKINVDCx5p33_ASAP7_75t_R g4262 ( 
.A(n_3325),
.Y(n_4262)
);

CKINVDCx16_ASAP7_75t_R g4263 ( 
.A(n_3068),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_1086),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_3449),
.Y(n_4265)
);

CKINVDCx5p33_ASAP7_75t_R g4266 ( 
.A(n_1231),
.Y(n_4266)
);

CKINVDCx5p33_ASAP7_75t_R g4267 ( 
.A(n_2145),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_3101),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_2620),
.Y(n_4269)
);

CKINVDCx5p33_ASAP7_75t_R g4270 ( 
.A(n_494),
.Y(n_4270)
);

CKINVDCx5p33_ASAP7_75t_R g4271 ( 
.A(n_2673),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_2044),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_2989),
.Y(n_4273)
);

CKINVDCx5p33_ASAP7_75t_R g4274 ( 
.A(n_2041),
.Y(n_4274)
);

CKINVDCx20_ASAP7_75t_R g4275 ( 
.A(n_770),
.Y(n_4275)
);

CKINVDCx5p33_ASAP7_75t_R g4276 ( 
.A(n_3441),
.Y(n_4276)
);

CKINVDCx5p33_ASAP7_75t_R g4277 ( 
.A(n_918),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_1531),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_2348),
.Y(n_4279)
);

CKINVDCx5p33_ASAP7_75t_R g4280 ( 
.A(n_1263),
.Y(n_4280)
);

CKINVDCx5p33_ASAP7_75t_R g4281 ( 
.A(n_172),
.Y(n_4281)
);

CKINVDCx5p33_ASAP7_75t_R g4282 ( 
.A(n_3006),
.Y(n_4282)
);

CKINVDCx5p33_ASAP7_75t_R g4283 ( 
.A(n_2599),
.Y(n_4283)
);

CKINVDCx5p33_ASAP7_75t_R g4284 ( 
.A(n_3129),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_841),
.Y(n_4285)
);

CKINVDCx5p33_ASAP7_75t_R g4286 ( 
.A(n_3157),
.Y(n_4286)
);

CKINVDCx5p33_ASAP7_75t_R g4287 ( 
.A(n_1580),
.Y(n_4287)
);

CKINVDCx5p33_ASAP7_75t_R g4288 ( 
.A(n_2517),
.Y(n_4288)
);

CKINVDCx20_ASAP7_75t_R g4289 ( 
.A(n_2060),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_3340),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3281),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_2769),
.Y(n_4292)
);

CKINVDCx5p33_ASAP7_75t_R g4293 ( 
.A(n_1326),
.Y(n_4293)
);

CKINVDCx5p33_ASAP7_75t_R g4294 ( 
.A(n_3331),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_2147),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_790),
.Y(n_4296)
);

CKINVDCx20_ASAP7_75t_R g4297 ( 
.A(n_798),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_1230),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_42),
.Y(n_4299)
);

CKINVDCx5p33_ASAP7_75t_R g4300 ( 
.A(n_860),
.Y(n_4300)
);

CKINVDCx5p33_ASAP7_75t_R g4301 ( 
.A(n_3173),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_2469),
.Y(n_4302)
);

CKINVDCx5p33_ASAP7_75t_R g4303 ( 
.A(n_2999),
.Y(n_4303)
);

CKINVDCx5p33_ASAP7_75t_R g4304 ( 
.A(n_3341),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_1457),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_1779),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_3540),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_2023),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_734),
.Y(n_4309)
);

CKINVDCx5p33_ASAP7_75t_R g4310 ( 
.A(n_1643),
.Y(n_4310)
);

CKINVDCx20_ASAP7_75t_R g4311 ( 
.A(n_3381),
.Y(n_4311)
);

CKINVDCx5p33_ASAP7_75t_R g4312 ( 
.A(n_1568),
.Y(n_4312)
);

CKINVDCx5p33_ASAP7_75t_R g4313 ( 
.A(n_2578),
.Y(n_4313)
);

CKINVDCx5p33_ASAP7_75t_R g4314 ( 
.A(n_3212),
.Y(n_4314)
);

INVx2_ASAP7_75t_SL g4315 ( 
.A(n_2970),
.Y(n_4315)
);

CKINVDCx5p33_ASAP7_75t_R g4316 ( 
.A(n_116),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_1577),
.Y(n_4317)
);

CKINVDCx5p33_ASAP7_75t_R g4318 ( 
.A(n_2207),
.Y(n_4318)
);

CKINVDCx5p33_ASAP7_75t_R g4319 ( 
.A(n_1007),
.Y(n_4319)
);

CKINVDCx5p33_ASAP7_75t_R g4320 ( 
.A(n_2436),
.Y(n_4320)
);

CKINVDCx5p33_ASAP7_75t_R g4321 ( 
.A(n_3293),
.Y(n_4321)
);

CKINVDCx20_ASAP7_75t_R g4322 ( 
.A(n_1870),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_1077),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_367),
.Y(n_4324)
);

CKINVDCx5p33_ASAP7_75t_R g4325 ( 
.A(n_2132),
.Y(n_4325)
);

BUFx6f_ASAP7_75t_L g4326 ( 
.A(n_3061),
.Y(n_4326)
);

CKINVDCx5p33_ASAP7_75t_R g4327 ( 
.A(n_2930),
.Y(n_4327)
);

BUFx6f_ASAP7_75t_L g4328 ( 
.A(n_1341),
.Y(n_4328)
);

CKINVDCx5p33_ASAP7_75t_R g4329 ( 
.A(n_2838),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3219),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_2655),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_286),
.Y(n_4332)
);

INVxp67_ASAP7_75t_L g4333 ( 
.A(n_616),
.Y(n_4333)
);

BUFx3_ASAP7_75t_L g4334 ( 
.A(n_712),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_3208),
.Y(n_4335)
);

CKINVDCx5p33_ASAP7_75t_R g4336 ( 
.A(n_3615),
.Y(n_4336)
);

CKINVDCx5p33_ASAP7_75t_R g4337 ( 
.A(n_3248),
.Y(n_4337)
);

CKINVDCx5p33_ASAP7_75t_R g4338 ( 
.A(n_3318),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_2812),
.Y(n_4339)
);

BUFx3_ASAP7_75t_L g4340 ( 
.A(n_2734),
.Y(n_4340)
);

CKINVDCx5p33_ASAP7_75t_R g4341 ( 
.A(n_976),
.Y(n_4341)
);

CKINVDCx20_ASAP7_75t_R g4342 ( 
.A(n_2464),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_3501),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_3210),
.Y(n_4344)
);

BUFx6f_ASAP7_75t_L g4345 ( 
.A(n_3338),
.Y(n_4345)
);

CKINVDCx5p33_ASAP7_75t_R g4346 ( 
.A(n_3178),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_2051),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_1211),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_968),
.Y(n_4349)
);

CKINVDCx5p33_ASAP7_75t_R g4350 ( 
.A(n_109),
.Y(n_4350)
);

BUFx3_ASAP7_75t_L g4351 ( 
.A(n_1223),
.Y(n_4351)
);

CKINVDCx5p33_ASAP7_75t_R g4352 ( 
.A(n_2004),
.Y(n_4352)
);

CKINVDCx5p33_ASAP7_75t_R g4353 ( 
.A(n_2947),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_764),
.Y(n_4354)
);

CKINVDCx20_ASAP7_75t_R g4355 ( 
.A(n_3321),
.Y(n_4355)
);

BUFx3_ASAP7_75t_L g4356 ( 
.A(n_34),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_3376),
.Y(n_4357)
);

BUFx6f_ASAP7_75t_L g4358 ( 
.A(n_296),
.Y(n_4358)
);

BUFx3_ASAP7_75t_L g4359 ( 
.A(n_2819),
.Y(n_4359)
);

CKINVDCx20_ASAP7_75t_R g4360 ( 
.A(n_1321),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3207),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_1871),
.Y(n_4362)
);

CKINVDCx5p33_ASAP7_75t_R g4363 ( 
.A(n_3121),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_3202),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_2103),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_3339),
.Y(n_4366)
);

CKINVDCx5p33_ASAP7_75t_R g4367 ( 
.A(n_1707),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_2960),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_172),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_3556),
.Y(n_4370)
);

INVx2_ASAP7_75t_SL g4371 ( 
.A(n_1082),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_1398),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_2429),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_1901),
.Y(n_4374)
);

CKINVDCx5p33_ASAP7_75t_R g4375 ( 
.A(n_2041),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_590),
.Y(n_4376)
);

BUFx8_ASAP7_75t_SL g4377 ( 
.A(n_1280),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_55),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_1419),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_942),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_1739),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_1580),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_2149),
.Y(n_4383)
);

CKINVDCx5p33_ASAP7_75t_R g4384 ( 
.A(n_800),
.Y(n_4384)
);

CKINVDCx5p33_ASAP7_75t_R g4385 ( 
.A(n_3507),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_1158),
.Y(n_4386)
);

BUFx3_ASAP7_75t_L g4387 ( 
.A(n_693),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_1922),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_2956),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_2258),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_3297),
.Y(n_4391)
);

BUFx6f_ASAP7_75t_L g4392 ( 
.A(n_3266),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_350),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_2323),
.Y(n_4394)
);

CKINVDCx5p33_ASAP7_75t_R g4395 ( 
.A(n_1721),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_2839),
.Y(n_4396)
);

CKINVDCx20_ASAP7_75t_R g4397 ( 
.A(n_2730),
.Y(n_4397)
);

CKINVDCx5p33_ASAP7_75t_R g4398 ( 
.A(n_701),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_2796),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_3170),
.Y(n_4400)
);

BUFx6f_ASAP7_75t_L g4401 ( 
.A(n_3323),
.Y(n_4401)
);

CKINVDCx5p33_ASAP7_75t_R g4402 ( 
.A(n_1522),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_2051),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_1186),
.Y(n_4404)
);

CKINVDCx5p33_ASAP7_75t_R g4405 ( 
.A(n_932),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_851),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_2832),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_984),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_2573),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_1295),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_1695),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_2456),
.Y(n_4412)
);

BUFx6f_ASAP7_75t_L g4413 ( 
.A(n_1618),
.Y(n_4413)
);

CKINVDCx5p33_ASAP7_75t_R g4414 ( 
.A(n_22),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_1411),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_909),
.Y(n_4416)
);

CKINVDCx5p33_ASAP7_75t_R g4417 ( 
.A(n_1321),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_3037),
.Y(n_4418)
);

INVx1_ASAP7_75t_SL g4419 ( 
.A(n_991),
.Y(n_4419)
);

CKINVDCx5p33_ASAP7_75t_R g4420 ( 
.A(n_3252),
.Y(n_4420)
);

CKINVDCx16_ASAP7_75t_R g4421 ( 
.A(n_3235),
.Y(n_4421)
);

CKINVDCx5p33_ASAP7_75t_R g4422 ( 
.A(n_3573),
.Y(n_4422)
);

CKINVDCx5p33_ASAP7_75t_R g4423 ( 
.A(n_1498),
.Y(n_4423)
);

CKINVDCx5p33_ASAP7_75t_R g4424 ( 
.A(n_1770),
.Y(n_4424)
);

CKINVDCx5p33_ASAP7_75t_R g4425 ( 
.A(n_1970),
.Y(n_4425)
);

CKINVDCx5p33_ASAP7_75t_R g4426 ( 
.A(n_1918),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_1500),
.Y(n_4427)
);

CKINVDCx5p33_ASAP7_75t_R g4428 ( 
.A(n_3211),
.Y(n_4428)
);

CKINVDCx5p33_ASAP7_75t_R g4429 ( 
.A(n_445),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_2848),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_2462),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_1460),
.Y(n_4432)
);

CKINVDCx20_ASAP7_75t_R g4433 ( 
.A(n_1259),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_3075),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_975),
.Y(n_4435)
);

BUFx3_ASAP7_75t_L g4436 ( 
.A(n_430),
.Y(n_4436)
);

CKINVDCx5p33_ASAP7_75t_R g4437 ( 
.A(n_3163),
.Y(n_4437)
);

CKINVDCx5p33_ASAP7_75t_R g4438 ( 
.A(n_3300),
.Y(n_4438)
);

CKINVDCx5p33_ASAP7_75t_R g4439 ( 
.A(n_3436),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3038),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3458),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_3396),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_2805),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_783),
.Y(n_4444)
);

CKINVDCx5p33_ASAP7_75t_R g4445 ( 
.A(n_88),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_1380),
.Y(n_4446)
);

INVx1_ASAP7_75t_SL g4447 ( 
.A(n_2881),
.Y(n_4447)
);

BUFx3_ASAP7_75t_L g4448 ( 
.A(n_1569),
.Y(n_4448)
);

CKINVDCx16_ASAP7_75t_R g4449 ( 
.A(n_3327),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_1326),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_397),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_2488),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_1071),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_818),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_89),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_687),
.Y(n_4456)
);

CKINVDCx5p33_ASAP7_75t_R g4457 ( 
.A(n_2583),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_2299),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_1259),
.Y(n_4459)
);

CKINVDCx5p33_ASAP7_75t_R g4460 ( 
.A(n_1980),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_3272),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_2207),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_2100),
.Y(n_4463)
);

BUFx10_ASAP7_75t_L g4464 ( 
.A(n_944),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_352),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_2945),
.Y(n_4466)
);

CKINVDCx5p33_ASAP7_75t_R g4467 ( 
.A(n_1522),
.Y(n_4467)
);

CKINVDCx5p33_ASAP7_75t_R g4468 ( 
.A(n_350),
.Y(n_4468)
);

CKINVDCx20_ASAP7_75t_R g4469 ( 
.A(n_2477),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_3255),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_1517),
.Y(n_4471)
);

BUFx8_ASAP7_75t_SL g4472 ( 
.A(n_2285),
.Y(n_4472)
);

INVx1_ASAP7_75t_SL g4473 ( 
.A(n_1031),
.Y(n_4473)
);

BUFx10_ASAP7_75t_L g4474 ( 
.A(n_443),
.Y(n_4474)
);

CKINVDCx20_ASAP7_75t_R g4475 ( 
.A(n_497),
.Y(n_4475)
);

CKINVDCx5p33_ASAP7_75t_R g4476 ( 
.A(n_2791),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_2313),
.Y(n_4477)
);

CKINVDCx5p33_ASAP7_75t_R g4478 ( 
.A(n_3363),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_1103),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_1225),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_2131),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_865),
.Y(n_4482)
);

CKINVDCx5p33_ASAP7_75t_R g4483 ( 
.A(n_3248),
.Y(n_4483)
);

BUFx10_ASAP7_75t_L g4484 ( 
.A(n_254),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_2893),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_560),
.Y(n_4486)
);

CKINVDCx20_ASAP7_75t_R g4487 ( 
.A(n_351),
.Y(n_4487)
);

CKINVDCx5p33_ASAP7_75t_R g4488 ( 
.A(n_3049),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_2548),
.Y(n_4489)
);

HB1xp67_ASAP7_75t_L g4490 ( 
.A(n_75),
.Y(n_4490)
);

INVx1_ASAP7_75t_SL g4491 ( 
.A(n_3580),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_622),
.Y(n_4492)
);

CKINVDCx5p33_ASAP7_75t_R g4493 ( 
.A(n_2085),
.Y(n_4493)
);

CKINVDCx5p33_ASAP7_75t_R g4494 ( 
.A(n_200),
.Y(n_4494)
);

CKINVDCx5p33_ASAP7_75t_R g4495 ( 
.A(n_2400),
.Y(n_4495)
);

CKINVDCx5p33_ASAP7_75t_R g4496 ( 
.A(n_1125),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_2894),
.Y(n_4497)
);

CKINVDCx5p33_ASAP7_75t_R g4498 ( 
.A(n_2523),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_1986),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_3329),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_3256),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_3386),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_1830),
.Y(n_4503)
);

CKINVDCx14_ASAP7_75t_R g4504 ( 
.A(n_3132),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_949),
.Y(n_4505)
);

CKINVDCx5p33_ASAP7_75t_R g4506 ( 
.A(n_2140),
.Y(n_4506)
);

CKINVDCx5p33_ASAP7_75t_R g4507 ( 
.A(n_1542),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_876),
.Y(n_4508)
);

CKINVDCx5p33_ASAP7_75t_R g4509 ( 
.A(n_1788),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_1037),
.Y(n_4510)
);

CKINVDCx5p33_ASAP7_75t_R g4511 ( 
.A(n_2390),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_3425),
.Y(n_4512)
);

CKINVDCx5p33_ASAP7_75t_R g4513 ( 
.A(n_1155),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_3152),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_1894),
.Y(n_4515)
);

CKINVDCx5p33_ASAP7_75t_R g4516 ( 
.A(n_1324),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_3260),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_769),
.Y(n_4518)
);

CKINVDCx5p33_ASAP7_75t_R g4519 ( 
.A(n_386),
.Y(n_4519)
);

CKINVDCx5p33_ASAP7_75t_R g4520 ( 
.A(n_2110),
.Y(n_4520)
);

CKINVDCx5p33_ASAP7_75t_R g4521 ( 
.A(n_2337),
.Y(n_4521)
);

CKINVDCx5p33_ASAP7_75t_R g4522 ( 
.A(n_1663),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_581),
.Y(n_4523)
);

INVx2_ASAP7_75t_SL g4524 ( 
.A(n_2502),
.Y(n_4524)
);

CKINVDCx5p33_ASAP7_75t_R g4525 ( 
.A(n_810),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3229),
.Y(n_4526)
);

CKINVDCx5p33_ASAP7_75t_R g4527 ( 
.A(n_3219),
.Y(n_4527)
);

BUFx10_ASAP7_75t_L g4528 ( 
.A(n_2375),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_94),
.Y(n_4529)
);

CKINVDCx5p33_ASAP7_75t_R g4530 ( 
.A(n_2043),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_2821),
.Y(n_4531)
);

CKINVDCx5p33_ASAP7_75t_R g4532 ( 
.A(n_3223),
.Y(n_4532)
);

BUFx2_ASAP7_75t_SL g4533 ( 
.A(n_1122),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_1755),
.Y(n_4534)
);

CKINVDCx20_ASAP7_75t_R g4535 ( 
.A(n_2700),
.Y(n_4535)
);

CKINVDCx16_ASAP7_75t_R g4536 ( 
.A(n_3462),
.Y(n_4536)
);

CKINVDCx5p33_ASAP7_75t_R g4537 ( 
.A(n_3246),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_602),
.Y(n_4538)
);

BUFx10_ASAP7_75t_L g4539 ( 
.A(n_1967),
.Y(n_4539)
);

CKINVDCx5p33_ASAP7_75t_R g4540 ( 
.A(n_440),
.Y(n_4540)
);

INVx1_ASAP7_75t_SL g4541 ( 
.A(n_2128),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_1860),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_2513),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3250),
.Y(n_4544)
);

INVx1_ASAP7_75t_SL g4545 ( 
.A(n_2337),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_2307),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_3289),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_3260),
.Y(n_4548)
);

CKINVDCx5p33_ASAP7_75t_R g4549 ( 
.A(n_2370),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_252),
.Y(n_4550)
);

CKINVDCx5p33_ASAP7_75t_R g4551 ( 
.A(n_2606),
.Y(n_4551)
);

CKINVDCx20_ASAP7_75t_R g4552 ( 
.A(n_59),
.Y(n_4552)
);

CKINVDCx5p33_ASAP7_75t_R g4553 ( 
.A(n_2297),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_3290),
.Y(n_4554)
);

CKINVDCx5p33_ASAP7_75t_R g4555 ( 
.A(n_2100),
.Y(n_4555)
);

BUFx2_ASAP7_75t_L g4556 ( 
.A(n_3191),
.Y(n_4556)
);

CKINVDCx5p33_ASAP7_75t_R g4557 ( 
.A(n_3451),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_1971),
.Y(n_4558)
);

CKINVDCx5p33_ASAP7_75t_R g4559 ( 
.A(n_2048),
.Y(n_4559)
);

CKINVDCx20_ASAP7_75t_R g4560 ( 
.A(n_749),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_668),
.Y(n_4561)
);

CKINVDCx20_ASAP7_75t_R g4562 ( 
.A(n_1803),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_697),
.Y(n_4563)
);

CKINVDCx5p33_ASAP7_75t_R g4564 ( 
.A(n_1537),
.Y(n_4564)
);

CKINVDCx20_ASAP7_75t_R g4565 ( 
.A(n_2526),
.Y(n_4565)
);

CKINVDCx5p33_ASAP7_75t_R g4566 ( 
.A(n_2402),
.Y(n_4566)
);

CKINVDCx5p33_ASAP7_75t_R g4567 ( 
.A(n_3363),
.Y(n_4567)
);

CKINVDCx5p33_ASAP7_75t_R g4568 ( 
.A(n_1945),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_3162),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_1240),
.Y(n_4570)
);

CKINVDCx20_ASAP7_75t_R g4571 ( 
.A(n_1342),
.Y(n_4571)
);

CKINVDCx5p33_ASAP7_75t_R g4572 ( 
.A(n_2520),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_2519),
.Y(n_4573)
);

INVx1_ASAP7_75t_SL g4574 ( 
.A(n_1294),
.Y(n_4574)
);

CKINVDCx5p33_ASAP7_75t_R g4575 ( 
.A(n_1270),
.Y(n_4575)
);

CKINVDCx5p33_ASAP7_75t_R g4576 ( 
.A(n_456),
.Y(n_4576)
);

CKINVDCx5p33_ASAP7_75t_R g4577 ( 
.A(n_3043),
.Y(n_4577)
);

CKINVDCx20_ASAP7_75t_R g4578 ( 
.A(n_2886),
.Y(n_4578)
);

CKINVDCx5p33_ASAP7_75t_R g4579 ( 
.A(n_2054),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_3484),
.Y(n_4580)
);

CKINVDCx5p33_ASAP7_75t_R g4581 ( 
.A(n_40),
.Y(n_4581)
);

CKINVDCx5p33_ASAP7_75t_R g4582 ( 
.A(n_2781),
.Y(n_4582)
);

CKINVDCx5p33_ASAP7_75t_R g4583 ( 
.A(n_3226),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_2130),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_1417),
.Y(n_4585)
);

CKINVDCx20_ASAP7_75t_R g4586 ( 
.A(n_3343),
.Y(n_4586)
);

INVx1_ASAP7_75t_SL g4587 ( 
.A(n_1506),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_1116),
.Y(n_4588)
);

CKINVDCx20_ASAP7_75t_R g4589 ( 
.A(n_3085),
.Y(n_4589)
);

CKINVDCx5p33_ASAP7_75t_R g4590 ( 
.A(n_739),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_3628),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_2995),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_2759),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_3245),
.Y(n_4594)
);

CKINVDCx5p33_ASAP7_75t_R g4595 ( 
.A(n_1885),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_2099),
.Y(n_4596)
);

INVxp67_ASAP7_75t_SL g4597 ( 
.A(n_990),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_1284),
.Y(n_4598)
);

CKINVDCx5p33_ASAP7_75t_R g4599 ( 
.A(n_2127),
.Y(n_4599)
);

CKINVDCx16_ASAP7_75t_R g4600 ( 
.A(n_935),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_1021),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_347),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_3314),
.Y(n_4603)
);

CKINVDCx5p33_ASAP7_75t_R g4604 ( 
.A(n_493),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_302),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_574),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_1660),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_586),
.Y(n_4608)
);

CKINVDCx20_ASAP7_75t_R g4609 ( 
.A(n_835),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_3232),
.Y(n_4610)
);

CKINVDCx16_ASAP7_75t_R g4611 ( 
.A(n_243),
.Y(n_4611)
);

BUFx10_ASAP7_75t_L g4612 ( 
.A(n_920),
.Y(n_4612)
);

CKINVDCx5p33_ASAP7_75t_R g4613 ( 
.A(n_2449),
.Y(n_4613)
);

CKINVDCx5p33_ASAP7_75t_R g4614 ( 
.A(n_1926),
.Y(n_4614)
);

CKINVDCx5p33_ASAP7_75t_R g4615 ( 
.A(n_1780),
.Y(n_4615)
);

INVxp67_ASAP7_75t_L g4616 ( 
.A(n_538),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_57),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_3320),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_2475),
.Y(n_4619)
);

INVx1_ASAP7_75t_SL g4620 ( 
.A(n_3557),
.Y(n_4620)
);

CKINVDCx20_ASAP7_75t_R g4621 ( 
.A(n_2307),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_1379),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_147),
.Y(n_4623)
);

CKINVDCx5p33_ASAP7_75t_R g4624 ( 
.A(n_2317),
.Y(n_4624)
);

CKINVDCx5p33_ASAP7_75t_R g4625 ( 
.A(n_14),
.Y(n_4625)
);

BUFx5_ASAP7_75t_L g4626 ( 
.A(n_572),
.Y(n_4626)
);

INVx2_ASAP7_75t_SL g4627 ( 
.A(n_903),
.Y(n_4627)
);

CKINVDCx5p33_ASAP7_75t_R g4628 ( 
.A(n_361),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_2228),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_1248),
.Y(n_4630)
);

INVx1_ASAP7_75t_SL g4631 ( 
.A(n_1633),
.Y(n_4631)
);

CKINVDCx5p33_ASAP7_75t_R g4632 ( 
.A(n_178),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_2733),
.Y(n_4633)
);

CKINVDCx5p33_ASAP7_75t_R g4634 ( 
.A(n_745),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_3181),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_2235),
.Y(n_4636)
);

BUFx6f_ASAP7_75t_L g4637 ( 
.A(n_1472),
.Y(n_4637)
);

CKINVDCx5p33_ASAP7_75t_R g4638 ( 
.A(n_3303),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_3218),
.Y(n_4639)
);

CKINVDCx5p33_ASAP7_75t_R g4640 ( 
.A(n_3239),
.Y(n_4640)
);

INVxp67_ASAP7_75t_L g4641 ( 
.A(n_2335),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_557),
.Y(n_4642)
);

CKINVDCx5p33_ASAP7_75t_R g4643 ( 
.A(n_860),
.Y(n_4643)
);

CKINVDCx5p33_ASAP7_75t_R g4644 ( 
.A(n_2470),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_242),
.Y(n_4645)
);

CKINVDCx5p33_ASAP7_75t_R g4646 ( 
.A(n_3334),
.Y(n_4646)
);

INVx1_ASAP7_75t_SL g4647 ( 
.A(n_909),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_1277),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_3321),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_1288),
.Y(n_4650)
);

CKINVDCx5p33_ASAP7_75t_R g4651 ( 
.A(n_1948),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_3287),
.Y(n_4652)
);

BUFx2_ASAP7_75t_SL g4653 ( 
.A(n_736),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_584),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_395),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_1884),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_144),
.Y(n_4657)
);

CKINVDCx5p33_ASAP7_75t_R g4658 ( 
.A(n_797),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_190),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_2728),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_3553),
.Y(n_4661)
);

INVx1_ASAP7_75t_SL g4662 ( 
.A(n_165),
.Y(n_4662)
);

INVx2_ASAP7_75t_SL g4663 ( 
.A(n_1380),
.Y(n_4663)
);

CKINVDCx5p33_ASAP7_75t_R g4664 ( 
.A(n_3274),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_2462),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_2389),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_3175),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_3010),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_1844),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_1432),
.Y(n_4670)
);

INVx1_ASAP7_75t_SL g4671 ( 
.A(n_993),
.Y(n_4671)
);

CKINVDCx5p33_ASAP7_75t_R g4672 ( 
.A(n_1553),
.Y(n_4672)
);

INVx1_ASAP7_75t_SL g4673 ( 
.A(n_1869),
.Y(n_4673)
);

CKINVDCx5p33_ASAP7_75t_R g4674 ( 
.A(n_3367),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_737),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_782),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_1221),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_1413),
.Y(n_4678)
);

CKINVDCx5p33_ASAP7_75t_R g4679 ( 
.A(n_144),
.Y(n_4679)
);

HB1xp67_ASAP7_75t_L g4680 ( 
.A(n_358),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_2060),
.Y(n_4681)
);

BUFx6f_ASAP7_75t_L g4682 ( 
.A(n_2825),
.Y(n_4682)
);

BUFx2_ASAP7_75t_L g4683 ( 
.A(n_217),
.Y(n_4683)
);

CKINVDCx5p33_ASAP7_75t_R g4684 ( 
.A(n_848),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_2864),
.Y(n_4685)
);

CKINVDCx5p33_ASAP7_75t_R g4686 ( 
.A(n_3298),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_2272),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_3374),
.Y(n_4688)
);

CKINVDCx5p33_ASAP7_75t_R g4689 ( 
.A(n_1329),
.Y(n_4689)
);

CKINVDCx5p33_ASAP7_75t_R g4690 ( 
.A(n_1273),
.Y(n_4690)
);

CKINVDCx5p33_ASAP7_75t_R g4691 ( 
.A(n_1529),
.Y(n_4691)
);

CKINVDCx5p33_ASAP7_75t_R g4692 ( 
.A(n_2000),
.Y(n_4692)
);

CKINVDCx5p33_ASAP7_75t_R g4693 ( 
.A(n_3311),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_3203),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_3358),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_2043),
.Y(n_4696)
);

CKINVDCx5p33_ASAP7_75t_R g4697 ( 
.A(n_564),
.Y(n_4697)
);

CKINVDCx5p33_ASAP7_75t_R g4698 ( 
.A(n_290),
.Y(n_4698)
);

INVx2_ASAP7_75t_L g4699 ( 
.A(n_2635),
.Y(n_4699)
);

CKINVDCx5p33_ASAP7_75t_R g4700 ( 
.A(n_3038),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_195),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_567),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_494),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_2116),
.Y(n_4704)
);

CKINVDCx5p33_ASAP7_75t_R g4705 ( 
.A(n_679),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_2157),
.Y(n_4706)
);

CKINVDCx5p33_ASAP7_75t_R g4707 ( 
.A(n_348),
.Y(n_4707)
);

CKINVDCx5p33_ASAP7_75t_R g4708 ( 
.A(n_183),
.Y(n_4708)
);

CKINVDCx20_ASAP7_75t_R g4709 ( 
.A(n_3265),
.Y(n_4709)
);

CKINVDCx16_ASAP7_75t_R g4710 ( 
.A(n_3345),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_249),
.Y(n_4711)
);

CKINVDCx5p33_ASAP7_75t_R g4712 ( 
.A(n_3301),
.Y(n_4712)
);

CKINVDCx5p33_ASAP7_75t_R g4713 ( 
.A(n_2454),
.Y(n_4713)
);

CKINVDCx5p33_ASAP7_75t_R g4714 ( 
.A(n_2712),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_438),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_1724),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_1278),
.Y(n_4717)
);

BUFx3_ASAP7_75t_L g4718 ( 
.A(n_3520),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_3251),
.Y(n_4719)
);

CKINVDCx5p33_ASAP7_75t_R g4720 ( 
.A(n_2171),
.Y(n_4720)
);

CKINVDCx5p33_ASAP7_75t_R g4721 ( 
.A(n_1350),
.Y(n_4721)
);

CKINVDCx5p33_ASAP7_75t_R g4722 ( 
.A(n_474),
.Y(n_4722)
);

CKINVDCx16_ASAP7_75t_R g4723 ( 
.A(n_1266),
.Y(n_4723)
);

BUFx10_ASAP7_75t_L g4724 ( 
.A(n_3295),
.Y(n_4724)
);

CKINVDCx5p33_ASAP7_75t_R g4725 ( 
.A(n_3228),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_1469),
.Y(n_4726)
);

BUFx6f_ASAP7_75t_L g4727 ( 
.A(n_1460),
.Y(n_4727)
);

CKINVDCx5p33_ASAP7_75t_R g4728 ( 
.A(n_1409),
.Y(n_4728)
);

CKINVDCx5p33_ASAP7_75t_R g4729 ( 
.A(n_2001),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_3263),
.Y(n_4730)
);

CKINVDCx5p33_ASAP7_75t_R g4731 ( 
.A(n_3309),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_757),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_2643),
.Y(n_4733)
);

CKINVDCx20_ASAP7_75t_R g4734 ( 
.A(n_3206),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_1709),
.Y(n_4735)
);

CKINVDCx5p33_ASAP7_75t_R g4736 ( 
.A(n_524),
.Y(n_4736)
);

CKINVDCx5p33_ASAP7_75t_R g4737 ( 
.A(n_1184),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_1097),
.Y(n_4738)
);

CKINVDCx5p33_ASAP7_75t_R g4739 ( 
.A(n_954),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_2391),
.Y(n_4740)
);

CKINVDCx5p33_ASAP7_75t_R g4741 ( 
.A(n_2492),
.Y(n_4741)
);

CKINVDCx5p33_ASAP7_75t_R g4742 ( 
.A(n_3306),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_107),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_2363),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_560),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_2391),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_3118),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_129),
.Y(n_4748)
);

CKINVDCx5p33_ASAP7_75t_R g4749 ( 
.A(n_1833),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_87),
.Y(n_4750)
);

INVxp67_ASAP7_75t_L g4751 ( 
.A(n_3305),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_1738),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_861),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_1795),
.Y(n_4754)
);

CKINVDCx5p33_ASAP7_75t_R g4755 ( 
.A(n_2407),
.Y(n_4755)
);

CKINVDCx5p33_ASAP7_75t_R g4756 ( 
.A(n_3622),
.Y(n_4756)
);

BUFx6f_ASAP7_75t_L g4757 ( 
.A(n_1387),
.Y(n_4757)
);

CKINVDCx20_ASAP7_75t_R g4758 ( 
.A(n_963),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_1374),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_1184),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_2209),
.Y(n_4761)
);

CKINVDCx5p33_ASAP7_75t_R g4762 ( 
.A(n_2625),
.Y(n_4762)
);

BUFx2_ASAP7_75t_L g4763 ( 
.A(n_1466),
.Y(n_4763)
);

CKINVDCx20_ASAP7_75t_R g4764 ( 
.A(n_2389),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_981),
.Y(n_4765)
);

INVx2_ASAP7_75t_SL g4766 ( 
.A(n_3207),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_448),
.Y(n_4767)
);

CKINVDCx5p33_ASAP7_75t_R g4768 ( 
.A(n_3264),
.Y(n_4768)
);

CKINVDCx5p33_ASAP7_75t_R g4769 ( 
.A(n_2594),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_1004),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_1772),
.Y(n_4771)
);

CKINVDCx5p33_ASAP7_75t_R g4772 ( 
.A(n_3314),
.Y(n_4772)
);

CKINVDCx5p33_ASAP7_75t_R g4773 ( 
.A(n_1761),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_1604),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_3167),
.Y(n_4775)
);

CKINVDCx20_ASAP7_75t_R g4776 ( 
.A(n_1458),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_2697),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_375),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_3347),
.Y(n_4779)
);

CKINVDCx20_ASAP7_75t_R g4780 ( 
.A(n_1622),
.Y(n_4780)
);

BUFx6f_ASAP7_75t_L g4781 ( 
.A(n_2369),
.Y(n_4781)
);

CKINVDCx5p33_ASAP7_75t_R g4782 ( 
.A(n_323),
.Y(n_4782)
);

BUFx2_ASAP7_75t_L g4783 ( 
.A(n_3315),
.Y(n_4783)
);

BUFx10_ASAP7_75t_L g4784 ( 
.A(n_3322),
.Y(n_4784)
);

BUFx3_ASAP7_75t_L g4785 ( 
.A(n_2704),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_711),
.Y(n_4786)
);

CKINVDCx5p33_ASAP7_75t_R g4787 ( 
.A(n_1669),
.Y(n_4787)
);

CKINVDCx5p33_ASAP7_75t_R g4788 ( 
.A(n_1816),
.Y(n_4788)
);

CKINVDCx5p33_ASAP7_75t_R g4789 ( 
.A(n_2710),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_3177),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_2406),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_1529),
.Y(n_4792)
);

CKINVDCx5p33_ASAP7_75t_R g4793 ( 
.A(n_2440),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_1402),
.Y(n_4794)
);

CKINVDCx5p33_ASAP7_75t_R g4795 ( 
.A(n_3),
.Y(n_4795)
);

CKINVDCx5p33_ASAP7_75t_R g4796 ( 
.A(n_1301),
.Y(n_4796)
);

CKINVDCx5p33_ASAP7_75t_R g4797 ( 
.A(n_753),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_3214),
.Y(n_4798)
);

CKINVDCx5p33_ASAP7_75t_R g4799 ( 
.A(n_2990),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_3506),
.Y(n_4800)
);

INVxp67_ASAP7_75t_SL g4801 ( 
.A(n_2177),
.Y(n_4801)
);

BUFx3_ASAP7_75t_L g4802 ( 
.A(n_3115),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_3216),
.Y(n_4803)
);

BUFx3_ASAP7_75t_L g4804 ( 
.A(n_1069),
.Y(n_4804)
);

CKINVDCx5p33_ASAP7_75t_R g4805 ( 
.A(n_1174),
.Y(n_4805)
);

BUFx10_ASAP7_75t_L g4806 ( 
.A(n_2196),
.Y(n_4806)
);

CKINVDCx5p33_ASAP7_75t_R g4807 ( 
.A(n_499),
.Y(n_4807)
);

CKINVDCx5p33_ASAP7_75t_R g4808 ( 
.A(n_3231),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_3285),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_1338),
.Y(n_4810)
);

CKINVDCx5p33_ASAP7_75t_R g4811 ( 
.A(n_2889),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_2129),
.Y(n_4812)
);

CKINVDCx5p33_ASAP7_75t_R g4813 ( 
.A(n_520),
.Y(n_4813)
);

CKINVDCx5p33_ASAP7_75t_R g4814 ( 
.A(n_3182),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_2694),
.Y(n_4815)
);

CKINVDCx5p33_ASAP7_75t_R g4816 ( 
.A(n_3276),
.Y(n_4816)
);

INVxp67_ASAP7_75t_L g4817 ( 
.A(n_2664),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_3333),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_1338),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_1608),
.Y(n_4820)
);

CKINVDCx5p33_ASAP7_75t_R g4821 ( 
.A(n_1666),
.Y(n_4821)
);

CKINVDCx5p33_ASAP7_75t_R g4822 ( 
.A(n_1667),
.Y(n_4822)
);

CKINVDCx20_ASAP7_75t_R g4823 ( 
.A(n_3225),
.Y(n_4823)
);

CKINVDCx5p33_ASAP7_75t_R g4824 ( 
.A(n_3112),
.Y(n_4824)
);

CKINVDCx5p33_ASAP7_75t_R g4825 ( 
.A(n_3186),
.Y(n_4825)
);

INVx1_ASAP7_75t_SL g4826 ( 
.A(n_503),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_3337),
.Y(n_4827)
);

CKINVDCx5p33_ASAP7_75t_R g4828 ( 
.A(n_1246),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_167),
.Y(n_4829)
);

CKINVDCx5p33_ASAP7_75t_R g4830 ( 
.A(n_1944),
.Y(n_4830)
);

CKINVDCx5p33_ASAP7_75t_R g4831 ( 
.A(n_3183),
.Y(n_4831)
);

CKINVDCx5p33_ASAP7_75t_R g4832 ( 
.A(n_821),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_1795),
.Y(n_4833)
);

CKINVDCx5p33_ASAP7_75t_R g4834 ( 
.A(n_2467),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_437),
.Y(n_4835)
);

BUFx2_ASAP7_75t_L g4836 ( 
.A(n_3310),
.Y(n_4836)
);

CKINVDCx5p33_ASAP7_75t_R g4837 ( 
.A(n_1164),
.Y(n_4837)
);

CKINVDCx5p33_ASAP7_75t_R g4838 ( 
.A(n_2407),
.Y(n_4838)
);

CKINVDCx20_ASAP7_75t_R g4839 ( 
.A(n_368),
.Y(n_4839)
);

BUFx6f_ASAP7_75t_L g4840 ( 
.A(n_292),
.Y(n_4840)
);

CKINVDCx5p33_ASAP7_75t_R g4841 ( 
.A(n_69),
.Y(n_4841)
);

CKINVDCx5p33_ASAP7_75t_R g4842 ( 
.A(n_3319),
.Y(n_4842)
);

BUFx2_ASAP7_75t_R g4843 ( 
.A(n_1444),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_1243),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_3070),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_1091),
.Y(n_4846)
);

BUFx3_ASAP7_75t_L g4847 ( 
.A(n_1668),
.Y(n_4847)
);

CKINVDCx20_ASAP7_75t_R g4848 ( 
.A(n_1447),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_586),
.Y(n_4849)
);

CKINVDCx5p33_ASAP7_75t_R g4850 ( 
.A(n_2392),
.Y(n_4850)
);

INVxp67_ASAP7_75t_L g4851 ( 
.A(n_676),
.Y(n_4851)
);

BUFx3_ASAP7_75t_L g4852 ( 
.A(n_2682),
.Y(n_4852)
);

CKINVDCx5p33_ASAP7_75t_R g4853 ( 
.A(n_2500),
.Y(n_4853)
);

BUFx3_ASAP7_75t_L g4854 ( 
.A(n_3599),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_3193),
.Y(n_4855)
);

CKINVDCx5p33_ASAP7_75t_R g4856 ( 
.A(n_2102),
.Y(n_4856)
);

CKINVDCx5p33_ASAP7_75t_R g4857 ( 
.A(n_977),
.Y(n_4857)
);

CKINVDCx5p33_ASAP7_75t_R g4858 ( 
.A(n_2519),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_1858),
.Y(n_4859)
);

CKINVDCx20_ASAP7_75t_R g4860 ( 
.A(n_1150),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_940),
.Y(n_4861)
);

CKINVDCx5p33_ASAP7_75t_R g4862 ( 
.A(n_2786),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_3045),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_713),
.Y(n_4864)
);

CKINVDCx5p33_ASAP7_75t_R g4865 ( 
.A(n_2843),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_2496),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_3169),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_749),
.Y(n_4868)
);

INVx1_ASAP7_75t_SL g4869 ( 
.A(n_3288),
.Y(n_4869)
);

CKINVDCx5p33_ASAP7_75t_R g4870 ( 
.A(n_1730),
.Y(n_4870)
);

CKINVDCx20_ASAP7_75t_R g4871 ( 
.A(n_3043),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_3209),
.Y(n_4872)
);

CKINVDCx5p33_ASAP7_75t_R g4873 ( 
.A(n_1901),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_1167),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_3526),
.Y(n_4875)
);

CKINVDCx5p33_ASAP7_75t_R g4876 ( 
.A(n_1261),
.Y(n_4876)
);

CKINVDCx16_ASAP7_75t_R g4877 ( 
.A(n_1018),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_3292),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_1845),
.Y(n_4879)
);

CKINVDCx20_ASAP7_75t_R g4880 ( 
.A(n_594),
.Y(n_4880)
);

CKINVDCx5p33_ASAP7_75t_R g4881 ( 
.A(n_3460),
.Y(n_4881)
);

CKINVDCx5p33_ASAP7_75t_R g4882 ( 
.A(n_3334),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_1904),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_606),
.Y(n_4884)
);

CKINVDCx5p33_ASAP7_75t_R g4885 ( 
.A(n_2195),
.Y(n_4885)
);

CKINVDCx5p33_ASAP7_75t_R g4886 ( 
.A(n_2873),
.Y(n_4886)
);

INVxp67_ASAP7_75t_L g4887 ( 
.A(n_2055),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_2909),
.Y(n_4888)
);

CKINVDCx5p33_ASAP7_75t_R g4889 ( 
.A(n_3269),
.Y(n_4889)
);

CKINVDCx20_ASAP7_75t_R g4890 ( 
.A(n_3221),
.Y(n_4890)
);

CKINVDCx5p33_ASAP7_75t_R g4891 ( 
.A(n_3537),
.Y(n_4891)
);

CKINVDCx20_ASAP7_75t_R g4892 ( 
.A(n_768),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_558),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_1382),
.Y(n_4894)
);

CKINVDCx20_ASAP7_75t_R g4895 ( 
.A(n_3132),
.Y(n_4895)
);

CKINVDCx16_ASAP7_75t_R g4896 ( 
.A(n_1683),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_133),
.Y(n_4897)
);

CKINVDCx14_ASAP7_75t_R g4898 ( 
.A(n_1924),
.Y(n_4898)
);

BUFx3_ASAP7_75t_L g4899 ( 
.A(n_1105),
.Y(n_4899)
);

CKINVDCx5p33_ASAP7_75t_R g4900 ( 
.A(n_3304),
.Y(n_4900)
);

CKINVDCx5p33_ASAP7_75t_R g4901 ( 
.A(n_2714),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_3273),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_2152),
.Y(n_4903)
);

CKINVDCx20_ASAP7_75t_R g4904 ( 
.A(n_2512),
.Y(n_4904)
);

CKINVDCx5p33_ASAP7_75t_R g4905 ( 
.A(n_2761),
.Y(n_4905)
);

CKINVDCx5p33_ASAP7_75t_R g4906 ( 
.A(n_3033),
.Y(n_4906)
);

CKINVDCx14_ASAP7_75t_R g4907 ( 
.A(n_1762),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_1500),
.Y(n_4908)
);

HB1xp67_ASAP7_75t_L g4909 ( 
.A(n_2794),
.Y(n_4909)
);

INVx1_ASAP7_75t_SL g4910 ( 
.A(n_1100),
.Y(n_4910)
);

CKINVDCx5p33_ASAP7_75t_R g4911 ( 
.A(n_2597),
.Y(n_4911)
);

CKINVDCx5p33_ASAP7_75t_R g4912 ( 
.A(n_1510),
.Y(n_4912)
);

CKINVDCx5p33_ASAP7_75t_R g4913 ( 
.A(n_374),
.Y(n_4913)
);

CKINVDCx20_ASAP7_75t_R g4914 ( 
.A(n_274),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_2172),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_2949),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_1294),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_2930),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_724),
.Y(n_4919)
);

CKINVDCx20_ASAP7_75t_R g4920 ( 
.A(n_209),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_2709),
.Y(n_4921)
);

CKINVDCx5p33_ASAP7_75t_R g4922 ( 
.A(n_3277),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_2317),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_3172),
.Y(n_4924)
);

CKINVDCx5p33_ASAP7_75t_R g4925 ( 
.A(n_3342),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_849),
.Y(n_4926)
);

CKINVDCx5p33_ASAP7_75t_R g4927 ( 
.A(n_66),
.Y(n_4927)
);

CKINVDCx5p33_ASAP7_75t_R g4928 ( 
.A(n_173),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_3099),
.Y(n_4929)
);

CKINVDCx20_ASAP7_75t_R g4930 ( 
.A(n_2522),
.Y(n_4930)
);

CKINVDCx5p33_ASAP7_75t_R g4931 ( 
.A(n_3244),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_2994),
.Y(n_4932)
);

CKINVDCx5p33_ASAP7_75t_R g4933 ( 
.A(n_3054),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_1589),
.Y(n_4934)
);

CKINVDCx5p33_ASAP7_75t_R g4935 ( 
.A(n_176),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_2103),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_478),
.Y(n_4937)
);

CKINVDCx5p33_ASAP7_75t_R g4938 ( 
.A(n_2530),
.Y(n_4938)
);

CKINVDCx5p33_ASAP7_75t_R g4939 ( 
.A(n_2872),
.Y(n_4939)
);

CKINVDCx5p33_ASAP7_75t_R g4940 ( 
.A(n_3285),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_2446),
.Y(n_4941)
);

BUFx2_ASAP7_75t_L g4942 ( 
.A(n_934),
.Y(n_4942)
);

CKINVDCx5p33_ASAP7_75t_R g4943 ( 
.A(n_803),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_2191),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_2071),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_2541),
.Y(n_4946)
);

CKINVDCx5p33_ASAP7_75t_R g4947 ( 
.A(n_2751),
.Y(n_4947)
);

CKINVDCx5p33_ASAP7_75t_R g4948 ( 
.A(n_2725),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_3427),
.Y(n_4949)
);

CKINVDCx5p33_ASAP7_75t_R g4950 ( 
.A(n_171),
.Y(n_4950)
);

CKINVDCx5p33_ASAP7_75t_R g4951 ( 
.A(n_603),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_1762),
.Y(n_4952)
);

CKINVDCx20_ASAP7_75t_R g4953 ( 
.A(n_1703),
.Y(n_4953)
);

BUFx6f_ASAP7_75t_L g4954 ( 
.A(n_3455),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_1972),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_2141),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_665),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_268),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_159),
.Y(n_4959)
);

CKINVDCx5p33_ASAP7_75t_R g4960 ( 
.A(n_2441),
.Y(n_4960)
);

BUFx6f_ASAP7_75t_L g4961 ( 
.A(n_348),
.Y(n_4961)
);

CKINVDCx5p33_ASAP7_75t_R g4962 ( 
.A(n_3479),
.Y(n_4962)
);

CKINVDCx5p33_ASAP7_75t_R g4963 ( 
.A(n_294),
.Y(n_4963)
);

BUFx6f_ASAP7_75t_L g4964 ( 
.A(n_97),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_1750),
.Y(n_4965)
);

CKINVDCx5p33_ASAP7_75t_R g4966 ( 
.A(n_222),
.Y(n_4966)
);

CKINVDCx5p33_ASAP7_75t_R g4967 ( 
.A(n_2753),
.Y(n_4967)
);

CKINVDCx5p33_ASAP7_75t_R g4968 ( 
.A(n_2110),
.Y(n_4968)
);

CKINVDCx5p33_ASAP7_75t_R g4969 ( 
.A(n_2841),
.Y(n_4969)
);

BUFx2_ASAP7_75t_L g4970 ( 
.A(n_2888),
.Y(n_4970)
);

CKINVDCx14_ASAP7_75t_R g4971 ( 
.A(n_3291),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_3270),
.Y(n_4972)
);

CKINVDCx5p33_ASAP7_75t_R g4973 ( 
.A(n_1515),
.Y(n_4973)
);

CKINVDCx5p33_ASAP7_75t_R g4974 ( 
.A(n_1016),
.Y(n_4974)
);

CKINVDCx5p33_ASAP7_75t_R g4975 ( 
.A(n_1577),
.Y(n_4975)
);

CKINVDCx5p33_ASAP7_75t_R g4976 ( 
.A(n_3033),
.Y(n_4976)
);

CKINVDCx5p33_ASAP7_75t_R g4977 ( 
.A(n_770),
.Y(n_4977)
);

INVx2_ASAP7_75t_SL g4978 ( 
.A(n_1665),
.Y(n_4978)
);

CKINVDCx20_ASAP7_75t_R g4979 ( 
.A(n_3184),
.Y(n_4979)
);

INVx2_ASAP7_75t_L g4980 ( 
.A(n_2010),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_103),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_3283),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_999),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_181),
.Y(n_4984)
);

CKINVDCx5p33_ASAP7_75t_R g4985 ( 
.A(n_90),
.Y(n_4985)
);

CKINVDCx5p33_ASAP7_75t_R g4986 ( 
.A(n_2342),
.Y(n_4986)
);

CKINVDCx16_ASAP7_75t_R g4987 ( 
.A(n_1225),
.Y(n_4987)
);

BUFx10_ASAP7_75t_L g4988 ( 
.A(n_1200),
.Y(n_4988)
);

CKINVDCx5p33_ASAP7_75t_R g4989 ( 
.A(n_273),
.Y(n_4989)
);

BUFx2_ASAP7_75t_SL g4990 ( 
.A(n_3353),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_2854),
.Y(n_4991)
);

BUFx10_ASAP7_75t_L g4992 ( 
.A(n_2835),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_3287),
.Y(n_4993)
);

CKINVDCx5p33_ASAP7_75t_R g4994 ( 
.A(n_1296),
.Y(n_4994)
);

CKINVDCx16_ASAP7_75t_R g4995 ( 
.A(n_359),
.Y(n_4995)
);

CKINVDCx5p33_ASAP7_75t_R g4996 ( 
.A(n_853),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_3456),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_2853),
.Y(n_4998)
);

BUFx10_ASAP7_75t_L g4999 ( 
.A(n_3230),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_3527),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_2119),
.Y(n_5001)
);

CKINVDCx5p33_ASAP7_75t_R g5002 ( 
.A(n_1262),
.Y(n_5002)
);

CKINVDCx5p33_ASAP7_75t_R g5003 ( 
.A(n_1315),
.Y(n_5003)
);

CKINVDCx5p33_ASAP7_75t_R g5004 ( 
.A(n_1235),
.Y(n_5004)
);

CKINVDCx5p33_ASAP7_75t_R g5005 ( 
.A(n_985),
.Y(n_5005)
);

CKINVDCx5p33_ASAP7_75t_R g5006 ( 
.A(n_1607),
.Y(n_5006)
);

CKINVDCx5p33_ASAP7_75t_R g5007 ( 
.A(n_1203),
.Y(n_5007)
);

CKINVDCx5p33_ASAP7_75t_R g5008 ( 
.A(n_1575),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_2991),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_477),
.Y(n_5010)
);

CKINVDCx5p33_ASAP7_75t_R g5011 ( 
.A(n_1296),
.Y(n_5011)
);

CKINVDCx5p33_ASAP7_75t_R g5012 ( 
.A(n_687),
.Y(n_5012)
);

CKINVDCx20_ASAP7_75t_R g5013 ( 
.A(n_2867),
.Y(n_5013)
);

CKINVDCx5p33_ASAP7_75t_R g5014 ( 
.A(n_2485),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_132),
.Y(n_5015)
);

CKINVDCx5p33_ASAP7_75t_R g5016 ( 
.A(n_3036),
.Y(n_5016)
);

CKINVDCx5p33_ASAP7_75t_R g5017 ( 
.A(n_3274),
.Y(n_5017)
);

CKINVDCx5p33_ASAP7_75t_R g5018 ( 
.A(n_1571),
.Y(n_5018)
);

CKINVDCx5p33_ASAP7_75t_R g5019 ( 
.A(n_2906),
.Y(n_5019)
);

CKINVDCx5p33_ASAP7_75t_R g5020 ( 
.A(n_2348),
.Y(n_5020)
);

CKINVDCx5p33_ASAP7_75t_R g5021 ( 
.A(n_2659),
.Y(n_5021)
);

CKINVDCx5p33_ASAP7_75t_R g5022 ( 
.A(n_2003),
.Y(n_5022)
);

CKINVDCx5p33_ASAP7_75t_R g5023 ( 
.A(n_1907),
.Y(n_5023)
);

CKINVDCx5p33_ASAP7_75t_R g5024 ( 
.A(n_207),
.Y(n_5024)
);

CKINVDCx5p33_ASAP7_75t_R g5025 ( 
.A(n_2360),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_3204),
.Y(n_5026)
);

CKINVDCx5p33_ASAP7_75t_R g5027 ( 
.A(n_3213),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_3075),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_88),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_1244),
.Y(n_5030)
);

CKINVDCx5p33_ASAP7_75t_R g5031 ( 
.A(n_2285),
.Y(n_5031)
);

INVx2_ASAP7_75t_SL g5032 ( 
.A(n_41),
.Y(n_5032)
);

CKINVDCx5p33_ASAP7_75t_R g5033 ( 
.A(n_3081),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_3550),
.Y(n_5034)
);

INVx2_ASAP7_75t_SL g5035 ( 
.A(n_1800),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_2727),
.Y(n_5036)
);

CKINVDCx5p33_ASAP7_75t_R g5037 ( 
.A(n_834),
.Y(n_5037)
);

BUFx8_ASAP7_75t_SL g5038 ( 
.A(n_1877),
.Y(n_5038)
);

CKINVDCx5p33_ASAP7_75t_R g5039 ( 
.A(n_3236),
.Y(n_5039)
);

CKINVDCx5p33_ASAP7_75t_R g5040 ( 
.A(n_1613),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_514),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_3682),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_3682),
.Y(n_5043)
);

INVx2_ASAP7_75t_L g5044 ( 
.A(n_3682),
.Y(n_5044)
);

NOR2xp67_ASAP7_75t_L g5045 ( 
.A(n_3661),
.B(n_0),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_3682),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_3682),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_3858),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_3858),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_3858),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_3858),
.Y(n_5051)
);

CKINVDCx16_ASAP7_75t_R g5052 ( 
.A(n_3650),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_3858),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4019),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_3679),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4019),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4019),
.Y(n_5057)
);

BUFx3_ASAP7_75t_L g5058 ( 
.A(n_3698),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4019),
.Y(n_5059)
);

BUFx10_ASAP7_75t_L g5060 ( 
.A(n_3810),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4019),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4192),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4197),
.Y(n_5063)
);

BUFx2_ASAP7_75t_L g5064 ( 
.A(n_4377),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4192),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4192),
.Y(n_5066)
);

CKINVDCx5p33_ASAP7_75t_R g5067 ( 
.A(n_4472),
.Y(n_5067)
);

CKINVDCx5p33_ASAP7_75t_R g5068 ( 
.A(n_5038),
.Y(n_5068)
);

BUFx2_ASAP7_75t_L g5069 ( 
.A(n_3761),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4192),
.Y(n_5070)
);

BUFx2_ASAP7_75t_L g5071 ( 
.A(n_3908),
.Y(n_5071)
);

INVxp67_ASAP7_75t_SL g5072 ( 
.A(n_4580),
.Y(n_5072)
);

INVx2_ASAP7_75t_SL g5073 ( 
.A(n_3633),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4192),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4626),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4626),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4626),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4626),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_3635),
.Y(n_5079)
);

CKINVDCx5p33_ASAP7_75t_R g5080 ( 
.A(n_3669),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_3703),
.Y(n_5081)
);

INVx1_ASAP7_75t_SL g5082 ( 
.A(n_4028),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4626),
.Y(n_5083)
);

CKINVDCx5p33_ASAP7_75t_R g5084 ( 
.A(n_3719),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_3661),
.Y(n_5085)
);

INVx2_ASAP7_75t_SL g5086 ( 
.A(n_3633),
.Y(n_5086)
);

CKINVDCx5p33_ASAP7_75t_R g5087 ( 
.A(n_3771),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_3711),
.Y(n_5088)
);

BUFx6f_ASAP7_75t_L g5089 ( 
.A(n_3649),
.Y(n_5089)
);

INVx2_ASAP7_75t_SL g5090 ( 
.A(n_3738),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_3711),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_3649),
.Y(n_5092)
);

CKINVDCx5p33_ASAP7_75t_R g5093 ( 
.A(n_3806),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_3649),
.Y(n_5094)
);

CKINVDCx5p33_ASAP7_75t_R g5095 ( 
.A(n_3807),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_3673),
.Y(n_5096)
);

BUFx2_ASAP7_75t_L g5097 ( 
.A(n_4031),
.Y(n_5097)
);

CKINVDCx20_ASAP7_75t_R g5098 ( 
.A(n_3760),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_3673),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_3812),
.Y(n_5100)
);

CKINVDCx5p33_ASAP7_75t_R g5101 ( 
.A(n_3864),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_3673),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_3744),
.Y(n_5103)
);

INVx2_ASAP7_75t_L g5104 ( 
.A(n_3744),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_3744),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_3794),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_3794),
.Y(n_5107)
);

CKINVDCx5p33_ASAP7_75t_R g5108 ( 
.A(n_3867),
.Y(n_5108)
);

BUFx10_ASAP7_75t_L g5109 ( 
.A(n_3938),
.Y(n_5109)
);

CKINVDCx5p33_ASAP7_75t_R g5110 ( 
.A(n_3886),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_3794),
.Y(n_5111)
);

NOR2xp67_ASAP7_75t_L g5112 ( 
.A(n_4038),
.B(n_0),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_3916),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_3814),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_3814),
.Y(n_5115)
);

BUFx5_ASAP7_75t_L g5116 ( 
.A(n_3637),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_3814),
.Y(n_5117)
);

CKINVDCx16_ASAP7_75t_R g5118 ( 
.A(n_3740),
.Y(n_5118)
);

BUFx6f_ASAP7_75t_L g5119 ( 
.A(n_3815),
.Y(n_5119)
);

BUFx6f_ASAP7_75t_L g5120 ( 
.A(n_3815),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_3815),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_3852),
.Y(n_5122)
);

NOR2xp33_ASAP7_75t_L g5123 ( 
.A(n_3767),
.B(n_1),
.Y(n_5123)
);

OR2x2_ASAP7_75t_L g5124 ( 
.A(n_4109),
.B(n_1),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_3939),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_3852),
.Y(n_5126)
);

CKINVDCx5p33_ASAP7_75t_R g5127 ( 
.A(n_4012),
.Y(n_5127)
);

INVxp67_ASAP7_75t_SL g5128 ( 
.A(n_3726),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_3852),
.Y(n_5129)
);

CKINVDCx5p33_ASAP7_75t_R g5130 ( 
.A(n_4014),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_3919),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_3919),
.Y(n_5132)
);

CKINVDCx5p33_ASAP7_75t_R g5133 ( 
.A(n_4041),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_3919),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_3936),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_3936),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_4061),
.Y(n_5137)
);

CKINVDCx5p33_ASAP7_75t_R g5138 ( 
.A(n_4085),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_3936),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_3942),
.Y(n_5140)
);

CKINVDCx5p33_ASAP7_75t_R g5141 ( 
.A(n_4097),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_3942),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_3942),
.Y(n_5143)
);

CKINVDCx5p33_ASAP7_75t_R g5144 ( 
.A(n_4111),
.Y(n_5144)
);

CKINVDCx20_ASAP7_75t_R g5145 ( 
.A(n_3957),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_3962),
.Y(n_5146)
);

CKINVDCx5p33_ASAP7_75t_R g5147 ( 
.A(n_4118),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_3962),
.Y(n_5148)
);

BUFx3_ASAP7_75t_L g5149 ( 
.A(n_4718),
.Y(n_5149)
);

CKINVDCx5p33_ASAP7_75t_R g5150 ( 
.A(n_4121),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_3962),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_4152),
.Y(n_5152)
);

CKINVDCx20_ASAP7_75t_R g5153 ( 
.A(n_4170),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_3967),
.Y(n_5154)
);

CKINVDCx5p33_ASAP7_75t_R g5155 ( 
.A(n_4224),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_3967),
.Y(n_5156)
);

INVx3_ASAP7_75t_L g5157 ( 
.A(n_3658),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_3967),
.Y(n_5158)
);

BUFx3_ASAP7_75t_L g5159 ( 
.A(n_4854),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4009),
.Y(n_5160)
);

CKINVDCx5p33_ASAP7_75t_R g5161 ( 
.A(n_4234),
.Y(n_5161)
);

CKINVDCx5p33_ASAP7_75t_R g5162 ( 
.A(n_4276),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4009),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4009),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4053),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4053),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_4053),
.Y(n_5167)
);

INVxp67_ASAP7_75t_SL g5168 ( 
.A(n_4221),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4140),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4140),
.Y(n_5170)
);

NOR2xp67_ASAP7_75t_L g5171 ( 
.A(n_4167),
.B(n_2),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4140),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4153),
.Y(n_5173)
);

INVxp33_ASAP7_75t_SL g5174 ( 
.A(n_3966),
.Y(n_5174)
);

BUFx5_ASAP7_75t_L g5175 ( 
.A(n_3694),
.Y(n_5175)
);

CKINVDCx5p33_ASAP7_75t_R g5176 ( 
.A(n_4336),
.Y(n_5176)
);

INVx2_ASAP7_75t_SL g5177 ( 
.A(n_3738),
.Y(n_5177)
);

CKINVDCx5p33_ASAP7_75t_R g5178 ( 
.A(n_4343),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_4370),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4153),
.Y(n_5180)
);

CKINVDCx20_ASAP7_75t_R g5181 ( 
.A(n_4218),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_4153),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4182),
.Y(n_5183)
);

CKINVDCx20_ASAP7_75t_R g5184 ( 
.A(n_4311),
.Y(n_5184)
);

CKINVDCx5p33_ASAP7_75t_R g5185 ( 
.A(n_4385),
.Y(n_5185)
);

CKINVDCx5p33_ASAP7_75t_R g5186 ( 
.A(n_4422),
.Y(n_5186)
);

BUFx6f_ASAP7_75t_L g5187 ( 
.A(n_4182),
.Y(n_5187)
);

CKINVDCx5p33_ASAP7_75t_R g5188 ( 
.A(n_4439),
.Y(n_5188)
);

INVx1_ASAP7_75t_SL g5189 ( 
.A(n_4459),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4182),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_4442),
.Y(n_5191)
);

CKINVDCx5p33_ASAP7_75t_R g5192 ( 
.A(n_4557),
.Y(n_5192)
);

CKINVDCx5p33_ASAP7_75t_R g5193 ( 
.A(n_4756),
.Y(n_5193)
);

CKINVDCx5p33_ASAP7_75t_R g5194 ( 
.A(n_4881),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_4183),
.Y(n_5195)
);

CKINVDCx5p33_ASAP7_75t_R g5196 ( 
.A(n_4891),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4183),
.Y(n_5197)
);

CKINVDCx5p33_ASAP7_75t_R g5198 ( 
.A(n_4962),
.Y(n_5198)
);

CKINVDCx20_ASAP7_75t_R g5199 ( 
.A(n_3891),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_4997),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4183),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_4210),
.Y(n_5202)
);

CKINVDCx5p33_ASAP7_75t_R g5203 ( 
.A(n_5034),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_3952),
.Y(n_5204)
);

CKINVDCx5p33_ASAP7_75t_R g5205 ( 
.A(n_4011),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4210),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4210),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4305),
.Y(n_5208)
);

CKINVDCx5p33_ASAP7_75t_R g5209 ( 
.A(n_4228),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_4305),
.Y(n_5210)
);

CKINVDCx5p33_ASAP7_75t_R g5211 ( 
.A(n_4504),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_4898),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_4305),
.Y(n_5213)
);

CKINVDCx5p33_ASAP7_75t_R g5214 ( 
.A(n_4907),
.Y(n_5214)
);

BUFx10_ASAP7_75t_L g5215 ( 
.A(n_4101),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_4326),
.Y(n_5216)
);

CKINVDCx20_ASAP7_75t_R g5217 ( 
.A(n_4536),
.Y(n_5217)
);

CKINVDCx5p33_ASAP7_75t_R g5218 ( 
.A(n_4971),
.Y(n_5218)
);

INVx2_ASAP7_75t_SL g5219 ( 
.A(n_3795),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4326),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_4326),
.Y(n_5221)
);

INVx1_ASAP7_75t_SL g5222 ( 
.A(n_4556),
.Y(n_5222)
);

CKINVDCx16_ASAP7_75t_R g5223 ( 
.A(n_3825),
.Y(n_5223)
);

CKINVDCx5p33_ASAP7_75t_R g5224 ( 
.A(n_3888),
.Y(n_5224)
);

CKINVDCx5p33_ASAP7_75t_R g5225 ( 
.A(n_3935),
.Y(n_5225)
);

CKINVDCx5p33_ASAP7_75t_R g5226 ( 
.A(n_3950),
.Y(n_5226)
);

CKINVDCx5p33_ASAP7_75t_R g5227 ( 
.A(n_4079),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_4328),
.Y(n_5228)
);

CKINVDCx20_ASAP7_75t_R g5229 ( 
.A(n_4130),
.Y(n_5229)
);

BUFx6f_ASAP7_75t_L g5230 ( 
.A(n_4328),
.Y(n_5230)
);

CKINVDCx5p33_ASAP7_75t_R g5231 ( 
.A(n_4216),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_4235),
.Y(n_5232)
);

BUFx6f_ASAP7_75t_L g5233 ( 
.A(n_4328),
.Y(n_5233)
);

INVx2_ASAP7_75t_L g5234 ( 
.A(n_4345),
.Y(n_5234)
);

NOR2xp67_ASAP7_75t_L g5235 ( 
.A(n_4205),
.B(n_2),
.Y(n_5235)
);

CKINVDCx5p33_ASAP7_75t_R g5236 ( 
.A(n_4254),
.Y(n_5236)
);

CKINVDCx5p33_ASAP7_75t_R g5237 ( 
.A(n_4263),
.Y(n_5237)
);

CKINVDCx5p33_ASAP7_75t_R g5238 ( 
.A(n_4421),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_4345),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4345),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4358),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4358),
.Y(n_5242)
);

CKINVDCx5p33_ASAP7_75t_R g5243 ( 
.A(n_4449),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_4358),
.Y(n_5244)
);

CKINVDCx5p33_ASAP7_75t_R g5245 ( 
.A(n_4600),
.Y(n_5245)
);

BUFx2_ASAP7_75t_L g5246 ( 
.A(n_4683),
.Y(n_5246)
);

INVxp67_ASAP7_75t_SL g5247 ( 
.A(n_4154),
.Y(n_5247)
);

CKINVDCx5p33_ASAP7_75t_R g5248 ( 
.A(n_4611),
.Y(n_5248)
);

CKINVDCx5p33_ASAP7_75t_R g5249 ( 
.A(n_4710),
.Y(n_5249)
);

CKINVDCx5p33_ASAP7_75t_R g5250 ( 
.A(n_4723),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_4392),
.Y(n_5251)
);

CKINVDCx5p33_ASAP7_75t_R g5252 ( 
.A(n_4877),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_4392),
.Y(n_5253)
);

CKINVDCx5p33_ASAP7_75t_R g5254 ( 
.A(n_4896),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_4987),
.Y(n_5255)
);

CKINVDCx20_ASAP7_75t_R g5256 ( 
.A(n_4995),
.Y(n_5256)
);

INVx1_ASAP7_75t_SL g5257 ( 
.A(n_4763),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_4392),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_4401),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_4401),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_4401),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_4413),
.Y(n_5262)
);

CKINVDCx5p33_ASAP7_75t_R g5263 ( 
.A(n_5039),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_4413),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_4413),
.Y(n_5265)
);

CKINVDCx5p33_ASAP7_75t_R g5266 ( 
.A(n_3632),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_4637),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4637),
.Y(n_5268)
);

CKINVDCx14_ASAP7_75t_R g5269 ( 
.A(n_4783),
.Y(n_5269)
);

BUFx3_ASAP7_75t_L g5270 ( 
.A(n_3793),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_4637),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_4682),
.Y(n_5272)
);

CKINVDCx5p33_ASAP7_75t_R g5273 ( 
.A(n_5027),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_4682),
.Y(n_5274)
);

CKINVDCx5p33_ASAP7_75t_R g5275 ( 
.A(n_5030),
.Y(n_5275)
);

NOR2xp67_ASAP7_75t_L g5276 ( 
.A(n_4333),
.B(n_3),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_5031),
.Y(n_5277)
);

CKINVDCx5p33_ASAP7_75t_R g5278 ( 
.A(n_5033),
.Y(n_5278)
);

INVx1_ASAP7_75t_SL g5279 ( 
.A(n_4836),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4682),
.Y(n_5280)
);

INVxp67_ASAP7_75t_L g5281 ( 
.A(n_4942),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4727),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4727),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_5037),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4727),
.Y(n_5285)
);

CKINVDCx5p33_ASAP7_75t_R g5286 ( 
.A(n_5040),
.Y(n_5286)
);

BUFx5_ASAP7_75t_L g5287 ( 
.A(n_3710),
.Y(n_5287)
);

INVxp33_ASAP7_75t_L g5288 ( 
.A(n_4247),
.Y(n_5288)
);

CKINVDCx5p33_ASAP7_75t_R g5289 ( 
.A(n_3634),
.Y(n_5289)
);

NOR2xp67_ASAP7_75t_L g5290 ( 
.A(n_4616),
.B(n_4),
.Y(n_5290)
);

CKINVDCx14_ASAP7_75t_R g5291 ( 
.A(n_4970),
.Y(n_5291)
);

CKINVDCx20_ASAP7_75t_R g5292 ( 
.A(n_3659),
.Y(n_5292)
);

BUFx6f_ASAP7_75t_L g5293 ( 
.A(n_4757),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_4757),
.Y(n_5294)
);

INVx2_ASAP7_75t_L g5295 ( 
.A(n_4757),
.Y(n_5295)
);

CKINVDCx5p33_ASAP7_75t_R g5296 ( 
.A(n_5022),
.Y(n_5296)
);

CKINVDCx5p33_ASAP7_75t_R g5297 ( 
.A(n_5023),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_4781),
.Y(n_5298)
);

BUFx3_ASAP7_75t_L g5299 ( 
.A(n_3903),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_5025),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4781),
.Y(n_5301)
);

CKINVDCx5p33_ASAP7_75t_R g5302 ( 
.A(n_3636),
.Y(n_5302)
);

INVx2_ASAP7_75t_SL g5303 ( 
.A(n_3795),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4781),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4840),
.Y(n_5305)
);

CKINVDCx5p33_ASAP7_75t_R g5306 ( 
.A(n_3638),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_4840),
.Y(n_5307)
);

BUFx2_ASAP7_75t_L g5308 ( 
.A(n_3917),
.Y(n_5308)
);

CKINVDCx5p33_ASAP7_75t_R g5309 ( 
.A(n_3640),
.Y(n_5309)
);

CKINVDCx5p33_ASAP7_75t_R g5310 ( 
.A(n_3641),
.Y(n_5310)
);

CKINVDCx14_ASAP7_75t_R g5311 ( 
.A(n_3816),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_4840),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_4961),
.Y(n_5313)
);

INVxp67_ASAP7_75t_L g5314 ( 
.A(n_4490),
.Y(n_5314)
);

CKINVDCx16_ASAP7_75t_R g5315 ( 
.A(n_3816),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_4961),
.Y(n_5316)
);

CKINVDCx16_ASAP7_75t_R g5317 ( 
.A(n_3844),
.Y(n_5317)
);

CKINVDCx5p33_ASAP7_75t_R g5318 ( 
.A(n_5017),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_4961),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4964),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4964),
.Y(n_5321)
);

CKINVDCx5p33_ASAP7_75t_R g5322 ( 
.A(n_5019),
.Y(n_5322)
);

INVx2_ASAP7_75t_L g5323 ( 
.A(n_4964),
.Y(n_5323)
);

INVx1_ASAP7_75t_SL g5324 ( 
.A(n_3671),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_3940),
.Y(n_5325)
);

BUFx8_ASAP7_75t_SL g5326 ( 
.A(n_3675),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_3972),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_3991),
.Y(n_5328)
);

BUFx2_ASAP7_75t_L g5329 ( 
.A(n_4082),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4110),
.Y(n_5330)
);

CKINVDCx20_ASAP7_75t_R g5331 ( 
.A(n_3693),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4163),
.Y(n_5332)
);

INVxp67_ASAP7_75t_SL g5333 ( 
.A(n_4680),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_4169),
.Y(n_5334)
);

CKINVDCx5p33_ASAP7_75t_R g5335 ( 
.A(n_5014),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4292),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4334),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_4340),
.Y(n_5338)
);

BUFx6f_ASAP7_75t_L g5339 ( 
.A(n_4351),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_4356),
.Y(n_5340)
);

CKINVDCx5p33_ASAP7_75t_R g5341 ( 
.A(n_5024),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_4359),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4387),
.Y(n_5343)
);

CKINVDCx5p33_ASAP7_75t_R g5344 ( 
.A(n_3642),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_4436),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_4448),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4785),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_3895),
.B(n_4),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4802),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_4804),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4847),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_4852),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_4899),
.Y(n_5353)
);

CKINVDCx5p33_ASAP7_75t_R g5354 ( 
.A(n_5016),
.Y(n_5354)
);

NOR2xp67_ASAP7_75t_L g5355 ( 
.A(n_4641),
.B(n_5),
.Y(n_5355)
);

CKINVDCx5p33_ASAP7_75t_R g5356 ( 
.A(n_5020),
.Y(n_5356)
);

BUFx3_ASAP7_75t_L g5357 ( 
.A(n_3844),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5026),
.Y(n_5358)
);

INVx2_ASAP7_75t_L g5359 ( 
.A(n_3639),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_5029),
.Y(n_5360)
);

INVx2_ASAP7_75t_L g5361 ( 
.A(n_3644),
.Y(n_5361)
);

BUFx3_ASAP7_75t_L g5362 ( 
.A(n_3912),
.Y(n_5362)
);

INVx1_ASAP7_75t_SL g5363 ( 
.A(n_3801),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_3643),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_3646),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_3647),
.Y(n_5366)
);

CKINVDCx5p33_ASAP7_75t_R g5367 ( 
.A(n_5007),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5010),
.Y(n_5368)
);

CKINVDCx5p33_ASAP7_75t_R g5369 ( 
.A(n_5008),
.Y(n_5369)
);

INVx2_ASAP7_75t_SL g5370 ( 
.A(n_3912),
.Y(n_5370)
);

CKINVDCx20_ASAP7_75t_R g5371 ( 
.A(n_3716),
.Y(n_5371)
);

INVx2_ASAP7_75t_SL g5372 ( 
.A(n_3914),
.Y(n_5372)
);

CKINVDCx20_ASAP7_75t_R g5373 ( 
.A(n_3753),
.Y(n_5373)
);

BUFx10_ASAP7_75t_L g5374 ( 
.A(n_4738),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_5018),
.Y(n_5375)
);

CKINVDCx5p33_ASAP7_75t_R g5376 ( 
.A(n_5021),
.Y(n_5376)
);

BUFx2_ASAP7_75t_L g5377 ( 
.A(n_4868),
.Y(n_5377)
);

INVxp67_ASAP7_75t_L g5378 ( 
.A(n_4909),
.Y(n_5378)
);

INVx2_ASAP7_75t_L g5379 ( 
.A(n_3645),
.Y(n_5379)
);

CKINVDCx5p33_ASAP7_75t_R g5380 ( 
.A(n_3648),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5036),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_3652),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_3654),
.Y(n_5383)
);

CKINVDCx16_ASAP7_75t_R g5384 ( 
.A(n_3914),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5015),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5028),
.Y(n_5386)
);

INVx1_ASAP7_75t_SL g5387 ( 
.A(n_3818),
.Y(n_5387)
);

CKINVDCx5p33_ASAP7_75t_R g5388 ( 
.A(n_5003),
.Y(n_5388)
);

CKINVDCx5p33_ASAP7_75t_R g5389 ( 
.A(n_5004),
.Y(n_5389)
);

CKINVDCx5p33_ASAP7_75t_R g5390 ( 
.A(n_5005),
.Y(n_5390)
);

BUFx3_ASAP7_75t_L g5391 ( 
.A(n_3954),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5041),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_5006),
.Y(n_5393)
);

CKINVDCx5p33_ASAP7_75t_R g5394 ( 
.A(n_5009),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_3657),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_5012),
.Y(n_5396)
);

BUFx6f_ASAP7_75t_L g5397 ( 
.A(n_4954),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_3651),
.Y(n_5398)
);

INVxp67_ASAP7_75t_SL g5399 ( 
.A(n_3871),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_3653),
.Y(n_5400)
);

BUFx2_ASAP7_75t_L g5401 ( 
.A(n_3655),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4993),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_4991),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4998),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_3665),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_3666),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_3667),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_4996),
.Y(n_5408)
);

BUFx2_ASAP7_75t_L g5409 ( 
.A(n_3656),
.Y(n_5409)
);

CKINVDCx5p33_ASAP7_75t_R g5410 ( 
.A(n_5002),
.Y(n_5410)
);

CKINVDCx5p33_ASAP7_75t_R g5411 ( 
.A(n_5011),
.Y(n_5411)
);

CKINVDCx20_ASAP7_75t_R g5412 ( 
.A(n_3809),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_3670),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_3674),
.Y(n_5414)
);

HB1xp67_ASAP7_75t_L g5415 ( 
.A(n_3660),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_3685),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_3686),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_4985),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_4983),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_4984),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_3704),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_3708),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_4989),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_3713),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_4994),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_3714),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_3718),
.Y(n_5427)
);

CKINVDCx5p33_ASAP7_75t_R g5428 ( 
.A(n_3663),
.Y(n_5428)
);

CKINVDCx5p33_ASAP7_75t_R g5429 ( 
.A(n_3664),
.Y(n_5429)
);

BUFx2_ASAP7_75t_SL g5430 ( 
.A(n_4253),
.Y(n_5430)
);

BUFx10_ASAP7_75t_L g5431 ( 
.A(n_3668),
.Y(n_5431)
);

INVx3_ASAP7_75t_L g5432 ( 
.A(n_3954),
.Y(n_5432)
);

CKINVDCx5p33_ASAP7_75t_R g5433 ( 
.A(n_3672),
.Y(n_5433)
);

CKINVDCx5p33_ASAP7_75t_R g5434 ( 
.A(n_4981),
.Y(n_5434)
);

CKINVDCx20_ASAP7_75t_R g5435 ( 
.A(n_3826),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_4982),
.Y(n_5436)
);

HB1xp67_ASAP7_75t_L g5437 ( 
.A(n_4986),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_3722),
.Y(n_5438)
);

CKINVDCx5p33_ASAP7_75t_R g5439 ( 
.A(n_3676),
.Y(n_5439)
);

CKINVDCx20_ASAP7_75t_R g5440 ( 
.A(n_3829),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_3723),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_3727),
.Y(n_5442)
);

CKINVDCx20_ASAP7_75t_R g5443 ( 
.A(n_3854),
.Y(n_5443)
);

BUFx2_ASAP7_75t_L g5444 ( 
.A(n_3677),
.Y(n_5444)
);

CKINVDCx5p33_ASAP7_75t_R g5445 ( 
.A(n_3678),
.Y(n_5445)
);

BUFx10_ASAP7_75t_L g5446 ( 
.A(n_3681),
.Y(n_5446)
);

CKINVDCx5p33_ASAP7_75t_R g5447 ( 
.A(n_3683),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_3730),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_3735),
.Y(n_5449)
);

BUFx6f_ASAP7_75t_L g5450 ( 
.A(n_4954),
.Y(n_5450)
);

INVx1_ASAP7_75t_SL g5451 ( 
.A(n_4115),
.Y(n_5451)
);

BUFx3_ASAP7_75t_L g5452 ( 
.A(n_3987),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_3745),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_3746),
.Y(n_5454)
);

INVx1_ASAP7_75t_SL g5455 ( 
.A(n_3985),
.Y(n_5455)
);

CKINVDCx5p33_ASAP7_75t_R g5456 ( 
.A(n_3684),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_3752),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_3754),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_3759),
.Y(n_5459)
);

OR2x2_ASAP7_75t_L g5460 ( 
.A(n_3712),
.B(n_5),
.Y(n_5460)
);

INVx2_ASAP7_75t_L g5461 ( 
.A(n_3762),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_3769),
.Y(n_5462)
);

CKINVDCx20_ASAP7_75t_R g5463 ( 
.A(n_3860),
.Y(n_5463)
);

BUFx6f_ASAP7_75t_L g5464 ( 
.A(n_4954),
.Y(n_5464)
);

INVx2_ASAP7_75t_L g5465 ( 
.A(n_3770),
.Y(n_5465)
);

INVx1_ASAP7_75t_SL g5466 ( 
.A(n_3969),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_3780),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_3783),
.Y(n_5468)
);

BUFx2_ASAP7_75t_SL g5469 ( 
.A(n_4265),
.Y(n_5469)
);

CKINVDCx5p33_ASAP7_75t_R g5470 ( 
.A(n_4977),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_3788),
.Y(n_5471)
);

BUFx6f_ASAP7_75t_L g5472 ( 
.A(n_3729),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_3796),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_3798),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_3802),
.Y(n_5475)
);

CKINVDCx16_ASAP7_75t_R g5476 ( 
.A(n_4992),
.Y(n_5476)
);

BUFx3_ASAP7_75t_L g5477 ( 
.A(n_3987),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_3805),
.Y(n_5478)
);

CKINVDCx5p33_ASAP7_75t_R g5479 ( 
.A(n_5079),
.Y(n_5479)
);

CKINVDCx20_ASAP7_75t_R g5480 ( 
.A(n_5098),
.Y(n_5480)
);

CKINVDCx20_ASAP7_75t_R g5481 ( 
.A(n_5145),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5397),
.Y(n_5482)
);

CKINVDCx16_ASAP7_75t_R g5483 ( 
.A(n_5052),
.Y(n_5483)
);

CKINVDCx5p33_ASAP7_75t_R g5484 ( 
.A(n_5080),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5397),
.Y(n_5485)
);

CKINVDCx5p33_ASAP7_75t_R g5486 ( 
.A(n_5081),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5450),
.Y(n_5487)
);

CKINVDCx14_ASAP7_75t_R g5488 ( 
.A(n_5311),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_5084),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5450),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5464),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5092),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_5464),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5089),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5089),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5119),
.Y(n_5496)
);

HB1xp67_ASAP7_75t_L g5497 ( 
.A(n_5224),
.Y(n_5497)
);

INVxp67_ASAP7_75t_SL g5498 ( 
.A(n_5058),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5119),
.Y(n_5499)
);

INVxp33_ASAP7_75t_L g5500 ( 
.A(n_5415),
.Y(n_5500)
);

INVxp67_ASAP7_75t_L g5501 ( 
.A(n_5437),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5120),
.Y(n_5502)
);

CKINVDCx16_ASAP7_75t_R g5503 ( 
.A(n_5118),
.Y(n_5503)
);

HB1xp67_ASAP7_75t_L g5504 ( 
.A(n_5225),
.Y(n_5504)
);

CKINVDCx5p33_ASAP7_75t_R g5505 ( 
.A(n_5087),
.Y(n_5505)
);

INVx2_ASAP7_75t_L g5506 ( 
.A(n_5104),
.Y(n_5506)
);

HB1xp67_ASAP7_75t_L g5507 ( 
.A(n_5226),
.Y(n_5507)
);

CKINVDCx5p33_ASAP7_75t_R g5508 ( 
.A(n_5093),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5120),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5187),
.Y(n_5510)
);

CKINVDCx20_ASAP7_75t_R g5511 ( 
.A(n_5153),
.Y(n_5511)
);

INVx1_ASAP7_75t_SL g5512 ( 
.A(n_5324),
.Y(n_5512)
);

CKINVDCx5p33_ASAP7_75t_R g5513 ( 
.A(n_5095),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5187),
.Y(n_5514)
);

CKINVDCx5p33_ASAP7_75t_R g5515 ( 
.A(n_5100),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5230),
.Y(n_5516)
);

CKINVDCx20_ASAP7_75t_R g5517 ( 
.A(n_5181),
.Y(n_5517)
);

INVxp33_ASAP7_75t_SL g5518 ( 
.A(n_5055),
.Y(n_5518)
);

CKINVDCx5p33_ASAP7_75t_R g5519 ( 
.A(n_5101),
.Y(n_5519)
);

INVxp67_ASAP7_75t_SL g5520 ( 
.A(n_5149),
.Y(n_5520)
);

CKINVDCx20_ASAP7_75t_R g5521 ( 
.A(n_5184),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5230),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5233),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5233),
.Y(n_5524)
);

INVxp33_ASAP7_75t_L g5525 ( 
.A(n_5326),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5293),
.Y(n_5526)
);

INVxp67_ASAP7_75t_SL g5527 ( 
.A(n_5159),
.Y(n_5527)
);

INVxp67_ASAP7_75t_SL g5528 ( 
.A(n_5128),
.Y(n_5528)
);

HB1xp67_ASAP7_75t_L g5529 ( 
.A(n_5227),
.Y(n_5529)
);

CKINVDCx5p33_ASAP7_75t_R g5530 ( 
.A(n_5108),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5293),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_5110),
.Y(n_5532)
);

CKINVDCx20_ASAP7_75t_R g5533 ( 
.A(n_5292),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5122),
.Y(n_5534)
);

CKINVDCx5p33_ASAP7_75t_R g5535 ( 
.A(n_5113),
.Y(n_5535)
);

CKINVDCx20_ASAP7_75t_R g5536 ( 
.A(n_5331),
.Y(n_5536)
);

CKINVDCx5p33_ASAP7_75t_R g5537 ( 
.A(n_5125),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5142),
.Y(n_5538)
);

CKINVDCx5p33_ASAP7_75t_R g5539 ( 
.A(n_5127),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5148),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_5182),
.Y(n_5541)
);

INVxp33_ASAP7_75t_SL g5542 ( 
.A(n_5063),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_5228),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5234),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_5253),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5260),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5261),
.Y(n_5547)
);

CKINVDCx5p33_ASAP7_75t_R g5548 ( 
.A(n_5130),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5295),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5298),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5313),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5323),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5094),
.Y(n_5553)
);

CKINVDCx20_ASAP7_75t_R g5554 ( 
.A(n_5371),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_5096),
.Y(n_5555)
);

CKINVDCx14_ASAP7_75t_R g5556 ( 
.A(n_5269),
.Y(n_5556)
);

INVxp33_ASAP7_75t_SL g5557 ( 
.A(n_5067),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5099),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5102),
.Y(n_5559)
);

CKINVDCx5p33_ASAP7_75t_R g5560 ( 
.A(n_5133),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_5103),
.Y(n_5561)
);

CKINVDCx5p33_ASAP7_75t_R g5562 ( 
.A(n_5137),
.Y(n_5562)
);

INVx2_ASAP7_75t_SL g5563 ( 
.A(n_5431),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5105),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5106),
.Y(n_5565)
);

CKINVDCx5p33_ASAP7_75t_R g5566 ( 
.A(n_5138),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5107),
.Y(n_5567)
);

CKINVDCx5p33_ASAP7_75t_R g5568 ( 
.A(n_5141),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_5144),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_5111),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5114),
.Y(n_5571)
);

INVx1_ASAP7_75t_SL g5572 ( 
.A(n_5363),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5115),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5117),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5121),
.Y(n_5575)
);

CKINVDCx5p33_ASAP7_75t_R g5576 ( 
.A(n_5147),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5126),
.Y(n_5577)
);

INVxp33_ASAP7_75t_SL g5578 ( 
.A(n_5068),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_5150),
.Y(n_5579)
);

CKINVDCx5p33_ASAP7_75t_R g5580 ( 
.A(n_5152),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5129),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5131),
.Y(n_5582)
);

CKINVDCx5p33_ASAP7_75t_R g5583 ( 
.A(n_5155),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_5132),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5134),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_5135),
.Y(n_5586)
);

INVxp67_ASAP7_75t_L g5587 ( 
.A(n_5401),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5136),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_5139),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5140),
.Y(n_5590)
);

CKINVDCx20_ASAP7_75t_R g5591 ( 
.A(n_5373),
.Y(n_5591)
);

INVxp67_ASAP7_75t_L g5592 ( 
.A(n_5409),
.Y(n_5592)
);

BUFx3_ASAP7_75t_L g5593 ( 
.A(n_5270),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_5143),
.Y(n_5594)
);

CKINVDCx16_ASAP7_75t_R g5595 ( 
.A(n_5223),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5146),
.Y(n_5596)
);

INVxp67_ASAP7_75t_L g5597 ( 
.A(n_5444),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5151),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5154),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5156),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5158),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_5161),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5160),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5163),
.Y(n_5604)
);

CKINVDCx20_ASAP7_75t_R g5605 ( 
.A(n_5412),
.Y(n_5605)
);

INVxp67_ASAP7_75t_SL g5606 ( 
.A(n_5157),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5164),
.Y(n_5607)
);

CKINVDCx20_ASAP7_75t_R g5608 ( 
.A(n_5435),
.Y(n_5608)
);

BUFx6f_ASAP7_75t_L g5609 ( 
.A(n_5339),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_5165),
.Y(n_5610)
);

BUFx3_ASAP7_75t_L g5611 ( 
.A(n_5299),
.Y(n_5611)
);

CKINVDCx5p33_ASAP7_75t_R g5612 ( 
.A(n_5162),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5166),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5167),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5169),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5170),
.Y(n_5616)
);

CKINVDCx5p33_ASAP7_75t_R g5617 ( 
.A(n_5176),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5172),
.Y(n_5618)
);

INVxp67_ASAP7_75t_L g5619 ( 
.A(n_5308),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5173),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5180),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5183),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5190),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5195),
.Y(n_5624)
);

CKINVDCx20_ASAP7_75t_R g5625 ( 
.A(n_5440),
.Y(n_5625)
);

CKINVDCx20_ASAP7_75t_R g5626 ( 
.A(n_5443),
.Y(n_5626)
);

CKINVDCx5p33_ASAP7_75t_R g5627 ( 
.A(n_5178),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5197),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5201),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5202),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5206),
.Y(n_5631)
);

INVxp33_ASAP7_75t_SL g5632 ( 
.A(n_5231),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5207),
.Y(n_5633)
);

INVxp67_ASAP7_75t_L g5634 ( 
.A(n_5329),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5208),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5210),
.Y(n_5636)
);

INVxp67_ASAP7_75t_SL g5637 ( 
.A(n_5339),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_5179),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5213),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5216),
.Y(n_5640)
);

CKINVDCx20_ASAP7_75t_R g5641 ( 
.A(n_5463),
.Y(n_5641)
);

INVxp67_ASAP7_75t_SL g5642 ( 
.A(n_5432),
.Y(n_5642)
);

INVxp67_ASAP7_75t_L g5643 ( 
.A(n_5357),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5220),
.Y(n_5644)
);

INVxp67_ASAP7_75t_SL g5645 ( 
.A(n_5123),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5221),
.Y(n_5646)
);

CKINVDCx20_ASAP7_75t_R g5647 ( 
.A(n_5199),
.Y(n_5647)
);

CKINVDCx20_ASAP7_75t_R g5648 ( 
.A(n_5217),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_5239),
.Y(n_5649)
);

HB1xp67_ASAP7_75t_L g5650 ( 
.A(n_5232),
.Y(n_5650)
);

CKINVDCx20_ASAP7_75t_R g5651 ( 
.A(n_5229),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5240),
.Y(n_5652)
);

CKINVDCx5p33_ASAP7_75t_R g5653 ( 
.A(n_5185),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5241),
.Y(n_5654)
);

HB1xp67_ASAP7_75t_L g5655 ( 
.A(n_5236),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5242),
.Y(n_5656)
);

CKINVDCx20_ASAP7_75t_R g5657 ( 
.A(n_5256),
.Y(n_5657)
);

INVxp33_ASAP7_75t_SL g5658 ( 
.A(n_5237),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5244),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5251),
.Y(n_5660)
);

CKINVDCx20_ASAP7_75t_R g5661 ( 
.A(n_5186),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5258),
.Y(n_5662)
);

CKINVDCx20_ASAP7_75t_R g5663 ( 
.A(n_5188),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5259),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5262),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5264),
.Y(n_5666)
);

CKINVDCx5p33_ASAP7_75t_R g5667 ( 
.A(n_5191),
.Y(n_5667)
);

HB1xp67_ASAP7_75t_L g5668 ( 
.A(n_5238),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5265),
.Y(n_5669)
);

HB1xp67_ASAP7_75t_L g5670 ( 
.A(n_5243),
.Y(n_5670)
);

CKINVDCx5p33_ASAP7_75t_R g5671 ( 
.A(n_5192),
.Y(n_5671)
);

INVxp67_ASAP7_75t_SL g5672 ( 
.A(n_5399),
.Y(n_5672)
);

CKINVDCx5p33_ASAP7_75t_R g5673 ( 
.A(n_5193),
.Y(n_5673)
);

CKINVDCx5p33_ASAP7_75t_R g5674 ( 
.A(n_5194),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5267),
.Y(n_5675)
);

BUFx6f_ASAP7_75t_L g5676 ( 
.A(n_5472),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5268),
.Y(n_5677)
);

HB1xp67_ASAP7_75t_L g5678 ( 
.A(n_5245),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5271),
.Y(n_5679)
);

INVxp33_ASAP7_75t_SL g5680 ( 
.A(n_5248),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5272),
.Y(n_5681)
);

INVx1_ASAP7_75t_L g5682 ( 
.A(n_5274),
.Y(n_5682)
);

INVxp67_ASAP7_75t_L g5683 ( 
.A(n_5362),
.Y(n_5683)
);

BUFx6f_ASAP7_75t_L g5684 ( 
.A(n_5472),
.Y(n_5684)
);

CKINVDCx5p33_ASAP7_75t_R g5685 ( 
.A(n_5196),
.Y(n_5685)
);

INVxp33_ASAP7_75t_L g5686 ( 
.A(n_5288),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5280),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5282),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_5283),
.Y(n_5689)
);

CKINVDCx5p33_ASAP7_75t_R g5690 ( 
.A(n_5198),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_5285),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5294),
.Y(n_5692)
);

INVxp67_ASAP7_75t_SL g5693 ( 
.A(n_5338),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5301),
.Y(n_5694)
);

CKINVDCx20_ASAP7_75t_R g5695 ( 
.A(n_5200),
.Y(n_5695)
);

HB1xp67_ASAP7_75t_L g5696 ( 
.A(n_5249),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_5304),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5305),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_5203),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5307),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_5312),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5316),
.Y(n_5702)
);

BUFx6f_ASAP7_75t_L g5703 ( 
.A(n_5319),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5320),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5321),
.Y(n_5705)
);

INVxp67_ASAP7_75t_L g5706 ( 
.A(n_5391),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5042),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5043),
.Y(n_5708)
);

CKINVDCx20_ASAP7_75t_R g5709 ( 
.A(n_5250),
.Y(n_5709)
);

BUFx3_ASAP7_75t_L g5710 ( 
.A(n_5325),
.Y(n_5710)
);

CKINVDCx5p33_ASAP7_75t_R g5711 ( 
.A(n_5263),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5044),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5046),
.Y(n_5713)
);

INVx2_ASAP7_75t_L g5714 ( 
.A(n_5047),
.Y(n_5714)
);

CKINVDCx5p33_ASAP7_75t_R g5715 ( 
.A(n_5266),
.Y(n_5715)
);

CKINVDCx16_ASAP7_75t_R g5716 ( 
.A(n_5315),
.Y(n_5716)
);

INVxp33_ASAP7_75t_L g5717 ( 
.A(n_5069),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5048),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5049),
.Y(n_5719)
);

INVx2_ASAP7_75t_L g5720 ( 
.A(n_5050),
.Y(n_5720)
);

CKINVDCx5p33_ASAP7_75t_R g5721 ( 
.A(n_5273),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5051),
.Y(n_5722)
);

INVxp67_ASAP7_75t_SL g5723 ( 
.A(n_5168),
.Y(n_5723)
);

BUFx2_ASAP7_75t_L g5724 ( 
.A(n_5252),
.Y(n_5724)
);

INVx1_ASAP7_75t_SL g5725 ( 
.A(n_5387),
.Y(n_5725)
);

INVxp67_ASAP7_75t_SL g5726 ( 
.A(n_5452),
.Y(n_5726)
);

CKINVDCx5p33_ASAP7_75t_R g5727 ( 
.A(n_5275),
.Y(n_5727)
);

INVxp67_ASAP7_75t_SL g5728 ( 
.A(n_5477),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5053),
.Y(n_5729)
);

INVxp67_ASAP7_75t_SL g5730 ( 
.A(n_5327),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5054),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5056),
.Y(n_5732)
);

INVx2_ASAP7_75t_L g5733 ( 
.A(n_5057),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5059),
.Y(n_5734)
);

INVxp67_ASAP7_75t_SL g5735 ( 
.A(n_5328),
.Y(n_5735)
);

INVxp67_ASAP7_75t_L g5736 ( 
.A(n_5073),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5061),
.Y(n_5737)
);

CKINVDCx20_ASAP7_75t_R g5738 ( 
.A(n_5254),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5062),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5065),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5066),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_5070),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5074),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5075),
.Y(n_5744)
);

CKINVDCx5p33_ASAP7_75t_R g5745 ( 
.A(n_5277),
.Y(n_5745)
);

INVxp67_ASAP7_75t_SL g5746 ( 
.A(n_5330),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5076),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5077),
.Y(n_5748)
);

HB1xp67_ASAP7_75t_L g5749 ( 
.A(n_5255),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5078),
.Y(n_5750)
);

CKINVDCx14_ASAP7_75t_R g5751 ( 
.A(n_5291),
.Y(n_5751)
);

CKINVDCx5p33_ASAP7_75t_R g5752 ( 
.A(n_5278),
.Y(n_5752)
);

CKINVDCx20_ASAP7_75t_R g5753 ( 
.A(n_5451),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5083),
.Y(n_5754)
);

BUFx6f_ASAP7_75t_L g5755 ( 
.A(n_5359),
.Y(n_5755)
);

HB1xp67_ASAP7_75t_L g5756 ( 
.A(n_5284),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5085),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_5088),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5091),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5358),
.Y(n_5760)
);

CKINVDCx20_ASAP7_75t_R g5761 ( 
.A(n_5455),
.Y(n_5761)
);

INVxp33_ASAP7_75t_L g5762 ( 
.A(n_5071),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5360),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5368),
.Y(n_5764)
);

CKINVDCx5p33_ASAP7_75t_R g5765 ( 
.A(n_5286),
.Y(n_5765)
);

HB1xp67_ASAP7_75t_L g5766 ( 
.A(n_5289),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5381),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5383),
.Y(n_5768)
);

CKINVDCx20_ASAP7_75t_R g5769 ( 
.A(n_5466),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5385),
.Y(n_5770)
);

BUFx6f_ASAP7_75t_L g5771 ( 
.A(n_5361),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5386),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5392),
.Y(n_5773)
);

CKINVDCx20_ASAP7_75t_R g5774 ( 
.A(n_5296),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5395),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5402),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5404),
.Y(n_5777)
);

CKINVDCx20_ASAP7_75t_R g5778 ( 
.A(n_5297),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5405),
.Y(n_5779)
);

BUFx10_ASAP7_75t_L g5780 ( 
.A(n_5204),
.Y(n_5780)
);

CKINVDCx5p33_ASAP7_75t_R g5781 ( 
.A(n_5300),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5406),
.Y(n_5782)
);

BUFx2_ASAP7_75t_L g5783 ( 
.A(n_5302),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5413),
.Y(n_5784)
);

CKINVDCx5p33_ASAP7_75t_R g5785 ( 
.A(n_5306),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5414),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5416),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5417),
.Y(n_5788)
);

CKINVDCx5p33_ASAP7_75t_R g5789 ( 
.A(n_5309),
.Y(n_5789)
);

CKINVDCx16_ASAP7_75t_R g5790 ( 
.A(n_5317),
.Y(n_5790)
);

INVxp67_ASAP7_75t_SL g5791 ( 
.A(n_5332),
.Y(n_5791)
);

INVxp67_ASAP7_75t_L g5792 ( 
.A(n_5086),
.Y(n_5792)
);

CKINVDCx20_ASAP7_75t_R g5793 ( 
.A(n_5310),
.Y(n_5793)
);

CKINVDCx20_ASAP7_75t_R g5794 ( 
.A(n_5318),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5419),
.Y(n_5795)
);

CKINVDCx16_ASAP7_75t_R g5796 ( 
.A(n_5384),
.Y(n_5796)
);

INVx1_ASAP7_75t_L g5797 ( 
.A(n_5420),
.Y(n_5797)
);

BUFx6f_ASAP7_75t_L g5798 ( 
.A(n_5379),
.Y(n_5798)
);

CKINVDCx5p33_ASAP7_75t_R g5799 ( 
.A(n_5322),
.Y(n_5799)
);

BUFx5_ASAP7_75t_L g5800 ( 
.A(n_5421),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_5422),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5424),
.Y(n_5802)
);

INVxp33_ASAP7_75t_L g5803 ( 
.A(n_5097),
.Y(n_5803)
);

INVxp33_ASAP7_75t_SL g5804 ( 
.A(n_5205),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5426),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_5335),
.Y(n_5806)
);

INVxp33_ASAP7_75t_SL g5807 ( 
.A(n_5209),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5436),
.Y(n_5808)
);

CKINVDCx5p33_ASAP7_75t_R g5809 ( 
.A(n_5341),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5438),
.Y(n_5810)
);

CKINVDCx5p33_ASAP7_75t_R g5811 ( 
.A(n_5344),
.Y(n_5811)
);

BUFx6f_ASAP7_75t_L g5812 ( 
.A(n_5382),
.Y(n_5812)
);

CKINVDCx16_ASAP7_75t_R g5813 ( 
.A(n_5476),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5441),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5442),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5448),
.Y(n_5816)
);

CKINVDCx20_ASAP7_75t_R g5817 ( 
.A(n_5354),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5449),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_5453),
.Y(n_5819)
);

CKINVDCx5p33_ASAP7_75t_R g5820 ( 
.A(n_5356),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5454),
.Y(n_5821)
);

INVxp67_ASAP7_75t_SL g5822 ( 
.A(n_5334),
.Y(n_5822)
);

INVxp67_ASAP7_75t_L g5823 ( 
.A(n_5090),
.Y(n_5823)
);

INVxp67_ASAP7_75t_SL g5824 ( 
.A(n_5336),
.Y(n_5824)
);

CKINVDCx16_ASAP7_75t_R g5825 ( 
.A(n_5064),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_5457),
.Y(n_5826)
);

CKINVDCx5p33_ASAP7_75t_R g5827 ( 
.A(n_5364),
.Y(n_5827)
);

CKINVDCx16_ASAP7_75t_R g5828 ( 
.A(n_5446),
.Y(n_5828)
);

CKINVDCx5p33_ASAP7_75t_R g5829 ( 
.A(n_5365),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5458),
.Y(n_5830)
);

INVx1_ASAP7_75t_SL g5831 ( 
.A(n_5211),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5459),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5462),
.Y(n_5833)
);

CKINVDCx5p33_ASAP7_75t_R g5834 ( 
.A(n_5366),
.Y(n_5834)
);

INVxp67_ASAP7_75t_L g5835 ( 
.A(n_5177),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5467),
.Y(n_5836)
);

INVxp33_ASAP7_75t_SL g5837 ( 
.A(n_5212),
.Y(n_5837)
);

CKINVDCx20_ASAP7_75t_R g5838 ( 
.A(n_5367),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5468),
.Y(n_5839)
);

INVxp67_ASAP7_75t_SL g5840 ( 
.A(n_5337),
.Y(n_5840)
);

CKINVDCx20_ASAP7_75t_R g5841 ( 
.A(n_5369),
.Y(n_5841)
);

BUFx3_ASAP7_75t_L g5842 ( 
.A(n_5340),
.Y(n_5842)
);

BUFx3_ASAP7_75t_L g5843 ( 
.A(n_5342),
.Y(n_5843)
);

CKINVDCx5p33_ASAP7_75t_R g5844 ( 
.A(n_5375),
.Y(n_5844)
);

INVxp33_ASAP7_75t_SL g5845 ( 
.A(n_5214),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5407),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5471),
.Y(n_5847)
);

CKINVDCx16_ASAP7_75t_R g5848 ( 
.A(n_5082),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5473),
.Y(n_5849)
);

HB1xp67_ASAP7_75t_L g5850 ( 
.A(n_5376),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5474),
.Y(n_5851)
);

INVxp67_ASAP7_75t_SL g5852 ( 
.A(n_5343),
.Y(n_5852)
);

CKINVDCx5p33_ASAP7_75t_R g5853 ( 
.A(n_5380),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5475),
.Y(n_5854)
);

INVx2_ASAP7_75t_L g5855 ( 
.A(n_5427),
.Y(n_5855)
);

BUFx2_ASAP7_75t_L g5856 ( 
.A(n_5388),
.Y(n_5856)
);

HB1xp67_ASAP7_75t_L g5857 ( 
.A(n_5389),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5478),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5461),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5465),
.Y(n_5860)
);

CKINVDCx20_ASAP7_75t_R g5861 ( 
.A(n_5390),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_5393),
.Y(n_5862)
);

CKINVDCx5p33_ASAP7_75t_R g5863 ( 
.A(n_5394),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5345),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5346),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5347),
.Y(n_5866)
);

CKINVDCx5p33_ASAP7_75t_R g5867 ( 
.A(n_5396),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5349),
.Y(n_5868)
);

INVxp67_ASAP7_75t_L g5869 ( 
.A(n_5219),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5350),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5351),
.Y(n_5871)
);

CKINVDCx5p33_ASAP7_75t_R g5872 ( 
.A(n_5398),
.Y(n_5872)
);

INVxp67_ASAP7_75t_SL g5873 ( 
.A(n_5352),
.Y(n_5873)
);

CKINVDCx5p33_ASAP7_75t_R g5874 ( 
.A(n_5400),
.Y(n_5874)
);

CKINVDCx20_ASAP7_75t_R g5875 ( 
.A(n_5403),
.Y(n_5875)
);

INVxp67_ASAP7_75t_SL g5876 ( 
.A(n_5353),
.Y(n_5876)
);

INVxp67_ASAP7_75t_SL g5877 ( 
.A(n_5348),
.Y(n_5877)
);

INVxp67_ASAP7_75t_SL g5878 ( 
.A(n_5045),
.Y(n_5878)
);

CKINVDCx20_ASAP7_75t_R g5879 ( 
.A(n_5408),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5430),
.Y(n_5880)
);

CKINVDCx20_ASAP7_75t_R g5881 ( 
.A(n_5410),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5469),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5116),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5116),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5116),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5116),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5175),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5175),
.Y(n_5888)
);

INVxp67_ASAP7_75t_SL g5889 ( 
.A(n_5314),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_5411),
.Y(n_5890)
);

INVx3_ASAP7_75t_L g5891 ( 
.A(n_5460),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5175),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5175),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5287),
.Y(n_5894)
);

INVxp67_ASAP7_75t_L g5895 ( 
.A(n_5303),
.Y(n_5895)
);

BUFx3_ASAP7_75t_L g5896 ( 
.A(n_5418),
.Y(n_5896)
);

BUFx3_ASAP7_75t_L g5897 ( 
.A(n_5423),
.Y(n_5897)
);

INVxp67_ASAP7_75t_SL g5898 ( 
.A(n_5378),
.Y(n_5898)
);

CKINVDCx20_ASAP7_75t_R g5899 ( 
.A(n_5425),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5287),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5287),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5287),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5247),
.Y(n_5903)
);

CKINVDCx5p33_ASAP7_75t_R g5904 ( 
.A(n_5428),
.Y(n_5904)
);

CKINVDCx20_ASAP7_75t_R g5905 ( 
.A(n_5429),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5333),
.Y(n_5906)
);

INVxp67_ASAP7_75t_SL g5907 ( 
.A(n_5072),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5470),
.Y(n_5908)
);

CKINVDCx5p33_ASAP7_75t_R g5909 ( 
.A(n_5433),
.Y(n_5909)
);

INVxp67_ASAP7_75t_L g5910 ( 
.A(n_5370),
.Y(n_5910)
);

INVxp67_ASAP7_75t_SL g5911 ( 
.A(n_5281),
.Y(n_5911)
);

INVxp67_ASAP7_75t_SL g5912 ( 
.A(n_5124),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5434),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5456),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5439),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5447),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5445),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5112),
.Y(n_5918)
);

INVxp67_ASAP7_75t_SL g5919 ( 
.A(n_5171),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5235),
.Y(n_5920)
);

INVxp33_ASAP7_75t_SL g5921 ( 
.A(n_5218),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_5189),
.Y(n_5922)
);

CKINVDCx5p33_ASAP7_75t_R g5923 ( 
.A(n_5222),
.Y(n_5923)
);

CKINVDCx16_ASAP7_75t_R g5924 ( 
.A(n_5257),
.Y(n_5924)
);

CKINVDCx5p33_ASAP7_75t_R g5925 ( 
.A(n_5279),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5276),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5290),
.Y(n_5927)
);

INVx1_ASAP7_75t_L g5928 ( 
.A(n_5355),
.Y(n_5928)
);

HB1xp67_ASAP7_75t_L g5929 ( 
.A(n_5372),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5377),
.Y(n_5930)
);

HB1xp67_ASAP7_75t_L g5931 ( 
.A(n_5246),
.Y(n_5931)
);

CKINVDCx5p33_ASAP7_75t_R g5932 ( 
.A(n_5174),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5060),
.Y(n_5933)
);

CKINVDCx5p33_ASAP7_75t_R g5934 ( 
.A(n_5109),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5215),
.Y(n_5935)
);

INVxp67_ASAP7_75t_SL g5936 ( 
.A(n_5374),
.Y(n_5936)
);

CKINVDCx5p33_ASAP7_75t_R g5937 ( 
.A(n_5079),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5397),
.Y(n_5938)
);

CKINVDCx20_ASAP7_75t_R g5939 ( 
.A(n_5098),
.Y(n_5939)
);

CKINVDCx5p33_ASAP7_75t_R g5940 ( 
.A(n_5079),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5397),
.Y(n_5941)
);

CKINVDCx5p33_ASAP7_75t_R g5942 ( 
.A(n_5079),
.Y(n_5942)
);

INVxp33_ASAP7_75t_L g5943 ( 
.A(n_5415),
.Y(n_5943)
);

CKINVDCx16_ASAP7_75t_R g5944 ( 
.A(n_5052),
.Y(n_5944)
);

CKINVDCx20_ASAP7_75t_R g5945 ( 
.A(n_5098),
.Y(n_5945)
);

INVx1_ASAP7_75t_SL g5946 ( 
.A(n_5324),
.Y(n_5946)
);

BUFx2_ASAP7_75t_L g5947 ( 
.A(n_5229),
.Y(n_5947)
);

INVxp67_ASAP7_75t_L g5948 ( 
.A(n_5415),
.Y(n_5948)
);

CKINVDCx16_ASAP7_75t_R g5949 ( 
.A(n_5052),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5397),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5397),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5397),
.Y(n_5952)
);

INVxp67_ASAP7_75t_L g5953 ( 
.A(n_5415),
.Y(n_5953)
);

CKINVDCx5p33_ASAP7_75t_R g5954 ( 
.A(n_5079),
.Y(n_5954)
);

BUFx3_ASAP7_75t_L g5955 ( 
.A(n_5058),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5397),
.Y(n_5956)
);

CKINVDCx5p33_ASAP7_75t_R g5957 ( 
.A(n_5079),
.Y(n_5957)
);

INVxp67_ASAP7_75t_SL g5958 ( 
.A(n_5058),
.Y(n_5958)
);

CKINVDCx5p33_ASAP7_75t_R g5959 ( 
.A(n_5079),
.Y(n_5959)
);

BUFx2_ASAP7_75t_L g5960 ( 
.A(n_5229),
.Y(n_5960)
);

HB1xp67_ASAP7_75t_L g5961 ( 
.A(n_5224),
.Y(n_5961)
);

CKINVDCx20_ASAP7_75t_R g5962 ( 
.A(n_5098),
.Y(n_5962)
);

CKINVDCx20_ASAP7_75t_R g5963 ( 
.A(n_5098),
.Y(n_5963)
);

BUFx3_ASAP7_75t_L g5964 ( 
.A(n_5058),
.Y(n_5964)
);

CKINVDCx5p33_ASAP7_75t_R g5965 ( 
.A(n_5079),
.Y(n_5965)
);

INVxp67_ASAP7_75t_SL g5966 ( 
.A(n_5058),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5397),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5397),
.Y(n_5968)
);

BUFx2_ASAP7_75t_L g5969 ( 
.A(n_5229),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5397),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5397),
.Y(n_5971)
);

INVxp67_ASAP7_75t_SL g5972 ( 
.A(n_5058),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5397),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5397),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_5079),
.Y(n_5975)
);

INVxp33_ASAP7_75t_SL g5976 ( 
.A(n_5055),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5397),
.Y(n_5977)
);

CKINVDCx5p33_ASAP7_75t_R g5978 ( 
.A(n_5079),
.Y(n_5978)
);

CKINVDCx20_ASAP7_75t_R g5979 ( 
.A(n_5098),
.Y(n_5979)
);

INVx2_ASAP7_75t_L g5980 ( 
.A(n_5092),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5397),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5397),
.Y(n_5982)
);

CKINVDCx16_ASAP7_75t_R g5983 ( 
.A(n_5052),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5397),
.Y(n_5984)
);

INVxp67_ASAP7_75t_SL g5985 ( 
.A(n_5058),
.Y(n_5985)
);

INVxp67_ASAP7_75t_L g5986 ( 
.A(n_5415),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5397),
.Y(n_5987)
);

INVx2_ASAP7_75t_L g5988 ( 
.A(n_5492),
.Y(n_5988)
);

AND2x4_ASAP7_75t_L g5989 ( 
.A(n_5955),
.B(n_5964),
.Y(n_5989)
);

NOR2xp33_ASAP7_75t_L g5990 ( 
.A(n_5528),
.B(n_4066),
.Y(n_5990)
);

AND2x4_ASAP7_75t_L g5991 ( 
.A(n_5498),
.B(n_3662),
.Y(n_5991)
);

OAI22xp5_ASAP7_75t_L g5992 ( 
.A1(n_5645),
.A2(n_4751),
.B1(n_4851),
.B2(n_4817),
.Y(n_5992)
);

BUFx6f_ASAP7_75t_L g5993 ( 
.A(n_5609),
.Y(n_5993)
);

BUFx6f_ASAP7_75t_L g5994 ( 
.A(n_5609),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5760),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5763),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5506),
.Y(n_5997)
);

BUFx6f_ASAP7_75t_L g5998 ( 
.A(n_5609),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5541),
.Y(n_5999)
);

INVx5_ASAP7_75t_L g6000 ( 
.A(n_5483),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5764),
.Y(n_6001)
);

INVx2_ASAP7_75t_L g6002 ( 
.A(n_5980),
.Y(n_6002)
);

AND2x4_ASAP7_75t_L g6003 ( 
.A(n_5520),
.B(n_4597),
.Y(n_6003)
);

INVx3_ASAP7_75t_L g6004 ( 
.A(n_5676),
.Y(n_6004)
);

BUFx6f_ASAP7_75t_L g6005 ( 
.A(n_5676),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5767),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5768),
.Y(n_6007)
);

BUFx6f_ASAP7_75t_L g6008 ( 
.A(n_5676),
.Y(n_6008)
);

INVx2_ASAP7_75t_L g6009 ( 
.A(n_5712),
.Y(n_6009)
);

INVx2_ASAP7_75t_L g6010 ( 
.A(n_5714),
.Y(n_6010)
);

INVx2_ASAP7_75t_L g6011 ( 
.A(n_5720),
.Y(n_6011)
);

CKINVDCx14_ASAP7_75t_R g6012 ( 
.A(n_5488),
.Y(n_6012)
);

BUFx8_ASAP7_75t_L g6013 ( 
.A(n_5947),
.Y(n_6013)
);

BUFx6f_ASAP7_75t_L g6014 ( 
.A(n_5684),
.Y(n_6014)
);

INVx2_ASAP7_75t_L g6015 ( 
.A(n_5755),
.Y(n_6015)
);

AND2x4_ASAP7_75t_L g6016 ( 
.A(n_5527),
.B(n_4801),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5770),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5772),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5755),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5773),
.Y(n_6020)
);

BUFx8_ASAP7_75t_L g6021 ( 
.A(n_5960),
.Y(n_6021)
);

AND2x4_ASAP7_75t_L g6022 ( 
.A(n_5958),
.B(n_3724),
.Y(n_6022)
);

OA21x2_ASAP7_75t_L g6023 ( 
.A1(n_5883),
.A2(n_4591),
.B(n_4307),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5775),
.Y(n_6024)
);

OAI21x1_ASAP7_75t_L g6025 ( 
.A1(n_5884),
.A2(n_3910),
.B(n_3881),
.Y(n_6025)
);

BUFx6f_ASAP7_75t_L g6026 ( 
.A(n_5684),
.Y(n_6026)
);

CKINVDCx6p67_ASAP7_75t_R g6027 ( 
.A(n_5848),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5966),
.B(n_3763),
.Y(n_6028)
);

BUFx6f_ASAP7_75t_L g6029 ( 
.A(n_5684),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5755),
.Y(n_6030)
);

BUFx6f_ASAP7_75t_L g6031 ( 
.A(n_5771),
.Y(n_6031)
);

OAI22xp5_ASAP7_75t_SL g6032 ( 
.A1(n_5924),
.A2(n_3915),
.B1(n_3949),
.B2(n_3883),
.Y(n_6032)
);

BUFx2_ASAP7_75t_L g6033 ( 
.A(n_5922),
.Y(n_6033)
);

INVx2_ASAP7_75t_L g6034 ( 
.A(n_5771),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5776),
.Y(n_6035)
);

OAI22xp5_ASAP7_75t_L g6036 ( 
.A1(n_5912),
.A2(n_4887),
.B1(n_3689),
.B2(n_3690),
.Y(n_6036)
);

OAI22x1_ASAP7_75t_L g6037 ( 
.A1(n_5923),
.A2(n_4843),
.B1(n_3715),
.B2(n_3728),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5771),
.Y(n_6038)
);

INVx6_ASAP7_75t_L g6039 ( 
.A(n_5593),
.Y(n_6039)
);

INVx4_ASAP7_75t_L g6040 ( 
.A(n_5479),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5777),
.Y(n_6041)
);

NAND2xp5_ASAP7_75t_L g6042 ( 
.A(n_5877),
.B(n_3687),
.Y(n_6042)
);

BUFx6f_ASAP7_75t_L g6043 ( 
.A(n_5798),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5779),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5782),
.Y(n_6045)
);

INVx2_ASAP7_75t_L g6046 ( 
.A(n_5798),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5784),
.Y(n_6047)
);

BUFx6f_ASAP7_75t_L g6048 ( 
.A(n_5798),
.Y(n_6048)
);

OAI22x1_ASAP7_75t_SL g6049 ( 
.A1(n_5925),
.A2(n_3994),
.B1(n_3997),
.B2(n_3978),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5786),
.Y(n_6050)
);

OA21x2_ASAP7_75t_L g6051 ( 
.A1(n_5885),
.A2(n_3941),
.B(n_3933),
.Y(n_6051)
);

NAND2xp5_ASAP7_75t_L g6052 ( 
.A(n_5878),
.B(n_5880),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_5812),
.Y(n_6053)
);

BUFx2_ASAP7_75t_L g6054 ( 
.A(n_5753),
.Y(n_6054)
);

INVx6_ASAP7_75t_L g6055 ( 
.A(n_5611),
.Y(n_6055)
);

HB1xp67_ASAP7_75t_L g6056 ( 
.A(n_5512),
.Y(n_6056)
);

NAND2x1p5_ASAP7_75t_L g6057 ( 
.A(n_5896),
.B(n_4491),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5787),
.Y(n_6058)
);

OA21x2_ASAP7_75t_L g6059 ( 
.A1(n_5886),
.A2(n_4185),
.B(n_4133),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5812),
.Y(n_6060)
);

INVx5_ASAP7_75t_L g6061 ( 
.A(n_5503),
.Y(n_6061)
);

INVx5_ASAP7_75t_L g6062 ( 
.A(n_5595),
.Y(n_6062)
);

HB1xp67_ASAP7_75t_L g6063 ( 
.A(n_5572),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_5484),
.Y(n_6064)
);

INVx5_ASAP7_75t_L g6065 ( 
.A(n_5944),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_5788),
.Y(n_6066)
);

AOI22xp5_ASAP7_75t_L g6067 ( 
.A1(n_5501),
.A2(n_4620),
.B1(n_3733),
.B2(n_3737),
.Y(n_6067)
);

INVxp67_ASAP7_75t_L g6068 ( 
.A(n_5725),
.Y(n_6068)
);

NOR2xp33_ASAP7_75t_SL g6069 ( 
.A(n_5828),
.B(n_4026),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5795),
.Y(n_6070)
);

OAI22xp5_ASAP7_75t_L g6071 ( 
.A1(n_5891),
.A2(n_3688),
.B1(n_3692),
.B2(n_3691),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5797),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_5812),
.Y(n_6073)
);

INVx3_ASAP7_75t_L g6074 ( 
.A(n_5703),
.Y(n_6074)
);

INVx2_ASAP7_75t_L g6075 ( 
.A(n_5846),
.Y(n_6075)
);

HB1xp67_ASAP7_75t_L g6076 ( 
.A(n_5946),
.Y(n_6076)
);

OAI22xp5_ASAP7_75t_SL g6077 ( 
.A1(n_5761),
.A2(n_4062),
.B1(n_4195),
.B2(n_4057),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5801),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5802),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_5855),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5805),
.Y(n_6081)
);

INVx2_ASAP7_75t_L g6082 ( 
.A(n_5703),
.Y(n_6082)
);

AND2x4_ASAP7_75t_L g6083 ( 
.A(n_5972),
.B(n_3924),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5703),
.Y(n_6084)
);

BUFx6f_ASAP7_75t_L g6085 ( 
.A(n_5710),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5808),
.Y(n_6086)
);

BUFx6f_ASAP7_75t_L g6087 ( 
.A(n_5842),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5561),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5810),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5814),
.Y(n_6090)
);

AND2x6_ASAP7_75t_L g6091 ( 
.A(n_5908),
.B(n_3680),
.Y(n_6091)
);

OAI22xp5_ASAP7_75t_SL g6092 ( 
.A1(n_5769),
.A2(n_4236),
.B1(n_4243),
.B2(n_4215),
.Y(n_6092)
);

INVx2_ASAP7_75t_SL g6093 ( 
.A(n_5929),
.Y(n_6093)
);

BUFx6f_ASAP7_75t_L g6094 ( 
.A(n_5843),
.Y(n_6094)
);

HB1xp67_ASAP7_75t_L g6095 ( 
.A(n_5686),
.Y(n_6095)
);

INVx2_ASAP7_75t_L g6096 ( 
.A(n_5571),
.Y(n_6096)
);

OA21x2_ASAP7_75t_L g6097 ( 
.A1(n_5887),
.A2(n_4255),
.B(n_4200),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5815),
.Y(n_6098)
);

INVx5_ASAP7_75t_L g6099 ( 
.A(n_5949),
.Y(n_6099)
);

BUFx6f_ASAP7_75t_L g6100 ( 
.A(n_5482),
.Y(n_6100)
);

INVx2_ASAP7_75t_L g6101 ( 
.A(n_5600),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5816),
.Y(n_6102)
);

NAND2xp5_ASAP7_75t_L g6103 ( 
.A(n_5882),
.B(n_4441),
.Y(n_6103)
);

INVx4_ASAP7_75t_L g6104 ( 
.A(n_5486),
.Y(n_6104)
);

INVxp67_ASAP7_75t_L g6105 ( 
.A(n_5931),
.Y(n_6105)
);

INVx2_ASAP7_75t_L g6106 ( 
.A(n_5697),
.Y(n_6106)
);

INVx4_ASAP7_75t_L g6107 ( 
.A(n_5489),
.Y(n_6107)
);

INVx5_ASAP7_75t_L g6108 ( 
.A(n_5983),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5889),
.B(n_4001),
.Y(n_6109)
);

NAND2xp5_ASAP7_75t_L g6110 ( 
.A(n_5672),
.B(n_4502),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_5919),
.B(n_5723),
.Y(n_6111)
);

OAI21x1_ASAP7_75t_L g6112 ( 
.A1(n_5888),
.A2(n_5893),
.B(n_5892),
.Y(n_6112)
);

BUFx6f_ASAP7_75t_L g6113 ( 
.A(n_5485),
.Y(n_6113)
);

CKINVDCx5p33_ASAP7_75t_R g6114 ( 
.A(n_5505),
.Y(n_6114)
);

AND2x4_ASAP7_75t_L g6115 ( 
.A(n_5985),
.B(n_3965),
.Y(n_6115)
);

INVx2_ASAP7_75t_L g6116 ( 
.A(n_5553),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5555),
.Y(n_6117)
);

INVx2_ASAP7_75t_L g6118 ( 
.A(n_5558),
.Y(n_6118)
);

INVx3_ASAP7_75t_L g6119 ( 
.A(n_5733),
.Y(n_6119)
);

BUFx8_ASAP7_75t_L g6120 ( 
.A(n_5969),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_5907),
.B(n_4512),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5818),
.Y(n_6122)
);

CKINVDCx5p33_ASAP7_75t_R g6123 ( 
.A(n_5508),
.Y(n_6123)
);

NAND2xp5_ASAP7_75t_L g6124 ( 
.A(n_5606),
.B(n_5707),
.Y(n_6124)
);

INVx2_ASAP7_75t_L g6125 ( 
.A(n_5559),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5819),
.Y(n_6126)
);

AND2x2_ASAP7_75t_L g6127 ( 
.A(n_5898),
.B(n_4001),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5821),
.Y(n_6128)
);

CKINVDCx5p33_ASAP7_75t_R g6129 ( 
.A(n_5513),
.Y(n_6129)
);

AND2x4_ASAP7_75t_L g6130 ( 
.A(n_5642),
.B(n_3990),
.Y(n_6130)
);

BUFx2_ASAP7_75t_L g6131 ( 
.A(n_5619),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_5564),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_5565),
.Y(n_6133)
);

AOI22xp5_ASAP7_75t_SL g6134 ( 
.A1(n_5932),
.A2(n_4289),
.B1(n_4297),
.B2(n_4275),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_5567),
.Y(n_6135)
);

BUFx6f_ASAP7_75t_L g6136 ( 
.A(n_5487),
.Y(n_6136)
);

OA21x2_ASAP7_75t_L g6137 ( 
.A1(n_5894),
.A2(n_4800),
.B(n_4661),
.Y(n_6137)
);

BUFx6f_ASAP7_75t_L g6138 ( 
.A(n_5490),
.Y(n_6138)
);

INVx3_ASAP7_75t_L g6139 ( 
.A(n_5491),
.Y(n_6139)
);

CKINVDCx16_ASAP7_75t_R g6140 ( 
.A(n_5716),
.Y(n_6140)
);

AOI22xp5_ASAP7_75t_L g6141 ( 
.A1(n_5948),
.A2(n_3772),
.B1(n_3859),
.B2(n_3750),
.Y(n_6141)
);

NAND2xp5_ASAP7_75t_L g6142 ( 
.A(n_5708),
.B(n_4875),
.Y(n_6142)
);

BUFx6f_ASAP7_75t_L g6143 ( 
.A(n_5987),
.Y(n_6143)
);

BUFx6f_ASAP7_75t_L g6144 ( 
.A(n_5493),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5826),
.Y(n_6145)
);

INVx3_ASAP7_75t_L g6146 ( 
.A(n_5938),
.Y(n_6146)
);

BUFx2_ASAP7_75t_L g6147 ( 
.A(n_5634),
.Y(n_6147)
);

BUFx3_ASAP7_75t_L g6148 ( 
.A(n_5661),
.Y(n_6148)
);

OAI21x1_ASAP7_75t_L g6149 ( 
.A1(n_5900),
.A2(n_5000),
.B(n_4949),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_5500),
.B(n_4212),
.Y(n_6150)
);

BUFx6f_ASAP7_75t_L g6151 ( 
.A(n_5941),
.Y(n_6151)
);

OA21x2_ASAP7_75t_L g6152 ( 
.A1(n_5901),
.A2(n_3819),
.B(n_3817),
.Y(n_6152)
);

AND2x4_ASAP7_75t_L g6153 ( 
.A(n_5637),
.B(n_4027),
.Y(n_6153)
);

OAI21x1_ASAP7_75t_L g6154 ( 
.A1(n_5902),
.A2(n_3758),
.B(n_3741),
.Y(n_6154)
);

AOI22xp5_ASAP7_75t_L g6155 ( 
.A1(n_5953),
.A2(n_3946),
.B1(n_3992),
.B2(n_3929),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5830),
.Y(n_6156)
);

OAI22xp5_ASAP7_75t_L g6157 ( 
.A1(n_5891),
.A2(n_5914),
.B1(n_5915),
.B2(n_5913),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5832),
.Y(n_6158)
);

INVx2_ASAP7_75t_L g6159 ( 
.A(n_5570),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5833),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_5573),
.Y(n_6161)
);

OA21x2_ASAP7_75t_L g6162 ( 
.A1(n_5713),
.A2(n_3823),
.B(n_3821),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_5574),
.Y(n_6163)
);

AND2x4_ASAP7_75t_L g6164 ( 
.A(n_5726),
.B(n_4090),
.Y(n_6164)
);

INVxp67_ASAP7_75t_L g6165 ( 
.A(n_5911),
.Y(n_6165)
);

CKINVDCx5p33_ASAP7_75t_R g6166 ( 
.A(n_5515),
.Y(n_6166)
);

INVx2_ASAP7_75t_L g6167 ( 
.A(n_5575),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5836),
.Y(n_6168)
);

AND2x4_ASAP7_75t_L g6169 ( 
.A(n_5728),
.B(n_4135),
.Y(n_6169)
);

INVx3_ASAP7_75t_L g6170 ( 
.A(n_5950),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_5577),
.Y(n_6171)
);

INVx4_ASAP7_75t_L g6172 ( 
.A(n_5519),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_5581),
.Y(n_6173)
);

AND2x4_ASAP7_75t_L g6174 ( 
.A(n_5693),
.B(n_4141),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5839),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5582),
.Y(n_6176)
);

AND2x4_ASAP7_75t_L g6177 ( 
.A(n_5916),
.B(n_4315),
.Y(n_6177)
);

AOI22xp5_ASAP7_75t_SL g6178 ( 
.A1(n_5774),
.A2(n_4342),
.B1(n_4355),
.B2(n_4322),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5847),
.Y(n_6179)
);

INVx6_ASAP7_75t_L g6180 ( 
.A(n_5780),
.Y(n_6180)
);

INVx2_ASAP7_75t_L g6181 ( 
.A(n_5584),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5849),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5851),
.Y(n_6183)
);

BUFx3_ASAP7_75t_L g6184 ( 
.A(n_5663),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_5854),
.Y(n_6185)
);

OAI22x1_ASAP7_75t_L g6186 ( 
.A1(n_5986),
.A2(n_4007),
.B1(n_4060),
.B2(n_3993),
.Y(n_6186)
);

INVx2_ASAP7_75t_L g6187 ( 
.A(n_5585),
.Y(n_6187)
);

BUFx8_ASAP7_75t_SL g6188 ( 
.A(n_5533),
.Y(n_6188)
);

OAI22xp33_ASAP7_75t_R g6189 ( 
.A1(n_5930),
.A2(n_4164),
.B1(n_4190),
.B2(n_4065),
.Y(n_6189)
);

INVx3_ASAP7_75t_L g6190 ( 
.A(n_5951),
.Y(n_6190)
);

BUFx12f_ASAP7_75t_L g6191 ( 
.A(n_5780),
.Y(n_6191)
);

INVx2_ASAP7_75t_L g6192 ( 
.A(n_5586),
.Y(n_6192)
);

BUFx2_ASAP7_75t_L g6193 ( 
.A(n_5651),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_5858),
.Y(n_6194)
);

BUFx6f_ASAP7_75t_L g6195 ( 
.A(n_5984),
.Y(n_6195)
);

OAI22xp5_ASAP7_75t_SL g6196 ( 
.A1(n_5657),
.A2(n_4397),
.B1(n_4433),
.B2(n_4360),
.Y(n_6196)
);

AND2x2_ASAP7_75t_L g6197 ( 
.A(n_5943),
.B(n_4212),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_5588),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_5589),
.Y(n_6199)
);

OAI21x1_ASAP7_75t_L g6200 ( 
.A1(n_5718),
.A2(n_3830),
.B(n_3768),
.Y(n_6200)
);

CKINVDCx16_ASAP7_75t_R g6201 ( 
.A(n_5790),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_5590),
.Y(n_6202)
);

CKINVDCx6p67_ASAP7_75t_R g6203 ( 
.A(n_5796),
.Y(n_6203)
);

INVx6_ASAP7_75t_L g6204 ( 
.A(n_5825),
.Y(n_6204)
);

NAND2xp5_ASAP7_75t_L g6205 ( 
.A(n_5719),
.B(n_4371),
.Y(n_6205)
);

BUFx12f_ASAP7_75t_L g6206 ( 
.A(n_5711),
.Y(n_6206)
);

AOI22xp5_ASAP7_75t_L g6207 ( 
.A1(n_5587),
.A2(n_4447),
.B1(n_4473),
.B2(n_4419),
.Y(n_6207)
);

NOR2x1_ASAP7_75t_L g6208 ( 
.A(n_5897),
.B(n_4533),
.Y(n_6208)
);

BUFx6f_ASAP7_75t_L g6209 ( 
.A(n_5982),
.Y(n_6209)
);

BUFx6f_ASAP7_75t_L g6210 ( 
.A(n_5952),
.Y(n_6210)
);

CKINVDCx5p33_ASAP7_75t_R g6211 ( 
.A(n_5530),
.Y(n_6211)
);

INVx2_ASAP7_75t_L g6212 ( 
.A(n_5594),
.Y(n_6212)
);

BUFx6f_ASAP7_75t_L g6213 ( 
.A(n_5981),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_L g6214 ( 
.A(n_5722),
.B(n_4524),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_5729),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_5596),
.Y(n_6216)
);

AOI22xp5_ASAP7_75t_L g6217 ( 
.A1(n_5592),
.A2(n_5597),
.B1(n_5917),
.B2(n_5906),
.Y(n_6217)
);

INVx2_ASAP7_75t_L g6218 ( 
.A(n_5598),
.Y(n_6218)
);

HB1xp67_ASAP7_75t_L g6219 ( 
.A(n_5643),
.Y(n_6219)
);

BUFx2_ASAP7_75t_L g6220 ( 
.A(n_5709),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_5532),
.Y(n_6221)
);

CKINVDCx5p33_ASAP7_75t_R g6222 ( 
.A(n_5535),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5731),
.Y(n_6223)
);

INVx3_ASAP7_75t_L g6224 ( 
.A(n_5956),
.Y(n_6224)
);

AND2x4_ASAP7_75t_L g6225 ( 
.A(n_5730),
.B(n_4627),
.Y(n_6225)
);

INVx2_ASAP7_75t_L g6226 ( 
.A(n_5599),
.Y(n_6226)
);

INVx2_ASAP7_75t_L g6227 ( 
.A(n_5601),
.Y(n_6227)
);

BUFx2_ASAP7_75t_L g6228 ( 
.A(n_5738),
.Y(n_6228)
);

INVx1_ASAP7_75t_SL g6229 ( 
.A(n_5536),
.Y(n_6229)
);

AND2x4_ASAP7_75t_L g6230 ( 
.A(n_5735),
.B(n_4663),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_5732),
.B(n_4766),
.Y(n_6231)
);

NAND2xp5_ASAP7_75t_SL g6232 ( 
.A(n_5537),
.B(n_5539),
.Y(n_6232)
);

BUFx12f_ASAP7_75t_L g6233 ( 
.A(n_5715),
.Y(n_6233)
);

BUFx8_ASAP7_75t_L g6234 ( 
.A(n_5724),
.Y(n_6234)
);

INVx4_ASAP7_75t_L g6235 ( 
.A(n_5548),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_5734),
.Y(n_6236)
);

BUFx6f_ASAP7_75t_L g6237 ( 
.A(n_5967),
.Y(n_6237)
);

OAI22xp5_ASAP7_75t_L g6238 ( 
.A1(n_5903),
.A2(n_5831),
.B1(n_5920),
.B2(n_5918),
.Y(n_6238)
);

OA21x2_ASAP7_75t_L g6239 ( 
.A1(n_5737),
.A2(n_3832),
.B(n_3827),
.Y(n_6239)
);

INVx1_ASAP7_75t_L g6240 ( 
.A(n_5739),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5740),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5603),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_5604),
.Y(n_6243)
);

BUFx6f_ASAP7_75t_L g6244 ( 
.A(n_5968),
.Y(n_6244)
);

HB1xp67_ASAP7_75t_L g6245 ( 
.A(n_5683),
.Y(n_6245)
);

BUFx6f_ASAP7_75t_L g6246 ( 
.A(n_5970),
.Y(n_6246)
);

BUFx2_ASAP7_75t_L g6247 ( 
.A(n_5556),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5607),
.Y(n_6248)
);

BUFx3_ASAP7_75t_L g6249 ( 
.A(n_5695),
.Y(n_6249)
);

OAI22xp5_ASAP7_75t_SL g6250 ( 
.A1(n_5647),
.A2(n_4475),
.B1(n_4487),
.B2(n_4469),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5741),
.Y(n_6251)
);

INVx2_ASAP7_75t_L g6252 ( 
.A(n_5610),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5742),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_5743),
.B(n_4978),
.Y(n_6254)
);

BUFx6f_ASAP7_75t_L g6255 ( 
.A(n_5971),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5744),
.Y(n_6256)
);

NAND2xp5_ASAP7_75t_L g6257 ( 
.A(n_5747),
.B(n_5032),
.Y(n_6257)
);

OAI22xp5_ASAP7_75t_L g6258 ( 
.A1(n_5926),
.A2(n_3696),
.B1(n_3697),
.B2(n_3695),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_5613),
.Y(n_6259)
);

INVx2_ASAP7_75t_L g6260 ( 
.A(n_5614),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5615),
.Y(n_6261)
);

BUFx6f_ASAP7_75t_L g6262 ( 
.A(n_5973),
.Y(n_6262)
);

NOR2xp33_ASAP7_75t_L g6263 ( 
.A(n_5560),
.B(n_5035),
.Y(n_6263)
);

INVx3_ASAP7_75t_L g6264 ( 
.A(n_5974),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5748),
.Y(n_6265)
);

BUFx8_ASAP7_75t_L g6266 ( 
.A(n_5563),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_5750),
.B(n_4136),
.Y(n_6267)
);

BUFx6f_ASAP7_75t_L g6268 ( 
.A(n_5977),
.Y(n_6268)
);

NAND2xp5_ASAP7_75t_L g6269 ( 
.A(n_5754),
.B(n_3835),
.Y(n_6269)
);

NAND2xp5_ASAP7_75t_L g6270 ( 
.A(n_5800),
.B(n_3926),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5864),
.Y(n_6271)
);

AND2x4_ASAP7_75t_L g6272 ( 
.A(n_5746),
.B(n_3838),
.Y(n_6272)
);

AOI22xp5_ASAP7_75t_L g6273 ( 
.A1(n_5562),
.A2(n_5568),
.B1(n_5569),
.B2(n_5566),
.Y(n_6273)
);

HB1xp67_ASAP7_75t_L g6274 ( 
.A(n_5706),
.Y(n_6274)
);

INVx5_ASAP7_75t_L g6275 ( 
.A(n_5813),
.Y(n_6275)
);

OA21x2_ASAP7_75t_L g6276 ( 
.A1(n_5927),
.A2(n_3840),
.B(n_3839),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_5865),
.Y(n_6277)
);

HB1xp67_ASAP7_75t_L g6278 ( 
.A(n_5736),
.Y(n_6278)
);

BUFx6f_ASAP7_75t_L g6279 ( 
.A(n_5494),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_5866),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_5800),
.B(n_3934),
.Y(n_6281)
);

BUFx12f_ASAP7_75t_L g6282 ( 
.A(n_5721),
.Y(n_6282)
);

AND2x4_ASAP7_75t_L g6283 ( 
.A(n_5791),
.B(n_3842),
.Y(n_6283)
);

INVx1_ASAP7_75t_L g6284 ( 
.A(n_5868),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_5616),
.Y(n_6285)
);

OA21x2_ASAP7_75t_L g6286 ( 
.A1(n_5928),
.A2(n_3846),
.B(n_3843),
.Y(n_6286)
);

AND2x4_ASAP7_75t_L g6287 ( 
.A(n_5822),
.B(n_3850),
.Y(n_6287)
);

NAND2xp5_ASAP7_75t_L g6288 ( 
.A(n_5800),
.B(n_3951),
.Y(n_6288)
);

BUFx6f_ASAP7_75t_L g6289 ( 
.A(n_5495),
.Y(n_6289)
);

BUFx12f_ASAP7_75t_L g6290 ( 
.A(n_5727),
.Y(n_6290)
);

NAND2xp5_ASAP7_75t_L g6291 ( 
.A(n_5800),
.B(n_3958),
.Y(n_6291)
);

INVx5_ASAP7_75t_L g6292 ( 
.A(n_5783),
.Y(n_6292)
);

OA21x2_ASAP7_75t_L g6293 ( 
.A1(n_5824),
.A2(n_5852),
.B(n_5840),
.Y(n_6293)
);

INVx2_ASAP7_75t_L g6294 ( 
.A(n_5618),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_5620),
.Y(n_6295)
);

AND2x4_ASAP7_75t_L g6296 ( 
.A(n_5873),
.B(n_3855),
.Y(n_6296)
);

INVx3_ASAP7_75t_L g6297 ( 
.A(n_5496),
.Y(n_6297)
);

INVx2_ASAP7_75t_L g6298 ( 
.A(n_5621),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_5870),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5871),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5757),
.Y(n_6301)
);

INVx3_ASAP7_75t_L g6302 ( 
.A(n_5499),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_5800),
.B(n_3988),
.Y(n_6303)
);

BUFx8_ASAP7_75t_L g6304 ( 
.A(n_5856),
.Y(n_6304)
);

OA21x2_ASAP7_75t_L g6305 ( 
.A1(n_5876),
.A2(n_3863),
.B(n_3856),
.Y(n_6305)
);

INVxp67_ASAP7_75t_L g6306 ( 
.A(n_5933),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_5622),
.Y(n_6307)
);

INVx2_ASAP7_75t_L g6308 ( 
.A(n_5623),
.Y(n_6308)
);

OA21x2_ASAP7_75t_L g6309 ( 
.A1(n_5758),
.A2(n_3866),
.B(n_3865),
.Y(n_6309)
);

BUFx6f_ASAP7_75t_L g6310 ( 
.A(n_5502),
.Y(n_6310)
);

BUFx2_ASAP7_75t_L g6311 ( 
.A(n_5751),
.Y(n_6311)
);

NOR2xp33_ASAP7_75t_L g6312 ( 
.A(n_5576),
.B(n_3699),
.Y(n_6312)
);

NAND2xp5_ASAP7_75t_L g6313 ( 
.A(n_5759),
.B(n_4023),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_L g6314 ( 
.A(n_5624),
.B(n_4029),
.Y(n_6314)
);

CKINVDCx5p33_ASAP7_75t_R g6315 ( 
.A(n_5579),
.Y(n_6315)
);

CKINVDCx6p67_ASAP7_75t_R g6316 ( 
.A(n_5648),
.Y(n_6316)
);

INVx2_ASAP7_75t_L g6317 ( 
.A(n_5628),
.Y(n_6317)
);

INVx2_ASAP7_75t_L g6318 ( 
.A(n_5629),
.Y(n_6318)
);

INVx2_ASAP7_75t_L g6319 ( 
.A(n_5630),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_5631),
.Y(n_6320)
);

INVx2_ASAP7_75t_L g6321 ( 
.A(n_5633),
.Y(n_6321)
);

BUFx8_ASAP7_75t_L g6322 ( 
.A(n_5935),
.Y(n_6322)
);

INVx4_ASAP7_75t_L g6323 ( 
.A(n_5580),
.Y(n_6323)
);

AOI22xp5_ASAP7_75t_L g6324 ( 
.A1(n_5583),
.A2(n_5612),
.B1(n_5617),
.B2(n_5602),
.Y(n_6324)
);

INVx2_ASAP7_75t_L g6325 ( 
.A(n_5635),
.Y(n_6325)
);

INVx3_ASAP7_75t_L g6326 ( 
.A(n_5509),
.Y(n_6326)
);

AND2x2_ASAP7_75t_SL g6327 ( 
.A(n_5497),
.B(n_4032),
.Y(n_6327)
);

INVx2_ASAP7_75t_L g6328 ( 
.A(n_5636),
.Y(n_6328)
);

AND2x4_ASAP7_75t_L g6329 ( 
.A(n_5936),
.B(n_3870),
.Y(n_6329)
);

BUFx6f_ASAP7_75t_L g6330 ( 
.A(n_5510),
.Y(n_6330)
);

AND2x2_ASAP7_75t_SL g6331 ( 
.A(n_5504),
.B(n_5507),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_5639),
.Y(n_6332)
);

AND2x2_ASAP7_75t_SL g6333 ( 
.A(n_5529),
.B(n_4044),
.Y(n_6333)
);

AND2x4_ASAP7_75t_L g6334 ( 
.A(n_5514),
.B(n_3877),
.Y(n_6334)
);

BUFx6f_ASAP7_75t_L g6335 ( 
.A(n_5516),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_5640),
.B(n_4059),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_5644),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_5646),
.Y(n_6338)
);

NAND2xp5_ASAP7_75t_L g6339 ( 
.A(n_5649),
.B(n_4107),
.Y(n_6339)
);

INVx5_ASAP7_75t_L g6340 ( 
.A(n_5518),
.Y(n_6340)
);

INVx3_ASAP7_75t_L g6341 ( 
.A(n_5522),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_L g6342 ( 
.A(n_5652),
.B(n_4117),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_5654),
.Y(n_6343)
);

INVx2_ASAP7_75t_L g6344 ( 
.A(n_5656),
.Y(n_6344)
);

AOI22xp5_ASAP7_75t_L g6345 ( 
.A1(n_5627),
.A2(n_4545),
.B1(n_4574),
.B2(n_4541),
.Y(n_6345)
);

INVx3_ASAP7_75t_L g6346 ( 
.A(n_5523),
.Y(n_6346)
);

BUFx6f_ASAP7_75t_L g6347 ( 
.A(n_5524),
.Y(n_6347)
);

AND2x4_ASAP7_75t_L g6348 ( 
.A(n_5526),
.B(n_3880),
.Y(n_6348)
);

AND2x6_ASAP7_75t_L g6349 ( 
.A(n_5531),
.B(n_4587),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_5659),
.Y(n_6350)
);

NOR2xp33_ASAP7_75t_L g6351 ( 
.A(n_5638),
.B(n_3700),
.Y(n_6351)
);

BUFx6f_ASAP7_75t_L g6352 ( 
.A(n_5660),
.Y(n_6352)
);

OAI21x1_ASAP7_75t_L g6353 ( 
.A1(n_5662),
.A2(n_4172),
.B(n_4127),
.Y(n_6353)
);

INVx2_ASAP7_75t_L g6354 ( 
.A(n_5664),
.Y(n_6354)
);

AND2x4_ASAP7_75t_L g6355 ( 
.A(n_5792),
.B(n_3884),
.Y(n_6355)
);

BUFx2_ASAP7_75t_L g6356 ( 
.A(n_5778),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_5665),
.Y(n_6357)
);

BUFx6f_ASAP7_75t_L g6358 ( 
.A(n_5666),
.Y(n_6358)
);

AND2x4_ASAP7_75t_L g6359 ( 
.A(n_5823),
.B(n_3898),
.Y(n_6359)
);

HB1xp67_ASAP7_75t_L g6360 ( 
.A(n_5835),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5669),
.Y(n_6361)
);

NAND2xp5_ASAP7_75t_SL g6362 ( 
.A(n_5653),
.B(n_3701),
.Y(n_6362)
);

AND2x4_ASAP7_75t_L g6363 ( 
.A(n_5869),
.B(n_3900),
.Y(n_6363)
);

INVx3_ASAP7_75t_L g6364 ( 
.A(n_5675),
.Y(n_6364)
);

AND2x4_ASAP7_75t_L g6365 ( 
.A(n_5895),
.B(n_3902),
.Y(n_6365)
);

INVx2_ASAP7_75t_L g6366 ( 
.A(n_5677),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_5679),
.Y(n_6367)
);

AND2x2_ASAP7_75t_L g6368 ( 
.A(n_5717),
.B(n_4242),
.Y(n_6368)
);

BUFx2_ASAP7_75t_L g6369 ( 
.A(n_5793),
.Y(n_6369)
);

AOI22xp5_ASAP7_75t_L g6370 ( 
.A1(n_5667),
.A2(n_4647),
.B1(n_4662),
.B2(n_4631),
.Y(n_6370)
);

INVx3_ASAP7_75t_L g6371 ( 
.A(n_5681),
.Y(n_6371)
);

OAI22x1_ASAP7_75t_R g6372 ( 
.A1(n_5554),
.A2(n_4552),
.B1(n_4560),
.B2(n_4535),
.Y(n_6372)
);

INVx6_ASAP7_75t_L g6373 ( 
.A(n_5591),
.Y(n_6373)
);

INVx6_ASAP7_75t_L g6374 ( 
.A(n_5605),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_5682),
.Y(n_6375)
);

NOR2xp33_ASAP7_75t_L g6376 ( 
.A(n_5671),
.B(n_3702),
.Y(n_6376)
);

BUFx12f_ASAP7_75t_L g6377 ( 
.A(n_5745),
.Y(n_6377)
);

INVx6_ASAP7_75t_L g6378 ( 
.A(n_5608),
.Y(n_6378)
);

CKINVDCx11_ASAP7_75t_R g6379 ( 
.A(n_5625),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_5687),
.Y(n_6380)
);

BUFx6f_ASAP7_75t_L g6381 ( 
.A(n_5688),
.Y(n_6381)
);

CKINVDCx6p67_ASAP7_75t_R g6382 ( 
.A(n_5794),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_5689),
.Y(n_6383)
);

HB1xp67_ASAP7_75t_L g6384 ( 
.A(n_5910),
.Y(n_6384)
);

BUFx12f_ASAP7_75t_L g6385 ( 
.A(n_5752),
.Y(n_6385)
);

AND2x6_ASAP7_75t_L g6386 ( 
.A(n_5691),
.B(n_4671),
.Y(n_6386)
);

INVx2_ASAP7_75t_L g6387 ( 
.A(n_5692),
.Y(n_6387)
);

BUFx6f_ASAP7_75t_L g6388 ( 
.A(n_5694),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_5698),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_5700),
.Y(n_6390)
);

BUFx12f_ASAP7_75t_L g6391 ( 
.A(n_5765),
.Y(n_6391)
);

BUFx2_ASAP7_75t_L g6392 ( 
.A(n_5817),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_5762),
.Y(n_6393)
);

INVx4_ASAP7_75t_L g6394 ( 
.A(n_5673),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_5701),
.Y(n_6395)
);

BUFx3_ASAP7_75t_L g6396 ( 
.A(n_5838),
.Y(n_6396)
);

INVxp67_ASAP7_75t_L g6397 ( 
.A(n_5650),
.Y(n_6397)
);

AND2x2_ASAP7_75t_SL g6398 ( 
.A(n_5655),
.B(n_4181),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_5702),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_5704),
.Y(n_6400)
);

BUFx3_ASAP7_75t_L g6401 ( 
.A(n_5841),
.Y(n_6401)
);

BUFx6f_ASAP7_75t_L g6402 ( 
.A(n_5705),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_5534),
.Y(n_6403)
);

HB1xp67_ASAP7_75t_L g6404 ( 
.A(n_5803),
.Y(n_6404)
);

OAI21x1_ASAP7_75t_L g6405 ( 
.A1(n_5538),
.A2(n_4249),
.B(n_4213),
.Y(n_6405)
);

INVx3_ASAP7_75t_L g6406 ( 
.A(n_5859),
.Y(n_6406)
);

NAND2xp5_ASAP7_75t_L g6407 ( 
.A(n_5540),
.B(n_4269),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_5543),
.B(n_4272),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_5860),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5544),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_5545),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_SL g6412 ( 
.A(n_5674),
.B(n_3705),
.Y(n_6412)
);

AND2x4_ASAP7_75t_L g6413 ( 
.A(n_5756),
.B(n_3904),
.Y(n_6413)
);

CKINVDCx5p33_ASAP7_75t_R g6414 ( 
.A(n_5685),
.Y(n_6414)
);

BUFx3_ASAP7_75t_L g6415 ( 
.A(n_5861),
.Y(n_6415)
);

BUFx12f_ASAP7_75t_L g6416 ( 
.A(n_5781),
.Y(n_6416)
);

HB1xp67_ASAP7_75t_L g6417 ( 
.A(n_5668),
.Y(n_6417)
);

BUFx6f_ASAP7_75t_L g6418 ( 
.A(n_5546),
.Y(n_6418)
);

BUFx8_ASAP7_75t_L g6419 ( 
.A(n_5626),
.Y(n_6419)
);

INVx6_ASAP7_75t_L g6420 ( 
.A(n_5641),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5547),
.Y(n_6421)
);

AND2x4_ASAP7_75t_L g6422 ( 
.A(n_5766),
.B(n_3913),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_5549),
.Y(n_6423)
);

INVx2_ASAP7_75t_L g6424 ( 
.A(n_5550),
.Y(n_6424)
);

AND2x4_ASAP7_75t_L g6425 ( 
.A(n_5850),
.B(n_3920),
.Y(n_6425)
);

AND2x4_ASAP7_75t_L g6426 ( 
.A(n_5857),
.B(n_3922),
.Y(n_6426)
);

OAI22x1_ASAP7_75t_L g6427 ( 
.A1(n_5934),
.A2(n_4826),
.B1(n_4869),
.B2(n_4673),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_5551),
.Y(n_6428)
);

OA21x2_ASAP7_75t_L g6429 ( 
.A1(n_5552),
.A2(n_3925),
.B(n_3923),
.Y(n_6429)
);

OAI21x1_ASAP7_75t_L g6430 ( 
.A1(n_5670),
.A2(n_4383),
.B(n_4278),
.Y(n_6430)
);

OAI22xp5_ASAP7_75t_L g6431 ( 
.A1(n_5690),
.A2(n_3707),
.B1(n_3709),
.B2(n_3706),
.Y(n_6431)
);

NAND2xp5_ASAP7_75t_L g6432 ( 
.A(n_5699),
.B(n_4443),
.Y(n_6432)
);

BUFx6f_ASAP7_75t_L g6433 ( 
.A(n_5785),
.Y(n_6433)
);

BUFx6f_ASAP7_75t_L g6434 ( 
.A(n_5789),
.Y(n_6434)
);

BUFx2_ASAP7_75t_L g6435 ( 
.A(n_5875),
.Y(n_6435)
);

BUFx6f_ASAP7_75t_L g6436 ( 
.A(n_5799),
.Y(n_6436)
);

INVx2_ASAP7_75t_L g6437 ( 
.A(n_5937),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5678),
.Y(n_6438)
);

BUFx2_ASAP7_75t_L g6439 ( 
.A(n_5879),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_5940),
.Y(n_6440)
);

AOI22xp5_ASAP7_75t_L g6441 ( 
.A1(n_5942),
.A2(n_4910),
.B1(n_3720),
.B2(n_3721),
.Y(n_6441)
);

NOR2x1_ASAP7_75t_L g6442 ( 
.A(n_5881),
.B(n_4653),
.Y(n_6442)
);

INVx2_ASAP7_75t_L g6443 ( 
.A(n_5954),
.Y(n_6443)
);

AND2x4_ASAP7_75t_L g6444 ( 
.A(n_5696),
.B(n_3927),
.Y(n_6444)
);

INVx4_ASAP7_75t_L g6445 ( 
.A(n_5957),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_5749),
.Y(n_6446)
);

BUFx12f_ASAP7_75t_L g6447 ( 
.A(n_5806),
.Y(n_6447)
);

INVx2_ASAP7_75t_L g6448 ( 
.A(n_5959),
.Y(n_6448)
);

BUFx6f_ASAP7_75t_L g6449 ( 
.A(n_5809),
.Y(n_6449)
);

BUFx6f_ASAP7_75t_L g6450 ( 
.A(n_5811),
.Y(n_6450)
);

NAND2xp5_ASAP7_75t_L g6451 ( 
.A(n_5965),
.B(n_4450),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_5961),
.Y(n_6452)
);

NAND2xp5_ASAP7_75t_L g6453 ( 
.A(n_5975),
.B(n_4451),
.Y(n_6453)
);

INVx5_ASAP7_75t_L g6454 ( 
.A(n_5542),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_5978),
.Y(n_6455)
);

INVx2_ASAP7_75t_L g6456 ( 
.A(n_5820),
.Y(n_6456)
);

OA21x2_ASAP7_75t_L g6457 ( 
.A1(n_5827),
.A2(n_3937),
.B(n_3931),
.Y(n_6457)
);

INVx6_ASAP7_75t_L g6458 ( 
.A(n_5557),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5829),
.Y(n_6459)
);

OAI22xp5_ASAP7_75t_SL g6460 ( 
.A1(n_5899),
.A2(n_4565),
.B1(n_4571),
.B2(n_4562),
.Y(n_6460)
);

OAI22xp5_ASAP7_75t_L g6461 ( 
.A1(n_5834),
.A2(n_3725),
.B1(n_3731),
.B2(n_3717),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_L g6462 ( 
.A(n_5844),
.B(n_4497),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5853),
.Y(n_6463)
);

INVx2_ASAP7_75t_L g6464 ( 
.A(n_5862),
.Y(n_6464)
);

INVx2_ASAP7_75t_L g6465 ( 
.A(n_5863),
.Y(n_6465)
);

AND2x2_ASAP7_75t_L g6466 ( 
.A(n_5867),
.B(n_4242),
.Y(n_6466)
);

OAI22xp5_ASAP7_75t_L g6467 ( 
.A1(n_5872),
.A2(n_3734),
.B1(n_3736),
.B2(n_3732),
.Y(n_6467)
);

NOR2xp33_ASAP7_75t_SL g6468 ( 
.A(n_5632),
.B(n_4578),
.Y(n_6468)
);

AOI22x1_ASAP7_75t_SL g6469 ( 
.A1(n_5480),
.A2(n_4589),
.B1(n_4609),
.B2(n_4586),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_5874),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_5890),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_5904),
.Y(n_6472)
);

BUFx6f_ASAP7_75t_L g6473 ( 
.A(n_5909),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_5804),
.B(n_4546),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_5807),
.Y(n_6475)
);

BUFx3_ASAP7_75t_L g6476 ( 
.A(n_5905),
.Y(n_6476)
);

AND2x2_ASAP7_75t_L g6477 ( 
.A(n_5525),
.B(n_4464),
.Y(n_6477)
);

BUFx6f_ASAP7_75t_L g6478 ( 
.A(n_5658),
.Y(n_6478)
);

OA21x2_ASAP7_75t_L g6479 ( 
.A1(n_5837),
.A2(n_3960),
.B(n_3948),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5845),
.Y(n_6480)
);

INVx2_ASAP7_75t_L g6481 ( 
.A(n_5481),
.Y(n_6481)
);

OA21x2_ASAP7_75t_L g6482 ( 
.A1(n_5921),
.A2(n_3971),
.B(n_3968),
.Y(n_6482)
);

CKINVDCx6p67_ASAP7_75t_R g6483 ( 
.A(n_5511),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_5680),
.Y(n_6484)
);

INVx2_ASAP7_75t_L g6485 ( 
.A(n_5517),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_5578),
.Y(n_6486)
);

BUFx6f_ASAP7_75t_L g6487 ( 
.A(n_5521),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_5939),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_5945),
.Y(n_6489)
);

OA21x2_ASAP7_75t_L g6490 ( 
.A1(n_5976),
.A2(n_3975),
.B(n_3974),
.Y(n_6490)
);

BUFx6f_ASAP7_75t_L g6491 ( 
.A(n_5962),
.Y(n_6491)
);

XOR2xp5_ASAP7_75t_L g6492 ( 
.A(n_5963),
.B(n_4621),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_5979),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_5760),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_5760),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_5760),
.Y(n_6496)
);

AND2x4_ASAP7_75t_L g6497 ( 
.A(n_5955),
.B(n_3977),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_5760),
.Y(n_6498)
);

INVx2_ASAP7_75t_SL g6499 ( 
.A(n_5922),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_5877),
.B(n_4569),
.Y(n_6500)
);

BUFx6f_ASAP7_75t_L g6501 ( 
.A(n_5609),
.Y(n_6501)
);

BUFx12f_ASAP7_75t_L g6502 ( 
.A(n_5922),
.Y(n_6502)
);

AND2x2_ASAP7_75t_L g6503 ( 
.A(n_5686),
.B(n_4464),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_5760),
.Y(n_6504)
);

NAND2xp5_ASAP7_75t_SL g6505 ( 
.A(n_5922),
.B(n_3739),
.Y(n_6505)
);

BUFx6f_ASAP7_75t_L g6506 ( 
.A(n_5609),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5492),
.Y(n_6507)
);

CKINVDCx5p33_ASAP7_75t_R g6508 ( 
.A(n_5479),
.Y(n_6508)
);

BUFx12f_ASAP7_75t_L g6509 ( 
.A(n_5922),
.Y(n_6509)
);

OAI22x1_ASAP7_75t_L g6510 ( 
.A1(n_5922),
.A2(n_3743),
.B1(n_3747),
.B2(n_3742),
.Y(n_6510)
);

CKINVDCx5p33_ASAP7_75t_R g6511 ( 
.A(n_5479),
.Y(n_6511)
);

INVx4_ASAP7_75t_L g6512 ( 
.A(n_5479),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_5492),
.Y(n_6513)
);

CKINVDCx5p33_ASAP7_75t_R g6514 ( 
.A(n_5479),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_5760),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_5760),
.Y(n_6516)
);

AND2x4_ASAP7_75t_L g6517 ( 
.A(n_5955),
.B(n_3980),
.Y(n_6517)
);

BUFx3_ASAP7_75t_L g6518 ( 
.A(n_5955),
.Y(n_6518)
);

INVx3_ASAP7_75t_L g6519 ( 
.A(n_5609),
.Y(n_6519)
);

BUFx6f_ASAP7_75t_L g6520 ( 
.A(n_5609),
.Y(n_6520)
);

OAI22xp5_ASAP7_75t_L g6521 ( 
.A1(n_5645),
.A2(n_3749),
.B1(n_3751),
.B2(n_3748),
.Y(n_6521)
);

BUFx6f_ASAP7_75t_L g6522 ( 
.A(n_5609),
.Y(n_6522)
);

BUFx6f_ASAP7_75t_L g6523 ( 
.A(n_5609),
.Y(n_6523)
);

INVx3_ASAP7_75t_L g6524 ( 
.A(n_5609),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_5760),
.Y(n_6525)
);

AND2x6_ASAP7_75t_L g6526 ( 
.A(n_5908),
.B(n_3983),
.Y(n_6526)
);

AOI22xp5_ASAP7_75t_L g6527 ( 
.A1(n_5645),
.A2(n_3756),
.B1(n_3757),
.B2(n_3755),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_SL g6528 ( 
.A(n_5922),
.B(n_3764),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_5760),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_5492),
.Y(n_6530)
);

AND2x4_ASAP7_75t_L g6531 ( 
.A(n_5955),
.B(n_3984),
.Y(n_6531)
);

AND2x4_ASAP7_75t_L g6532 ( 
.A(n_5955),
.B(n_3986),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_5492),
.Y(n_6533)
);

INVx3_ASAP7_75t_L g6534 ( 
.A(n_5609),
.Y(n_6534)
);

BUFx2_ASAP7_75t_L g6535 ( 
.A(n_5922),
.Y(n_6535)
);

BUFx2_ASAP7_75t_L g6536 ( 
.A(n_5922),
.Y(n_6536)
);

BUFx8_ASAP7_75t_L g6537 ( 
.A(n_5947),
.Y(n_6537)
);

BUFx6f_ASAP7_75t_L g6538 ( 
.A(n_5609),
.Y(n_6538)
);

BUFx6f_ASAP7_75t_L g6539 ( 
.A(n_5609),
.Y(n_6539)
);

AND2x4_ASAP7_75t_L g6540 ( 
.A(n_5955),
.B(n_3998),
.Y(n_6540)
);

BUFx6f_ASAP7_75t_L g6541 ( 
.A(n_5609),
.Y(n_6541)
);

BUFx3_ASAP7_75t_L g6542 ( 
.A(n_5955),
.Y(n_6542)
);

OAI21x1_ASAP7_75t_L g6543 ( 
.A1(n_5883),
.A2(n_4593),
.B(n_4588),
.Y(n_6543)
);

AND2x2_ASAP7_75t_SL g6544 ( 
.A(n_5848),
.B(n_4601),
.Y(n_6544)
);

AND2x2_ASAP7_75t_SL g6545 ( 
.A(n_5848),
.B(n_4623),
.Y(n_6545)
);

OAI22xp5_ASAP7_75t_L g6546 ( 
.A1(n_5645),
.A2(n_3766),
.B1(n_3773),
.B2(n_3765),
.Y(n_6546)
);

AND2x4_ASAP7_75t_L g6547 ( 
.A(n_5955),
.B(n_4002),
.Y(n_6547)
);

OAI22xp5_ASAP7_75t_L g6548 ( 
.A1(n_5645),
.A2(n_3775),
.B1(n_3776),
.B2(n_3774),
.Y(n_6548)
);

AND2x4_ASAP7_75t_L g6549 ( 
.A(n_5955),
.B(n_4003),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_5760),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_5686),
.B(n_4474),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_5877),
.B(n_4648),
.Y(n_6552)
);

NOR2xp33_ASAP7_75t_L g6553 ( 
.A(n_5528),
.B(n_3777),
.Y(n_6553)
);

INVxp67_ASAP7_75t_L g6554 ( 
.A(n_5922),
.Y(n_6554)
);

NAND2xp5_ASAP7_75t_SL g6555 ( 
.A(n_5922),
.B(n_3778),
.Y(n_6555)
);

AOI22xp5_ASAP7_75t_L g6556 ( 
.A1(n_5645),
.A2(n_3781),
.B1(n_3782),
.B2(n_3779),
.Y(n_6556)
);

BUFx6f_ASAP7_75t_L g6557 ( 
.A(n_5609),
.Y(n_6557)
);

BUFx6f_ASAP7_75t_L g6558 ( 
.A(n_5609),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_5686),
.B(n_4474),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_5492),
.Y(n_6560)
);

OAI21x1_ASAP7_75t_L g6561 ( 
.A1(n_5883),
.A2(n_4685),
.B(n_4660),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_5760),
.Y(n_6562)
);

OAI22xp5_ASAP7_75t_L g6563 ( 
.A1(n_5645),
.A2(n_3785),
.B1(n_3786),
.B2(n_3784),
.Y(n_6563)
);

NAND2xp5_ASAP7_75t_L g6564 ( 
.A(n_5877),
.B(n_4699),
.Y(n_6564)
);

BUFx6f_ASAP7_75t_L g6565 ( 
.A(n_5609),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_5760),
.Y(n_6566)
);

BUFx6f_ASAP7_75t_L g6567 ( 
.A(n_5609),
.Y(n_6567)
);

INVx1_ASAP7_75t_L g6568 ( 
.A(n_6566),
.Y(n_6568)
);

NAND2xp5_ASAP7_75t_L g6569 ( 
.A(n_6042),
.B(n_3787),
.Y(n_6569)
);

BUFx6f_ASAP7_75t_L g6570 ( 
.A(n_5993),
.Y(n_6570)
);

NAND2xp5_ASAP7_75t_L g6571 ( 
.A(n_6293),
.B(n_3789),
.Y(n_6571)
);

XNOR2xp5_ASAP7_75t_L g6572 ( 
.A(n_6492),
.B(n_4709),
.Y(n_6572)
);

INVxp67_ASAP7_75t_L g6573 ( 
.A(n_6056),
.Y(n_6573)
);

AND2x6_ASAP7_75t_L g6574 ( 
.A(n_6437),
.B(n_4016),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6562),
.Y(n_6575)
);

NOR2xp33_ASAP7_75t_L g6576 ( 
.A(n_6068),
.B(n_3790),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_5995),
.Y(n_6577)
);

NAND2xp5_ASAP7_75t_L g6578 ( 
.A(n_6111),
.B(n_3791),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5996),
.Y(n_6579)
);

INVx2_ASAP7_75t_L g6580 ( 
.A(n_6009),
.Y(n_6580)
);

BUFx6f_ASAP7_75t_L g6581 ( 
.A(n_5994),
.Y(n_6581)
);

CKINVDCx5p33_ASAP7_75t_R g6582 ( 
.A(n_6188),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6001),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6215),
.B(n_3792),
.Y(n_6584)
);

INVx3_ASAP7_75t_L g6585 ( 
.A(n_6085),
.Y(n_6585)
);

CKINVDCx5p33_ASAP7_75t_R g6586 ( 
.A(n_6064),
.Y(n_6586)
);

OAI22xp5_ASAP7_75t_SL g6587 ( 
.A1(n_6460),
.A2(n_4758),
.B1(n_4764),
.B2(n_4734),
.Y(n_6587)
);

INVx2_ASAP7_75t_L g6588 ( 
.A(n_6010),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6006),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6011),
.Y(n_6590)
);

HB1xp67_ASAP7_75t_L g6591 ( 
.A(n_6063),
.Y(n_6591)
);

BUFx6f_ASAP7_75t_L g6592 ( 
.A(n_5998),
.Y(n_6592)
);

INVx3_ASAP7_75t_L g6593 ( 
.A(n_6087),
.Y(n_6593)
);

BUFx2_ASAP7_75t_L g6594 ( 
.A(n_6076),
.Y(n_6594)
);

BUFx6f_ASAP7_75t_L g6595 ( 
.A(n_6501),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_6075),
.Y(n_6596)
);

INVx2_ASAP7_75t_L g6597 ( 
.A(n_6080),
.Y(n_6597)
);

AND2x2_ASAP7_75t_SL g6598 ( 
.A(n_6468),
.B(n_4715),
.Y(n_6598)
);

CKINVDCx5p33_ASAP7_75t_R g6599 ( 
.A(n_6114),
.Y(n_6599)
);

BUFx2_ASAP7_75t_L g6600 ( 
.A(n_6095),
.Y(n_6600)
);

XNOR2xp5_ASAP7_75t_L g6601 ( 
.A(n_6178),
.B(n_4776),
.Y(n_6601)
);

INVx2_ASAP7_75t_L g6602 ( 
.A(n_5988),
.Y(n_6602)
);

CKINVDCx5p33_ASAP7_75t_R g6603 ( 
.A(n_6123),
.Y(n_6603)
);

INVx3_ASAP7_75t_L g6604 ( 
.A(n_6094),
.Y(n_6604)
);

CKINVDCx5p33_ASAP7_75t_R g6605 ( 
.A(n_6129),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6007),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_6017),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6018),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6020),
.Y(n_6609)
);

INVx2_ASAP7_75t_L g6610 ( 
.A(n_5997),
.Y(n_6610)
);

NOR2xp33_ASAP7_75t_L g6611 ( 
.A(n_6165),
.B(n_3797),
.Y(n_6611)
);

AND2x4_ASAP7_75t_L g6612 ( 
.A(n_5989),
.B(n_4018),
.Y(n_6612)
);

CKINVDCx14_ASAP7_75t_R g6613 ( 
.A(n_6012),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6024),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6035),
.Y(n_6615)
);

INVx2_ASAP7_75t_L g6616 ( 
.A(n_5999),
.Y(n_6616)
);

AND2x4_ASAP7_75t_L g6617 ( 
.A(n_6518),
.B(n_4020),
.Y(n_6617)
);

BUFx3_ASAP7_75t_L g6618 ( 
.A(n_6039),
.Y(n_6618)
);

CKINVDCx5p33_ASAP7_75t_R g6619 ( 
.A(n_6166),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6223),
.B(n_3799),
.Y(n_6620)
);

CKINVDCx20_ASAP7_75t_R g6621 ( 
.A(n_6379),
.Y(n_6621)
);

CKINVDCx5p33_ASAP7_75t_R g6622 ( 
.A(n_6211),
.Y(n_6622)
);

CKINVDCx5p33_ASAP7_75t_R g6623 ( 
.A(n_6221),
.Y(n_6623)
);

CKINVDCx5p33_ASAP7_75t_R g6624 ( 
.A(n_6222),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6041),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_6044),
.Y(n_6626)
);

CKINVDCx5p33_ASAP7_75t_R g6627 ( 
.A(n_6315),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6045),
.Y(n_6628)
);

CKINVDCx20_ASAP7_75t_R g6629 ( 
.A(n_6419),
.Y(n_6629)
);

CKINVDCx5p33_ASAP7_75t_R g6630 ( 
.A(n_6414),
.Y(n_6630)
);

AND2x2_ASAP7_75t_SL g6631 ( 
.A(n_6033),
.B(n_4803),
.Y(n_6631)
);

CKINVDCx5p33_ASAP7_75t_R g6632 ( 
.A(n_6508),
.Y(n_6632)
);

HB1xp67_ASAP7_75t_L g6633 ( 
.A(n_6393),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6047),
.Y(n_6634)
);

CKINVDCx20_ASAP7_75t_R g6635 ( 
.A(n_6483),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6050),
.Y(n_6636)
);

INVx2_ASAP7_75t_L g6637 ( 
.A(n_6002),
.Y(n_6637)
);

CKINVDCx5p33_ASAP7_75t_R g6638 ( 
.A(n_6511),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6058),
.Y(n_6639)
);

NAND2xp5_ASAP7_75t_SL g6640 ( 
.A(n_6499),
.B(n_3800),
.Y(n_6640)
);

CKINVDCx20_ASAP7_75t_R g6641 ( 
.A(n_6316),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6507),
.Y(n_6642)
);

BUFx6f_ASAP7_75t_L g6643 ( 
.A(n_6506),
.Y(n_6643)
);

CKINVDCx20_ASAP7_75t_R g6644 ( 
.A(n_6382),
.Y(n_6644)
);

NAND2xp33_ASAP7_75t_L g6645 ( 
.A(n_6526),
.B(n_3803),
.Y(n_6645)
);

INVx3_ASAP7_75t_L g6646 ( 
.A(n_6520),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6513),
.Y(n_6647)
);

AND2x2_ASAP7_75t_L g6648 ( 
.A(n_6535),
.B(n_4484),
.Y(n_6648)
);

CKINVDCx5p33_ASAP7_75t_R g6649 ( 
.A(n_6514),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6530),
.Y(n_6650)
);

CKINVDCx20_ASAP7_75t_R g6651 ( 
.A(n_6140),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6066),
.Y(n_6652)
);

NOR2xp33_ASAP7_75t_L g6653 ( 
.A(n_6432),
.B(n_3804),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6070),
.Y(n_6654)
);

CKINVDCx5p33_ASAP7_75t_R g6655 ( 
.A(n_6206),
.Y(n_6655)
);

INVx2_ASAP7_75t_L g6656 ( 
.A(n_6533),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6560),
.Y(n_6657)
);

NOR3xp33_ASAP7_75t_L g6658 ( 
.A(n_6077),
.B(n_3811),
.C(n_3808),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_6088),
.Y(n_6659)
);

XNOR2xp5_ASAP7_75t_L g6660 ( 
.A(n_6273),
.B(n_4780),
.Y(n_6660)
);

CKINVDCx5p33_ASAP7_75t_R g6661 ( 
.A(n_6233),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6072),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6078),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6079),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_6096),
.Y(n_6665)
);

INVx1_ASAP7_75t_L g6666 ( 
.A(n_6081),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6101),
.Y(n_6667)
);

CKINVDCx8_ASAP7_75t_R g6668 ( 
.A(n_6000),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6086),
.Y(n_6669)
);

BUFx2_ASAP7_75t_L g6670 ( 
.A(n_6404),
.Y(n_6670)
);

CKINVDCx5p33_ASAP7_75t_R g6671 ( 
.A(n_6282),
.Y(n_6671)
);

INVx3_ASAP7_75t_L g6672 ( 
.A(n_6522),
.Y(n_6672)
);

NAND2xp33_ASAP7_75t_L g6673 ( 
.A(n_6526),
.B(n_3813),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6536),
.B(n_4484),
.Y(n_6674)
);

CKINVDCx5p33_ASAP7_75t_R g6675 ( 
.A(n_6290),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6089),
.Y(n_6676)
);

INVx2_ASAP7_75t_L g6677 ( 
.A(n_6106),
.Y(n_6677)
);

NAND2xp5_ASAP7_75t_L g6678 ( 
.A(n_6236),
.B(n_3820),
.Y(n_6678)
);

INVx2_ASAP7_75t_L g6679 ( 
.A(n_6403),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_5990),
.B(n_4528),
.Y(n_6680)
);

INVx2_ASAP7_75t_L g6681 ( 
.A(n_6411),
.Y(n_6681)
);

CKINVDCx5p33_ASAP7_75t_R g6682 ( 
.A(n_6377),
.Y(n_6682)
);

CKINVDCx5p33_ASAP7_75t_R g6683 ( 
.A(n_6385),
.Y(n_6683)
);

NAND2xp5_ASAP7_75t_L g6684 ( 
.A(n_6240),
.B(n_3822),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_6424),
.Y(n_6685)
);

CKINVDCx20_ASAP7_75t_R g6686 ( 
.A(n_6201),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6241),
.B(n_3824),
.Y(n_6687)
);

HB1xp67_ASAP7_75t_L g6688 ( 
.A(n_6503),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6090),
.Y(n_6689)
);

NAND2xp5_ASAP7_75t_L g6690 ( 
.A(n_6251),
.B(n_3828),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6098),
.Y(n_6691)
);

AND2x2_ASAP7_75t_L g6692 ( 
.A(n_6109),
.B(n_4528),
.Y(n_6692)
);

INVx2_ASAP7_75t_L g6693 ( 
.A(n_6116),
.Y(n_6693)
);

INVx2_ASAP7_75t_L g6694 ( 
.A(n_6117),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6102),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_L g6696 ( 
.A(n_6253),
.B(n_3831),
.Y(n_6696)
);

CKINVDCx5p33_ASAP7_75t_R g6697 ( 
.A(n_6391),
.Y(n_6697)
);

CKINVDCx5p33_ASAP7_75t_R g6698 ( 
.A(n_6416),
.Y(n_6698)
);

BUFx6f_ASAP7_75t_L g6699 ( 
.A(n_6523),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6122),
.Y(n_6700)
);

NAND2xp5_ASAP7_75t_L g6701 ( 
.A(n_6256),
.B(n_6265),
.Y(n_6701)
);

CKINVDCx20_ASAP7_75t_R g6702 ( 
.A(n_6027),
.Y(n_6702)
);

AND2x4_ASAP7_75t_L g6703 ( 
.A(n_6542),
.B(n_4024),
.Y(n_6703)
);

CKINVDCx5p33_ASAP7_75t_R g6704 ( 
.A(n_6447),
.Y(n_6704)
);

CKINVDCx5p33_ASAP7_75t_R g6705 ( 
.A(n_6502),
.Y(n_6705)
);

BUFx6f_ASAP7_75t_L g6706 ( 
.A(n_6538),
.Y(n_6706)
);

CKINVDCx5p33_ASAP7_75t_R g6707 ( 
.A(n_6509),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6126),
.Y(n_6708)
);

CKINVDCx20_ASAP7_75t_R g6709 ( 
.A(n_6203),
.Y(n_6709)
);

AND2x2_ASAP7_75t_L g6710 ( 
.A(n_6127),
.B(n_4539),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_6128),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6145),
.Y(n_6712)
);

INVx1_ASAP7_75t_L g6713 ( 
.A(n_6156),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6158),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6160),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6168),
.Y(n_6716)
);

INVx2_ASAP7_75t_L g6717 ( 
.A(n_6118),
.Y(n_6717)
);

NAND2xp5_ASAP7_75t_L g6718 ( 
.A(n_6052),
.B(n_3833),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6175),
.Y(n_6719)
);

NAND2xp5_ASAP7_75t_SL g6720 ( 
.A(n_6327),
.B(n_6333),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6179),
.Y(n_6721)
);

CKINVDCx5p33_ASAP7_75t_R g6722 ( 
.A(n_6433),
.Y(n_6722)
);

INVx3_ASAP7_75t_L g6723 ( 
.A(n_6539),
.Y(n_6723)
);

OA21x2_ASAP7_75t_L g6724 ( 
.A1(n_6112),
.A2(n_4035),
.B(n_4025),
.Y(n_6724)
);

CKINVDCx5p33_ASAP7_75t_R g6725 ( 
.A(n_6434),
.Y(n_6725)
);

INVx2_ASAP7_75t_L g6726 ( 
.A(n_6125),
.Y(n_6726)
);

HB1xp67_ASAP7_75t_L g6727 ( 
.A(n_6551),
.Y(n_6727)
);

NAND2x1p5_ASAP7_75t_L g6728 ( 
.A(n_6040),
.B(n_4036),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6182),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6183),
.Y(n_6730)
);

INVx2_ASAP7_75t_L g6731 ( 
.A(n_6132),
.Y(n_6731)
);

BUFx6f_ASAP7_75t_L g6732 ( 
.A(n_6541),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6185),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_6133),
.Y(n_6734)
);

CKINVDCx5p33_ASAP7_75t_R g6735 ( 
.A(n_6436),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6554),
.B(n_4539),
.Y(n_6736)
);

CKINVDCx5p33_ASAP7_75t_R g6737 ( 
.A(n_6449),
.Y(n_6737)
);

INVx3_ASAP7_75t_L g6738 ( 
.A(n_6557),
.Y(n_6738)
);

BUFx3_ASAP7_75t_L g6739 ( 
.A(n_6055),
.Y(n_6739)
);

AND2x2_ASAP7_75t_L g6740 ( 
.A(n_6559),
.B(n_4612),
.Y(n_6740)
);

CKINVDCx5p33_ASAP7_75t_R g6741 ( 
.A(n_6450),
.Y(n_6741)
);

AOI22xp5_ASAP7_75t_L g6742 ( 
.A1(n_6398),
.A2(n_6157),
.B1(n_6553),
.B2(n_6003),
.Y(n_6742)
);

INVx2_ASAP7_75t_L g6743 ( 
.A(n_6135),
.Y(n_6743)
);

CKINVDCx5p33_ASAP7_75t_R g6744 ( 
.A(n_6473),
.Y(n_6744)
);

AOI22xp5_ASAP7_75t_L g6745 ( 
.A1(n_5991),
.A2(n_4839),
.B1(n_4848),
.B2(n_4823),
.Y(n_6745)
);

AND2x2_ASAP7_75t_R g6746 ( 
.A(n_6372),
.B(n_4037),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_6194),
.Y(n_6747)
);

NOR2xp33_ASAP7_75t_R g6748 ( 
.A(n_6061),
.B(n_4860),
.Y(n_6748)
);

INVx2_ASAP7_75t_L g6749 ( 
.A(n_6159),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6494),
.Y(n_6750)
);

CKINVDCx5p33_ASAP7_75t_R g6751 ( 
.A(n_6373),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_6495),
.Y(n_6752)
);

OA21x2_ASAP7_75t_L g6753 ( 
.A1(n_6154),
.A2(n_4050),
.B(n_4042),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6161),
.Y(n_6754)
);

AND2x4_ASAP7_75t_L g6755 ( 
.A(n_6519),
.B(n_4051),
.Y(n_6755)
);

INVx1_ASAP7_75t_L g6756 ( 
.A(n_6496),
.Y(n_6756)
);

INVx2_ASAP7_75t_L g6757 ( 
.A(n_6163),
.Y(n_6757)
);

NOR2xp67_ASAP7_75t_L g6758 ( 
.A(n_6062),
.B(n_3378),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_6498),
.Y(n_6759)
);

NOR2xp33_ASAP7_75t_R g6760 ( 
.A(n_6065),
.B(n_4871),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6504),
.Y(n_6761)
);

CKINVDCx5p33_ASAP7_75t_R g6762 ( 
.A(n_6374),
.Y(n_6762)
);

CKINVDCx5p33_ASAP7_75t_R g6763 ( 
.A(n_6378),
.Y(n_6763)
);

CKINVDCx5p33_ASAP7_75t_R g6764 ( 
.A(n_6420),
.Y(n_6764)
);

CKINVDCx5p33_ASAP7_75t_R g6765 ( 
.A(n_6148),
.Y(n_6765)
);

NAND2xp5_ASAP7_75t_L g6766 ( 
.A(n_6500),
.B(n_3834),
.Y(n_6766)
);

INVx1_ASAP7_75t_L g6767 ( 
.A(n_6515),
.Y(n_6767)
);

NOR2xp33_ASAP7_75t_R g6768 ( 
.A(n_6099),
.B(n_4880),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6516),
.Y(n_6769)
);

INVx2_ASAP7_75t_L g6770 ( 
.A(n_6167),
.Y(n_6770)
);

INVx3_ASAP7_75t_L g6771 ( 
.A(n_6558),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6525),
.Y(n_6772)
);

INVx2_ASAP7_75t_L g6773 ( 
.A(n_6171),
.Y(n_6773)
);

HB1xp67_ASAP7_75t_L g6774 ( 
.A(n_6054),
.Y(n_6774)
);

BUFx2_ASAP7_75t_L g6775 ( 
.A(n_6131),
.Y(n_6775)
);

CKINVDCx20_ASAP7_75t_R g6776 ( 
.A(n_6193),
.Y(n_6776)
);

CKINVDCx5p33_ASAP7_75t_R g6777 ( 
.A(n_6184),
.Y(n_6777)
);

BUFx6f_ASAP7_75t_L g6778 ( 
.A(n_6565),
.Y(n_6778)
);

INVx2_ASAP7_75t_L g6779 ( 
.A(n_6173),
.Y(n_6779)
);

CKINVDCx5p33_ASAP7_75t_R g6780 ( 
.A(n_6249),
.Y(n_6780)
);

INVx2_ASAP7_75t_L g6781 ( 
.A(n_6176),
.Y(n_6781)
);

CKINVDCx5p33_ASAP7_75t_R g6782 ( 
.A(n_6396),
.Y(n_6782)
);

BUFx2_ASAP7_75t_L g6783 ( 
.A(n_6147),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6529),
.Y(n_6784)
);

CKINVDCx5p33_ASAP7_75t_R g6785 ( 
.A(n_6401),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6550),
.Y(n_6786)
);

CKINVDCx20_ASAP7_75t_R g6787 ( 
.A(n_6415),
.Y(n_6787)
);

CKINVDCx20_ASAP7_75t_R g6788 ( 
.A(n_6476),
.Y(n_6788)
);

CKINVDCx5p33_ASAP7_75t_R g6789 ( 
.A(n_6487),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_SL g6790 ( 
.A(n_6451),
.B(n_3836),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6301),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6150),
.B(n_4612),
.Y(n_6792)
);

BUFx6f_ASAP7_75t_L g6793 ( 
.A(n_6567),
.Y(n_6793)
);

CKINVDCx5p33_ASAP7_75t_R g6794 ( 
.A(n_6491),
.Y(n_6794)
);

CKINVDCx5p33_ASAP7_75t_R g6795 ( 
.A(n_6324),
.Y(n_6795)
);

CKINVDCx5p33_ASAP7_75t_R g6796 ( 
.A(n_6104),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_6320),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6337),
.Y(n_6798)
);

CKINVDCx20_ASAP7_75t_R g6799 ( 
.A(n_6013),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6343),
.Y(n_6800)
);

CKINVDCx20_ASAP7_75t_R g6801 ( 
.A(n_6021),
.Y(n_6801)
);

CKINVDCx16_ASAP7_75t_R g6802 ( 
.A(n_6069),
.Y(n_6802)
);

BUFx12f_ASAP7_75t_L g6803 ( 
.A(n_6120),
.Y(n_6803)
);

CKINVDCx20_ASAP7_75t_R g6804 ( 
.A(n_6537),
.Y(n_6804)
);

CKINVDCx5p33_ASAP7_75t_R g6805 ( 
.A(n_6107),
.Y(n_6805)
);

CKINVDCx16_ASAP7_75t_R g6806 ( 
.A(n_6196),
.Y(n_6806)
);

INVx3_ASAP7_75t_L g6807 ( 
.A(n_6005),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6361),
.Y(n_6808)
);

NAND2xp5_ASAP7_75t_L g6809 ( 
.A(n_6552),
.B(n_3837),
.Y(n_6809)
);

INVx2_ASAP7_75t_L g6810 ( 
.A(n_6181),
.Y(n_6810)
);

INVx1_ASAP7_75t_L g6811 ( 
.A(n_6367),
.Y(n_6811)
);

CKINVDCx5p33_ASAP7_75t_R g6812 ( 
.A(n_6172),
.Y(n_6812)
);

CKINVDCx5p33_ASAP7_75t_R g6813 ( 
.A(n_6235),
.Y(n_6813)
);

AND2x4_ASAP7_75t_L g6814 ( 
.A(n_6524),
.B(n_4054),
.Y(n_6814)
);

NAND2xp5_ASAP7_75t_SL g6815 ( 
.A(n_6453),
.B(n_3841),
.Y(n_6815)
);

NOR2xp33_ASAP7_75t_R g6816 ( 
.A(n_6108),
.B(n_4890),
.Y(n_6816)
);

INVx2_ASAP7_75t_L g6817 ( 
.A(n_6187),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6375),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6390),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6399),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6400),
.Y(n_6821)
);

INVx1_ASAP7_75t_L g6822 ( 
.A(n_6409),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6271),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6192),
.Y(n_6824)
);

INVx3_ASAP7_75t_L g6825 ( 
.A(n_6008),
.Y(n_6825)
);

CKINVDCx5p33_ASAP7_75t_R g6826 ( 
.A(n_6323),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6198),
.Y(n_6827)
);

CKINVDCx5p33_ASAP7_75t_R g6828 ( 
.A(n_6394),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6277),
.Y(n_6829)
);

AND2x4_ASAP7_75t_L g6830 ( 
.A(n_6534),
.B(n_4055),
.Y(n_6830)
);

CKINVDCx5p33_ASAP7_75t_R g6831 ( 
.A(n_6445),
.Y(n_6831)
);

CKINVDCx5p33_ASAP7_75t_R g6832 ( 
.A(n_6512),
.Y(n_6832)
);

CKINVDCx5p33_ASAP7_75t_R g6833 ( 
.A(n_6478),
.Y(n_6833)
);

CKINVDCx5p33_ASAP7_75t_R g6834 ( 
.A(n_6191),
.Y(n_6834)
);

INVx2_ASAP7_75t_L g6835 ( 
.A(n_6199),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_6564),
.B(n_6110),
.Y(n_6836)
);

NAND3xp33_ASAP7_75t_L g6837 ( 
.A(n_6527),
.B(n_6556),
.C(n_6263),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6280),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6284),
.Y(n_6839)
);

CKINVDCx5p33_ASAP7_75t_R g6840 ( 
.A(n_6180),
.Y(n_6840)
);

BUFx6f_ASAP7_75t_L g6841 ( 
.A(n_6014),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_6299),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_6202),
.Y(n_6843)
);

AND2x2_ASAP7_75t_L g6844 ( 
.A(n_6197),
.B(n_4724),
.Y(n_6844)
);

NOR2xp33_ASAP7_75t_L g6845 ( 
.A(n_6462),
.B(n_6312),
.Y(n_6845)
);

NAND2xp5_ASAP7_75t_L g6846 ( 
.A(n_6124),
.B(n_6121),
.Y(n_6846)
);

INVx3_ASAP7_75t_L g6847 ( 
.A(n_6026),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6300),
.Y(n_6848)
);

NAND2xp5_ASAP7_75t_L g6849 ( 
.A(n_6267),
.B(n_6479),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_6410),
.Y(n_6850)
);

AND2x4_ASAP7_75t_L g6851 ( 
.A(n_6497),
.B(n_6517),
.Y(n_6851)
);

INVx6_ASAP7_75t_L g6852 ( 
.A(n_6234),
.Y(n_6852)
);

AND2x2_ASAP7_75t_L g6853 ( 
.A(n_6368),
.B(n_4724),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6421),
.Y(n_6854)
);

CKINVDCx5p33_ASAP7_75t_R g6855 ( 
.A(n_6458),
.Y(n_6855)
);

HB1xp67_ASAP7_75t_L g6856 ( 
.A(n_6490),
.Y(n_6856)
);

CKINVDCx5p33_ASAP7_75t_R g6857 ( 
.A(n_6356),
.Y(n_6857)
);

INVx5_ASAP7_75t_L g6858 ( 
.A(n_6349),
.Y(n_6858)
);

CKINVDCx5p33_ASAP7_75t_R g6859 ( 
.A(n_6369),
.Y(n_6859)
);

BUFx6f_ASAP7_75t_L g6860 ( 
.A(n_6029),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6423),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6482),
.B(n_3845),
.Y(n_6862)
);

BUFx6f_ASAP7_75t_L g6863 ( 
.A(n_6031),
.Y(n_6863)
);

CKINVDCx5p33_ASAP7_75t_R g6864 ( 
.A(n_6392),
.Y(n_6864)
);

INVx3_ASAP7_75t_L g6865 ( 
.A(n_6100),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6428),
.Y(n_6866)
);

CKINVDCx5p33_ASAP7_75t_R g6867 ( 
.A(n_6435),
.Y(n_6867)
);

INVx2_ASAP7_75t_L g6868 ( 
.A(n_6212),
.Y(n_6868)
);

CKINVDCx16_ASAP7_75t_R g6869 ( 
.A(n_6250),
.Y(n_6869)
);

INVx2_ASAP7_75t_L g6870 ( 
.A(n_6216),
.Y(n_6870)
);

BUFx3_ASAP7_75t_L g6871 ( 
.A(n_6247),
.Y(n_6871)
);

INVx3_ASAP7_75t_L g6872 ( 
.A(n_6113),
.Y(n_6872)
);

AND2x2_ASAP7_75t_L g6873 ( 
.A(n_6093),
.B(n_4784),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6406),
.Y(n_6874)
);

BUFx2_ASAP7_75t_L g6875 ( 
.A(n_6105),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6544),
.B(n_4784),
.Y(n_6876)
);

INVx1_ASAP7_75t_SL g6877 ( 
.A(n_6204),
.Y(n_6877)
);

INVx2_ASAP7_75t_L g6878 ( 
.A(n_6218),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6226),
.Y(n_6879)
);

AND2x2_ASAP7_75t_L g6880 ( 
.A(n_6545),
.B(n_4806),
.Y(n_6880)
);

INVx2_ASAP7_75t_L g6881 ( 
.A(n_6227),
.Y(n_6881)
);

CKINVDCx5p33_ASAP7_75t_R g6882 ( 
.A(n_6439),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6242),
.Y(n_6883)
);

INVx3_ASAP7_75t_L g6884 ( 
.A(n_6136),
.Y(n_6884)
);

INVxp33_ASAP7_75t_L g6885 ( 
.A(n_6092),
.Y(n_6885)
);

INVx2_ASAP7_75t_L g6886 ( 
.A(n_6243),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6248),
.Y(n_6887)
);

CKINVDCx5p33_ASAP7_75t_R g6888 ( 
.A(n_6229),
.Y(n_6888)
);

INVx1_ASAP7_75t_L g6889 ( 
.A(n_6252),
.Y(n_6889)
);

NAND2xp5_ASAP7_75t_SL g6890 ( 
.A(n_6016),
.B(n_3847),
.Y(n_6890)
);

NOR2xp33_ASAP7_75t_L g6891 ( 
.A(n_6351),
.B(n_3848),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6259),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6260),
.Y(n_6893)
);

CKINVDCx5p33_ASAP7_75t_R g6894 ( 
.A(n_6340),
.Y(n_6894)
);

AND2x4_ASAP7_75t_L g6895 ( 
.A(n_6531),
.B(n_4064),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_6261),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_6103),
.B(n_3849),
.Y(n_6897)
);

BUFx3_ASAP7_75t_L g6898 ( 
.A(n_6311),
.Y(n_6898)
);

CKINVDCx5p33_ASAP7_75t_R g6899 ( 
.A(n_6454),
.Y(n_6899)
);

NAND2xp33_ASAP7_75t_L g6900 ( 
.A(n_6208),
.B(n_3851),
.Y(n_6900)
);

INVx2_ASAP7_75t_L g6901 ( 
.A(n_6285),
.Y(n_6901)
);

NAND2xp5_ASAP7_75t_SL g6902 ( 
.A(n_6474),
.B(n_3853),
.Y(n_6902)
);

BUFx2_ASAP7_75t_L g6903 ( 
.A(n_6091),
.Y(n_6903)
);

INVx3_ASAP7_75t_L g6904 ( 
.A(n_6138),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6294),
.Y(n_6905)
);

BUFx6f_ASAP7_75t_L g6906 ( 
.A(n_6043),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6295),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6298),
.Y(n_6908)
);

CKINVDCx5p33_ASAP7_75t_R g6909 ( 
.A(n_6220),
.Y(n_6909)
);

CKINVDCx5p33_ASAP7_75t_R g6910 ( 
.A(n_6228),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6307),
.Y(n_6911)
);

AND2x4_ASAP7_75t_L g6912 ( 
.A(n_6532),
.B(n_4069),
.Y(n_6912)
);

CKINVDCx5p33_ASAP7_75t_R g6913 ( 
.A(n_6275),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6305),
.B(n_3857),
.Y(n_6914)
);

CKINVDCx5p33_ASAP7_75t_R g6915 ( 
.A(n_6304),
.Y(n_6915)
);

NOR2xp33_ASAP7_75t_L g6916 ( 
.A(n_6376),
.B(n_3861),
.Y(n_6916)
);

NAND2xp5_ASAP7_75t_L g6917 ( 
.A(n_6015),
.B(n_6019),
.Y(n_6917)
);

INVx3_ASAP7_75t_L g6918 ( 
.A(n_6143),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_6308),
.Y(n_6919)
);

INVx2_ASAP7_75t_L g6920 ( 
.A(n_6317),
.Y(n_6920)
);

CKINVDCx5p33_ASAP7_75t_R g6921 ( 
.A(n_6292),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6318),
.Y(n_6922)
);

BUFx6f_ASAP7_75t_L g6923 ( 
.A(n_6048),
.Y(n_6923)
);

CKINVDCx5p33_ASAP7_75t_R g6924 ( 
.A(n_6440),
.Y(n_6924)
);

BUFx8_ASAP7_75t_L g6925 ( 
.A(n_6481),
.Y(n_6925)
);

BUFx6f_ASAP7_75t_L g6926 ( 
.A(n_6144),
.Y(n_6926)
);

BUFx3_ASAP7_75t_L g6927 ( 
.A(n_6540),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_L g6928 ( 
.A(n_6030),
.B(n_3862),
.Y(n_6928)
);

CKINVDCx5p33_ASAP7_75t_R g6929 ( 
.A(n_6443),
.Y(n_6929)
);

HB1xp67_ASAP7_75t_L g6930 ( 
.A(n_6457),
.Y(n_6930)
);

CKINVDCx5p33_ASAP7_75t_R g6931 ( 
.A(n_6448),
.Y(n_6931)
);

BUFx3_ASAP7_75t_L g6932 ( 
.A(n_6547),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6319),
.Y(n_6933)
);

INVx2_ASAP7_75t_L g6934 ( 
.A(n_6321),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_6034),
.B(n_3868),
.Y(n_6935)
);

INVx3_ASAP7_75t_L g6936 ( 
.A(n_6151),
.Y(n_6936)
);

INVx6_ASAP7_75t_L g6937 ( 
.A(n_6322),
.Y(n_6937)
);

CKINVDCx5p33_ASAP7_75t_R g6938 ( 
.A(n_6456),
.Y(n_6938)
);

NAND2xp5_ASAP7_75t_L g6939 ( 
.A(n_6038),
.B(n_3869),
.Y(n_6939)
);

CKINVDCx5p33_ASAP7_75t_R g6940 ( 
.A(n_6464),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6325),
.Y(n_6941)
);

BUFx2_ASAP7_75t_L g6942 ( 
.A(n_6091),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6328),
.Y(n_6943)
);

BUFx6f_ASAP7_75t_L g6944 ( 
.A(n_6195),
.Y(n_6944)
);

AND2x4_ASAP7_75t_L g6945 ( 
.A(n_6549),
.B(n_4072),
.Y(n_6945)
);

CKINVDCx5p33_ASAP7_75t_R g6946 ( 
.A(n_6465),
.Y(n_6946)
);

CKINVDCx20_ASAP7_75t_R g6947 ( 
.A(n_6232),
.Y(n_6947)
);

INVx3_ASAP7_75t_L g6948 ( 
.A(n_6209),
.Y(n_6948)
);

CKINVDCx20_ASAP7_75t_R g6949 ( 
.A(n_6417),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6332),
.Y(n_6950)
);

INVx2_ASAP7_75t_L g6951 ( 
.A(n_6338),
.Y(n_6951)
);

BUFx6f_ASAP7_75t_L g6952 ( 
.A(n_6210),
.Y(n_6952)
);

AOI22xp5_ASAP7_75t_L g6953 ( 
.A1(n_6238),
.A2(n_4895),
.B1(n_4904),
.B2(n_4892),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6344),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6350),
.Y(n_6955)
);

CKINVDCx5p33_ASAP7_75t_R g6956 ( 
.A(n_6266),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6046),
.B(n_3872),
.Y(n_6957)
);

CKINVDCx5p33_ASAP7_75t_R g6958 ( 
.A(n_6455),
.Y(n_6958)
);

INVx3_ASAP7_75t_L g6959 ( 
.A(n_6213),
.Y(n_6959)
);

BUFx6f_ASAP7_75t_L g6960 ( 
.A(n_6237),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6354),
.Y(n_6961)
);

NAND2xp5_ASAP7_75t_L g6962 ( 
.A(n_6053),
.B(n_3873),
.Y(n_6962)
);

HB1xp67_ASAP7_75t_L g6963 ( 
.A(n_6219),
.Y(n_6963)
);

HB1xp67_ASAP7_75t_L g6964 ( 
.A(n_6245),
.Y(n_6964)
);

BUFx6f_ASAP7_75t_L g6965 ( 
.A(n_6244),
.Y(n_6965)
);

BUFx2_ASAP7_75t_L g6966 ( 
.A(n_6349),
.Y(n_6966)
);

AND2x2_ASAP7_75t_L g6967 ( 
.A(n_6466),
.B(n_4806),
.Y(n_6967)
);

INVx2_ASAP7_75t_L g6968 ( 
.A(n_6357),
.Y(n_6968)
);

INVx2_ASAP7_75t_L g6969 ( 
.A(n_6366),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6380),
.Y(n_6970)
);

NAND2xp5_ASAP7_75t_L g6971 ( 
.A(n_6060),
.B(n_3874),
.Y(n_6971)
);

CKINVDCx5p33_ASAP7_75t_R g6972 ( 
.A(n_6459),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6383),
.Y(n_6973)
);

AND2x4_ASAP7_75t_L g6974 ( 
.A(n_6334),
.B(n_4077),
.Y(n_6974)
);

INVx2_ASAP7_75t_L g6975 ( 
.A(n_6387),
.Y(n_6975)
);

BUFx8_ASAP7_75t_L g6976 ( 
.A(n_6485),
.Y(n_6976)
);

NOR2xp33_ASAP7_75t_R g6977 ( 
.A(n_6484),
.B(n_4914),
.Y(n_6977)
);

CKINVDCx5p33_ASAP7_75t_R g6978 ( 
.A(n_6463),
.Y(n_6978)
);

BUFx2_ASAP7_75t_L g6979 ( 
.A(n_6386),
.Y(n_6979)
);

NOR2xp67_ASAP7_75t_L g6980 ( 
.A(n_6475),
.B(n_3379),
.Y(n_6980)
);

NAND2xp33_ASAP7_75t_R g6981 ( 
.A(n_6413),
.B(n_3875),
.Y(n_6981)
);

AND2x4_ASAP7_75t_L g6982 ( 
.A(n_6348),
.B(n_4081),
.Y(n_6982)
);

NAND2xp33_ASAP7_75t_SL g6983 ( 
.A(n_6510),
.B(n_4920),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6389),
.Y(n_6984)
);

HB1xp67_ASAP7_75t_L g6985 ( 
.A(n_6274),
.Y(n_6985)
);

NOR2xp33_ASAP7_75t_L g6986 ( 
.A(n_6505),
.B(n_3876),
.Y(n_6986)
);

CKINVDCx5p33_ASAP7_75t_R g6987 ( 
.A(n_6470),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6395),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6278),
.B(n_4988),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6364),
.Y(n_6990)
);

NOR2xp33_ASAP7_75t_R g6991 ( 
.A(n_6480),
.B(n_6486),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6371),
.Y(n_6992)
);

CKINVDCx20_ASAP7_75t_R g6993 ( 
.A(n_6488),
.Y(n_6993)
);

INVx2_ASAP7_75t_L g6994 ( 
.A(n_6119),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6309),
.Y(n_6995)
);

INVx2_ASAP7_75t_L g6996 ( 
.A(n_6418),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6073),
.Y(n_6997)
);

OAI21x1_ASAP7_75t_L g6998 ( 
.A1(n_6543),
.A2(n_4833),
.B(n_4819),
.Y(n_6998)
);

NOR2xp33_ASAP7_75t_L g6999 ( 
.A(n_6528),
.B(n_6555),
.Y(n_6999)
);

XNOR2xp5_ASAP7_75t_L g7000 ( 
.A(n_6134),
.B(n_4930),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6162),
.Y(n_7001)
);

INVx1_ASAP7_75t_L g7002 ( 
.A(n_6239),
.Y(n_7002)
);

CKINVDCx20_ASAP7_75t_R g7003 ( 
.A(n_6489),
.Y(n_7003)
);

INVxp67_ASAP7_75t_SL g7004 ( 
.A(n_6074),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6139),
.Y(n_7005)
);

BUFx3_ASAP7_75t_L g7006 ( 
.A(n_6004),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_6429),
.Y(n_7007)
);

CKINVDCx5p33_ASAP7_75t_R g7008 ( 
.A(n_6471),
.Y(n_7008)
);

BUFx6f_ASAP7_75t_L g7009 ( 
.A(n_6246),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6313),
.Y(n_7010)
);

AND2x2_ASAP7_75t_L g7011 ( 
.A(n_6360),
.B(n_4988),
.Y(n_7011)
);

INVx2_ASAP7_75t_L g7012 ( 
.A(n_6146),
.Y(n_7012)
);

AND2x2_ASAP7_75t_L g7013 ( 
.A(n_6384),
.B(n_4992),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6170),
.Y(n_7014)
);

CKINVDCx5p33_ASAP7_75t_R g7015 ( 
.A(n_6472),
.Y(n_7015)
);

OAI21x1_ASAP7_75t_L g7016 ( 
.A1(n_6561),
.A2(n_4859),
.B(n_4835),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6190),
.Y(n_7017)
);

INVx2_ASAP7_75t_L g7018 ( 
.A(n_6224),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6264),
.Y(n_7019)
);

CKINVDCx5p33_ASAP7_75t_R g7020 ( 
.A(n_6493),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6297),
.Y(n_7021)
);

CKINVDCx8_ASAP7_75t_R g7022 ( 
.A(n_6386),
.Y(n_7022)
);

HB1xp67_ASAP7_75t_L g7023 ( 
.A(n_6444),
.Y(n_7023)
);

CKINVDCx5p33_ASAP7_75t_R g7024 ( 
.A(n_6217),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6302),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6326),
.Y(n_7026)
);

CKINVDCx5p33_ASAP7_75t_R g7027 ( 
.A(n_6331),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6341),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6346),
.Y(n_7029)
);

CKINVDCx5p33_ASAP7_75t_R g7030 ( 
.A(n_6431),
.Y(n_7030)
);

INVx2_ASAP7_75t_L g7031 ( 
.A(n_6082),
.Y(n_7031)
);

CKINVDCx5p33_ASAP7_75t_R g7032 ( 
.A(n_6461),
.Y(n_7032)
);

NAND2xp5_ASAP7_75t_L g7033 ( 
.A(n_6225),
.B(n_6230),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6407),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6408),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6084),
.Y(n_7036)
);

BUFx10_ASAP7_75t_L g7037 ( 
.A(n_6177),
.Y(n_7037)
);

BUFx6f_ASAP7_75t_L g7038 ( 
.A(n_6255),
.Y(n_7038)
);

CKINVDCx5p33_ASAP7_75t_R g7039 ( 
.A(n_6467),
.Y(n_7039)
);

BUFx2_ASAP7_75t_L g7040 ( 
.A(n_6397),
.Y(n_7040)
);

NAND2xp5_ASAP7_75t_L g7041 ( 
.A(n_6130),
.B(n_6174),
.Y(n_7041)
);

INVx3_ASAP7_75t_L g7042 ( 
.A(n_6262),
.Y(n_7042)
);

CKINVDCx5p33_ASAP7_75t_R g7043 ( 
.A(n_6032),
.Y(n_7043)
);

NAND2xp5_ASAP7_75t_L g7044 ( 
.A(n_6270),
.B(n_3878),
.Y(n_7044)
);

CKINVDCx5p33_ASAP7_75t_R g7045 ( 
.A(n_6441),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6314),
.Y(n_7046)
);

CKINVDCx5p33_ASAP7_75t_R g7047 ( 
.A(n_6469),
.Y(n_7047)
);

NOR2x1_ASAP7_75t_L g7048 ( 
.A(n_6362),
.B(n_4990),
.Y(n_7048)
);

CKINVDCx5p33_ASAP7_75t_R g7049 ( 
.A(n_6438),
.Y(n_7049)
);

AND2x2_ASAP7_75t_SL g7050 ( 
.A(n_6477),
.B(n_4872),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6336),
.Y(n_7051)
);

INVx2_ASAP7_75t_L g7052 ( 
.A(n_6352),
.Y(n_7052)
);

BUFx6f_ASAP7_75t_L g7053 ( 
.A(n_6268),
.Y(n_7053)
);

AND2x4_ASAP7_75t_L g7054 ( 
.A(n_6153),
.B(n_4084),
.Y(n_7054)
);

INVx2_ASAP7_75t_L g7055 ( 
.A(n_6358),
.Y(n_7055)
);

CKINVDCx16_ASAP7_75t_R g7056 ( 
.A(n_6442),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6339),
.Y(n_7057)
);

CKINVDCx16_ASAP7_75t_R g7058 ( 
.A(n_6345),
.Y(n_7058)
);

CKINVDCx5p33_ASAP7_75t_R g7059 ( 
.A(n_6446),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6342),
.Y(n_7060)
);

INVx2_ASAP7_75t_L g7061 ( 
.A(n_6381),
.Y(n_7061)
);

INVx2_ASAP7_75t_L g7062 ( 
.A(n_6388),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6281),
.B(n_3879),
.Y(n_7063)
);

INVx2_ASAP7_75t_L g7064 ( 
.A(n_6402),
.Y(n_7064)
);

CKINVDCx20_ASAP7_75t_R g7065 ( 
.A(n_6412),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_6276),
.Y(n_7066)
);

AND2x2_ASAP7_75t_L g7067 ( 
.A(n_6355),
.B(n_4999),
.Y(n_7067)
);

BUFx6f_ASAP7_75t_L g7068 ( 
.A(n_6279),
.Y(n_7068)
);

AND2x4_ASAP7_75t_L g7069 ( 
.A(n_6289),
.B(n_4087),
.Y(n_7069)
);

CKINVDCx20_ASAP7_75t_R g7070 ( 
.A(n_6452),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_6286),
.Y(n_7071)
);

HB1xp67_ASAP7_75t_L g7072 ( 
.A(n_6422),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6269),
.Y(n_7073)
);

NAND2xp33_ASAP7_75t_R g7074 ( 
.A(n_6425),
.B(n_3882),
.Y(n_7074)
);

CKINVDCx5p33_ASAP7_75t_R g7075 ( 
.A(n_6521),
.Y(n_7075)
);

CKINVDCx20_ASAP7_75t_R g7076 ( 
.A(n_6306),
.Y(n_7076)
);

CKINVDCx5p33_ASAP7_75t_R g7077 ( 
.A(n_6546),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_L g7078 ( 
.A(n_6288),
.B(n_3885),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6152),
.Y(n_7079)
);

CKINVDCx5p33_ASAP7_75t_R g7080 ( 
.A(n_6548),
.Y(n_7080)
);

BUFx2_ASAP7_75t_L g7081 ( 
.A(n_6426),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_6205),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6214),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6231),
.Y(n_7084)
);

AND2x4_ASAP7_75t_L g7085 ( 
.A(n_6310),
.B(n_4092),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6254),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6257),
.Y(n_7087)
);

HB1xp67_ASAP7_75t_L g7088 ( 
.A(n_6329),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6291),
.B(n_3887),
.Y(n_7089)
);

INVx3_ASAP7_75t_L g7090 ( 
.A(n_6330),
.Y(n_7090)
);

BUFx6f_ASAP7_75t_L g7091 ( 
.A(n_6335),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6353),
.Y(n_7092)
);

AND2x4_ASAP7_75t_L g7093 ( 
.A(n_6347),
.B(n_4100),
.Y(n_7093)
);

INVx2_ASAP7_75t_L g7094 ( 
.A(n_6405),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6200),
.Y(n_7095)
);

AND2x6_ASAP7_75t_L g7096 ( 
.A(n_6164),
.B(n_4102),
.Y(n_7096)
);

INVx3_ASAP7_75t_L g7097 ( 
.A(n_6022),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_6051),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6272),
.Y(n_7099)
);

BUFx10_ASAP7_75t_L g7100 ( 
.A(n_6359),
.Y(n_7100)
);

CKINVDCx5p33_ASAP7_75t_R g7101 ( 
.A(n_6563),
.Y(n_7101)
);

INVx3_ASAP7_75t_L g7102 ( 
.A(n_6028),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6283),
.Y(n_7103)
);

AND2x6_ASAP7_75t_L g7104 ( 
.A(n_6169),
.B(n_4106),
.Y(n_7104)
);

AND2x2_ASAP7_75t_L g7105 ( 
.A(n_6363),
.B(n_4999),
.Y(n_7105)
);

INVx4_ASAP7_75t_L g7106 ( 
.A(n_6287),
.Y(n_7106)
);

HB1xp67_ASAP7_75t_L g7107 ( 
.A(n_6083),
.Y(n_7107)
);

NOR2xp33_ASAP7_75t_L g7108 ( 
.A(n_6071),
.B(n_3889),
.Y(n_7108)
);

CKINVDCx20_ASAP7_75t_R g7109 ( 
.A(n_6370),
.Y(n_7109)
);

AO21x2_ASAP7_75t_L g7110 ( 
.A1(n_6430),
.A2(n_4114),
.B(n_4113),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6296),
.Y(n_7111)
);

INVx3_ASAP7_75t_L g7112 ( 
.A(n_6115),
.Y(n_7112)
);

BUFx6f_ASAP7_75t_L g7113 ( 
.A(n_6365),
.Y(n_7113)
);

CKINVDCx20_ASAP7_75t_R g7114 ( 
.A(n_6207),
.Y(n_7114)
);

NOR2xp33_ASAP7_75t_R g7115 ( 
.A(n_6303),
.B(n_4953),
.Y(n_7115)
);

AND2x4_ASAP7_75t_L g7116 ( 
.A(n_6067),
.B(n_4116),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6142),
.Y(n_7117)
);

INVx2_ASAP7_75t_L g7118 ( 
.A(n_6059),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_6097),
.Y(n_7119)
);

NAND2xp5_ASAP7_75t_SL g7120 ( 
.A(n_6057),
.B(n_3890),
.Y(n_7120)
);

AND2x4_ASAP7_75t_L g7121 ( 
.A(n_6141),
.B(n_4119),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_L g7122 ( 
.A(n_6137),
.B(n_3892),
.Y(n_7122)
);

NOR2xp33_ASAP7_75t_L g7123 ( 
.A(n_6036),
.B(n_3893),
.Y(n_7123)
);

NAND2xp5_ASAP7_75t_SL g7124 ( 
.A(n_5992),
.B(n_3894),
.Y(n_7124)
);

INVxp67_ASAP7_75t_L g7125 ( 
.A(n_6258),
.Y(n_7125)
);

INVxp67_ASAP7_75t_L g7126 ( 
.A(n_6427),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6023),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6025),
.Y(n_7128)
);

AND2x2_ASAP7_75t_L g7129 ( 
.A(n_6155),
.B(n_4979),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_6580),
.Y(n_7130)
);

INVx3_ASAP7_75t_L g7131 ( 
.A(n_6926),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6568),
.Y(n_7132)
);

INVx2_ASAP7_75t_L g7133 ( 
.A(n_6588),
.Y(n_7133)
);

OAI21xp33_ASAP7_75t_SL g7134 ( 
.A1(n_7117),
.A2(n_6149),
.B(n_4123),
.Y(n_7134)
);

BUFx10_ASAP7_75t_L g7135 ( 
.A(n_6576),
.Y(n_7135)
);

INVx2_ASAP7_75t_L g7136 ( 
.A(n_6590),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_6596),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6597),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6602),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_6610),
.Y(n_7140)
);

NAND2xp33_ASAP7_75t_R g7141 ( 
.A(n_6977),
.B(n_6049),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6616),
.Y(n_7142)
);

NAND2xp33_ASAP7_75t_SL g7143 ( 
.A(n_6796),
.B(n_6186),
.Y(n_7143)
);

BUFx10_ASAP7_75t_L g7144 ( 
.A(n_6840),
.Y(n_7144)
);

INVx5_ASAP7_75t_L g7145 ( 
.A(n_6803),
.Y(n_7145)
);

CKINVDCx5p33_ASAP7_75t_R g7146 ( 
.A(n_6586),
.Y(n_7146)
);

INVx2_ASAP7_75t_L g7147 ( 
.A(n_6637),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6575),
.Y(n_7148)
);

INVx2_ASAP7_75t_L g7149 ( 
.A(n_6642),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_SL g7150 ( 
.A(n_6845),
.B(n_6742),
.Y(n_7150)
);

BUFx10_ASAP7_75t_L g7151 ( 
.A(n_6599),
.Y(n_7151)
);

BUFx6f_ASAP7_75t_SL g7152 ( 
.A(n_6871),
.Y(n_7152)
);

NOR2xp33_ASAP7_75t_L g7153 ( 
.A(n_6573),
.B(n_5013),
.Y(n_7153)
);

CKINVDCx5p33_ASAP7_75t_R g7154 ( 
.A(n_6603),
.Y(n_7154)
);

AOI22xp33_ASAP7_75t_L g7155 ( 
.A1(n_6856),
.A2(n_6189),
.B1(n_6037),
.B2(n_4903),
.Y(n_7155)
);

NOR2xp33_ASAP7_75t_L g7156 ( 
.A(n_6891),
.B(n_3896),
.Y(n_7156)
);

AND3x2_ASAP7_75t_L g7157 ( 
.A(n_6594),
.B(n_4126),
.C(n_4120),
.Y(n_7157)
);

NAND2xp5_ASAP7_75t_SL g7158 ( 
.A(n_6631),
.B(n_3897),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6846),
.B(n_3899),
.Y(n_7159)
);

AOI21x1_ASAP7_75t_L g7160 ( 
.A1(n_6849),
.A2(n_4131),
.B(n_4129),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6577),
.Y(n_7161)
);

INVx3_ASAP7_75t_L g7162 ( 
.A(n_6926),
.Y(n_7162)
);

INVx2_ASAP7_75t_L g7163 ( 
.A(n_6647),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_6836),
.B(n_3901),
.Y(n_7164)
);

NAND3xp33_ASAP7_75t_L g7165 ( 
.A(n_6916),
.B(n_7123),
.C(n_7108),
.Y(n_7165)
);

INVx6_ASAP7_75t_L g7166 ( 
.A(n_6925),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_SL g7167 ( 
.A(n_7050),
.B(n_3905),
.Y(n_7167)
);

NAND2xp5_ASAP7_75t_SL g7168 ( 
.A(n_6999),
.B(n_3906),
.Y(n_7168)
);

INVx3_ASAP7_75t_L g7169 ( 
.A(n_6944),
.Y(n_7169)
);

BUFx3_ASAP7_75t_L g7170 ( 
.A(n_6618),
.Y(n_7170)
);

INVx2_ASAP7_75t_SL g7171 ( 
.A(n_6591),
.Y(n_7171)
);

AOI21x1_ASAP7_75t_L g7172 ( 
.A1(n_7127),
.A2(n_4143),
.B(n_4132),
.Y(n_7172)
);

NAND2xp33_ASAP7_75t_SL g7173 ( 
.A(n_6805),
.B(n_3907),
.Y(n_7173)
);

BUFx10_ASAP7_75t_L g7174 ( 
.A(n_6605),
.Y(n_7174)
);

BUFx3_ASAP7_75t_L g7175 ( 
.A(n_6739),
.Y(n_7175)
);

AND2x6_ASAP7_75t_L g7176 ( 
.A(n_7066),
.B(n_4147),
.Y(n_7176)
);

BUFx6f_ASAP7_75t_L g7177 ( 
.A(n_6570),
.Y(n_7177)
);

INVx2_ASAP7_75t_SL g7178 ( 
.A(n_6775),
.Y(n_7178)
);

CKINVDCx20_ASAP7_75t_R g7179 ( 
.A(n_6651),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6579),
.Y(n_7180)
);

AOI22xp33_ASAP7_75t_L g7181 ( 
.A1(n_6837),
.A2(n_4908),
.B1(n_4915),
.B2(n_4888),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6650),
.Y(n_7182)
);

INVx2_ASAP7_75t_L g7183 ( 
.A(n_6656),
.Y(n_7183)
);

INVx1_ASAP7_75t_SL g7184 ( 
.A(n_6783),
.Y(n_7184)
);

INVx8_ASAP7_75t_L g7185 ( 
.A(n_6722),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6657),
.Y(n_7186)
);

NAND2xp5_ASAP7_75t_L g7187 ( 
.A(n_7010),
.B(n_3909),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_6583),
.Y(n_7188)
);

CKINVDCx20_ASAP7_75t_R g7189 ( 
.A(n_6686),
.Y(n_7189)
);

NOR2xp33_ASAP7_75t_L g7190 ( 
.A(n_6720),
.B(n_3911),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_SL g7191 ( 
.A(n_6924),
.B(n_3918),
.Y(n_7191)
);

INVx3_ASAP7_75t_L g7192 ( 
.A(n_6944),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_6589),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_6606),
.Y(n_7194)
);

NAND2xp33_ASAP7_75t_R g7195 ( 
.A(n_6748),
.B(n_3921),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_6607),
.Y(n_7196)
);

INVx3_ASAP7_75t_L g7197 ( 
.A(n_6952),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_L g7198 ( 
.A(n_7046),
.B(n_3928),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6608),
.Y(n_7199)
);

INVx1_ASAP7_75t_SL g7200 ( 
.A(n_6670),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6609),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6614),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_6659),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_6615),
.Y(n_7204)
);

NAND2xp5_ASAP7_75t_SL g7205 ( 
.A(n_6929),
.B(n_3930),
.Y(n_7205)
);

INVx2_ASAP7_75t_L g7206 ( 
.A(n_6665),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6625),
.Y(n_7207)
);

BUFx2_ASAP7_75t_L g7208 ( 
.A(n_6600),
.Y(n_7208)
);

NOR2xp33_ASAP7_75t_L g7209 ( 
.A(n_7125),
.B(n_3932),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_6626),
.Y(n_7210)
);

INVx2_ASAP7_75t_L g7211 ( 
.A(n_6667),
.Y(n_7211)
);

INVx2_ASAP7_75t_L g7212 ( 
.A(n_6677),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6628),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_SL g7214 ( 
.A(n_6931),
.B(n_3943),
.Y(n_7214)
);

NOR2xp33_ASAP7_75t_L g7215 ( 
.A(n_7024),
.B(n_3944),
.Y(n_7215)
);

INVx2_ASAP7_75t_SL g7216 ( 
.A(n_6633),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6634),
.Y(n_7217)
);

BUFx3_ASAP7_75t_L g7218 ( 
.A(n_6789),
.Y(n_7218)
);

INVx2_ASAP7_75t_L g7219 ( 
.A(n_6636),
.Y(n_7219)
);

AND2x2_ASAP7_75t_L g7220 ( 
.A(n_6680),
.B(n_3945),
.Y(n_7220)
);

INVx5_ASAP7_75t_L g7221 ( 
.A(n_6852),
.Y(n_7221)
);

INVx3_ASAP7_75t_L g7222 ( 
.A(n_6952),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6639),
.Y(n_7223)
);

INVx2_ASAP7_75t_L g7224 ( 
.A(n_6652),
.Y(n_7224)
);

AOI21x1_ASAP7_75t_L g7225 ( 
.A1(n_6571),
.A2(n_4155),
.B(n_4150),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_6654),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_6662),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6663),
.Y(n_7228)
);

INVx2_ASAP7_75t_SL g7229 ( 
.A(n_6617),
.Y(n_7229)
);

AND2x4_ASAP7_75t_L g7230 ( 
.A(n_6877),
.B(n_4157),
.Y(n_7230)
);

INVx2_ASAP7_75t_L g7231 ( 
.A(n_6664),
.Y(n_7231)
);

INVx2_ASAP7_75t_SL g7232 ( 
.A(n_6703),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_6666),
.Y(n_7233)
);

INVx2_ASAP7_75t_SL g7234 ( 
.A(n_6963),
.Y(n_7234)
);

INVx4_ASAP7_75t_L g7235 ( 
.A(n_6725),
.Y(n_7235)
);

BUFx3_ASAP7_75t_L g7236 ( 
.A(n_6794),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_6669),
.Y(n_7237)
);

NAND2xp33_ASAP7_75t_L g7238 ( 
.A(n_6812),
.B(n_3947),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_6676),
.Y(n_7239)
);

AND2x2_ASAP7_75t_L g7240 ( 
.A(n_6692),
.B(n_3953),
.Y(n_7240)
);

INVx1_ASAP7_75t_SL g7241 ( 
.A(n_6875),
.Y(n_7241)
);

NOR3xp33_ASAP7_75t_L g7242 ( 
.A(n_6587),
.B(n_3956),
.C(n_3955),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_6689),
.Y(n_7243)
);

INVx2_ASAP7_75t_L g7244 ( 
.A(n_6691),
.Y(n_7244)
);

INVx4_ASAP7_75t_L g7245 ( 
.A(n_6735),
.Y(n_7245)
);

BUFx10_ASAP7_75t_L g7246 ( 
.A(n_6619),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_6695),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_SL g7248 ( 
.A(n_6938),
.B(n_3959),
.Y(n_7248)
);

CKINVDCx5p33_ASAP7_75t_R g7249 ( 
.A(n_6622),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_6700),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_6708),
.Y(n_7251)
);

INVx2_ASAP7_75t_L g7252 ( 
.A(n_6711),
.Y(n_7252)
);

INVx3_ASAP7_75t_L g7253 ( 
.A(n_6960),
.Y(n_7253)
);

NOR2xp33_ASAP7_75t_L g7254 ( 
.A(n_6688),
.B(n_3961),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_6712),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_6713),
.Y(n_7256)
);

INVx2_ASAP7_75t_L g7257 ( 
.A(n_6714),
.Y(n_7257)
);

CKINVDCx6p67_ASAP7_75t_R g7258 ( 
.A(n_6858),
.Y(n_7258)
);

INVx2_ASAP7_75t_SL g7259 ( 
.A(n_6964),
.Y(n_7259)
);

NOR2xp33_ASAP7_75t_L g7260 ( 
.A(n_6727),
.B(n_3963),
.Y(n_7260)
);

INVx2_ASAP7_75t_L g7261 ( 
.A(n_6715),
.Y(n_7261)
);

NAND2xp5_ASAP7_75t_L g7262 ( 
.A(n_7051),
.B(n_3964),
.Y(n_7262)
);

NOR2xp33_ASAP7_75t_L g7263 ( 
.A(n_6888),
.B(n_3970),
.Y(n_7263)
);

NAND2xp5_ASAP7_75t_L g7264 ( 
.A(n_7057),
.B(n_3973),
.Y(n_7264)
);

INVx3_ASAP7_75t_L g7265 ( 
.A(n_6960),
.Y(n_7265)
);

AOI22xp33_ASAP7_75t_L g7266 ( 
.A1(n_7060),
.A2(n_4929),
.B1(n_4932),
.B2(n_4919),
.Y(n_7266)
);

NAND2xp5_ASAP7_75t_L g7267 ( 
.A(n_7073),
.B(n_3976),
.Y(n_7267)
);

BUFx3_ASAP7_75t_L g7268 ( 
.A(n_6855),
.Y(n_7268)
);

INVx2_ASAP7_75t_L g7269 ( 
.A(n_6716),
.Y(n_7269)
);

AND2x2_ASAP7_75t_SL g7270 ( 
.A(n_6806),
.B(n_4934),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_6719),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6721),
.Y(n_7272)
);

INVx3_ASAP7_75t_L g7273 ( 
.A(n_6965),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_SL g7274 ( 
.A(n_6940),
.B(n_3979),
.Y(n_7274)
);

INVx8_ASAP7_75t_L g7275 ( 
.A(n_6737),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_SL g7276 ( 
.A(n_6946),
.B(n_6598),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_SL g7277 ( 
.A(n_6569),
.B(n_3981),
.Y(n_7277)
);

NAND2xp5_ASAP7_75t_SL g7278 ( 
.A(n_6958),
.B(n_3982),
.Y(n_7278)
);

INVx2_ASAP7_75t_SL g7279 ( 
.A(n_6985),
.Y(n_7279)
);

OR2x2_ASAP7_75t_L g7280 ( 
.A(n_7040),
.B(n_3989),
.Y(n_7280)
);

AND2x2_ASAP7_75t_SL g7281 ( 
.A(n_6869),
.B(n_4945),
.Y(n_7281)
);

INVx2_ASAP7_75t_SL g7282 ( 
.A(n_6863),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_6729),
.Y(n_7283)
);

INVx3_ASAP7_75t_L g7284 ( 
.A(n_6965),
.Y(n_7284)
);

INVx3_ASAP7_75t_L g7285 ( 
.A(n_7009),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_SL g7286 ( 
.A(n_6972),
.B(n_3995),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6730),
.Y(n_7287)
);

BUFx6f_ASAP7_75t_L g7288 ( 
.A(n_6570),
.Y(n_7288)
);

INVx2_ASAP7_75t_L g7289 ( 
.A(n_6733),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_SL g7290 ( 
.A(n_6978),
.B(n_3996),
.Y(n_7290)
);

INVx5_ASAP7_75t_L g7291 ( 
.A(n_6937),
.Y(n_7291)
);

INVx1_ASAP7_75t_SL g7292 ( 
.A(n_6949),
.Y(n_7292)
);

INVx1_ASAP7_75t_SL g7293 ( 
.A(n_6833),
.Y(n_7293)
);

INVx5_ASAP7_75t_L g7294 ( 
.A(n_6574),
.Y(n_7294)
);

NAND2xp33_ASAP7_75t_L g7295 ( 
.A(n_6813),
.B(n_3999),
.Y(n_7295)
);

INVx2_ASAP7_75t_L g7296 ( 
.A(n_6747),
.Y(n_7296)
);

CKINVDCx5p33_ASAP7_75t_R g7297 ( 
.A(n_6623),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6750),
.Y(n_7298)
);

INVxp67_ASAP7_75t_SL g7299 ( 
.A(n_6863),
.Y(n_7299)
);

NAND2xp5_ASAP7_75t_SL g7300 ( 
.A(n_6987),
.B(n_4000),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_L g7301 ( 
.A(n_7034),
.B(n_4004),
.Y(n_7301)
);

NOR2x1p5_ASAP7_75t_L g7302 ( 
.A(n_6741),
.B(n_4005),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_6752),
.Y(n_7303)
);

NAND2xp5_ASAP7_75t_L g7304 ( 
.A(n_7035),
.B(n_6653),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_6756),
.Y(n_7305)
);

NAND2xp5_ASAP7_75t_L g7306 ( 
.A(n_7082),
.B(n_4006),
.Y(n_7306)
);

INVx2_ASAP7_75t_SL g7307 ( 
.A(n_6906),
.Y(n_7307)
);

NOR2xp33_ASAP7_75t_L g7308 ( 
.A(n_7049),
.B(n_4008),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_L g7309 ( 
.A(n_7083),
.B(n_7084),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_7086),
.B(n_4010),
.Y(n_7310)
);

INVx1_ASAP7_75t_L g7311 ( 
.A(n_6759),
.Y(n_7311)
);

INVx2_ASAP7_75t_L g7312 ( 
.A(n_6761),
.Y(n_7312)
);

NOR2xp33_ASAP7_75t_L g7313 ( 
.A(n_7059),
.B(n_4013),
.Y(n_7313)
);

INVx1_ASAP7_75t_L g7314 ( 
.A(n_6767),
.Y(n_7314)
);

AND2x2_ASAP7_75t_L g7315 ( 
.A(n_6710),
.B(n_4015),
.Y(n_7315)
);

INVx2_ASAP7_75t_L g7316 ( 
.A(n_6769),
.Y(n_7316)
);

INVx2_ASAP7_75t_L g7317 ( 
.A(n_6772),
.Y(n_7317)
);

NAND2xp5_ASAP7_75t_SL g7318 ( 
.A(n_7008),
.B(n_4017),
.Y(n_7318)
);

INVx4_ASAP7_75t_L g7319 ( 
.A(n_6744),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_6784),
.Y(n_7320)
);

INVx3_ASAP7_75t_L g7321 ( 
.A(n_7009),
.Y(n_7321)
);

BUFx10_ASAP7_75t_L g7322 ( 
.A(n_6624),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_L g7323 ( 
.A(n_7087),
.B(n_6578),
.Y(n_7323)
);

BUFx3_ASAP7_75t_L g7324 ( 
.A(n_6581),
.Y(n_7324)
);

INVxp67_ASAP7_75t_L g7325 ( 
.A(n_6873),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_6786),
.Y(n_7326)
);

INVx2_ASAP7_75t_L g7327 ( 
.A(n_6791),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_6797),
.Y(n_7328)
);

AND3x2_ASAP7_75t_L g7329 ( 
.A(n_6903),
.B(n_4165),
.C(n_4160),
.Y(n_7329)
);

INVx2_ASAP7_75t_L g7330 ( 
.A(n_6798),
.Y(n_7330)
);

CKINVDCx5p33_ASAP7_75t_R g7331 ( 
.A(n_6627),
.Y(n_7331)
);

INVx2_ASAP7_75t_L g7332 ( 
.A(n_6800),
.Y(n_7332)
);

INVx2_ASAP7_75t_L g7333 ( 
.A(n_6808),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_L g7334 ( 
.A(n_6766),
.B(n_4021),
.Y(n_7334)
);

INVx3_ASAP7_75t_L g7335 ( 
.A(n_7038),
.Y(n_7335)
);

CKINVDCx5p33_ASAP7_75t_R g7336 ( 
.A(n_6630),
.Y(n_7336)
);

BUFx3_ASAP7_75t_L g7337 ( 
.A(n_6581),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_6811),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6818),
.Y(n_7339)
);

INVx2_ASAP7_75t_SL g7340 ( 
.A(n_6906),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6819),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_6820),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_6740),
.B(n_4022),
.Y(n_7343)
);

INVx2_ASAP7_75t_L g7344 ( 
.A(n_6821),
.Y(n_7344)
);

NOR2xp33_ASAP7_75t_L g7345 ( 
.A(n_7015),
.B(n_4030),
.Y(n_7345)
);

NAND2xp5_ASAP7_75t_L g7346 ( 
.A(n_6809),
.B(n_4033),
.Y(n_7346)
);

AOI22xp33_ASAP7_75t_L g7347 ( 
.A1(n_7071),
.A2(n_5001),
.B1(n_4980),
.B2(n_4174),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_6823),
.Y(n_7348)
);

INVx1_ASAP7_75t_SL g7349 ( 
.A(n_6776),
.Y(n_7349)
);

INVx1_ASAP7_75t_L g7350 ( 
.A(n_6829),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_SL g7351 ( 
.A(n_6826),
.B(n_4034),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6838),
.Y(n_7352)
);

AND2x2_ASAP7_75t_L g7353 ( 
.A(n_6792),
.B(n_4039),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_6839),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_6842),
.Y(n_7355)
);

INVx2_ASAP7_75t_L g7356 ( 
.A(n_6848),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_6822),
.Y(n_7357)
);

OAI22xp33_ASAP7_75t_L g7358 ( 
.A1(n_7045),
.A2(n_4043),
.B1(n_4045),
.B2(n_4040),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_6850),
.Y(n_7359)
);

INVx4_ASAP7_75t_L g7360 ( 
.A(n_6751),
.Y(n_7360)
);

NOR2xp33_ASAP7_75t_L g7361 ( 
.A(n_6876),
.B(n_4046),
.Y(n_7361)
);

INVxp67_ASAP7_75t_SL g7362 ( 
.A(n_6923),
.Y(n_7362)
);

AND2x2_ASAP7_75t_L g7363 ( 
.A(n_6844),
.B(n_4047),
.Y(n_7363)
);

NOR2xp33_ASAP7_75t_L g7364 ( 
.A(n_6880),
.B(n_4048),
.Y(n_7364)
);

INVx2_ASAP7_75t_L g7365 ( 
.A(n_6854),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_6861),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_6718),
.B(n_4049),
.Y(n_7367)
);

AND3x2_ASAP7_75t_L g7368 ( 
.A(n_6942),
.B(n_4176),
.C(n_4173),
.Y(n_7368)
);

NAND2xp5_ASAP7_75t_L g7369 ( 
.A(n_7044),
.B(n_4052),
.Y(n_7369)
);

INVx2_ASAP7_75t_SL g7370 ( 
.A(n_6923),
.Y(n_7370)
);

INVx2_ASAP7_75t_SL g7371 ( 
.A(n_6612),
.Y(n_7371)
);

OAI22xp33_ASAP7_75t_L g7372 ( 
.A1(n_6885),
.A2(n_4058),
.B1(n_4063),
.B2(n_4056),
.Y(n_7372)
);

NAND2xp5_ASAP7_75t_L g7373 ( 
.A(n_7063),
.B(n_4067),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_L g7374 ( 
.A(n_7078),
.B(n_4068),
.Y(n_7374)
);

INVx2_ASAP7_75t_L g7375 ( 
.A(n_6866),
.Y(n_7375)
);

BUFx3_ASAP7_75t_L g7376 ( 
.A(n_6592),
.Y(n_7376)
);

NOR2xp33_ASAP7_75t_L g7377 ( 
.A(n_6611),
.B(n_4070),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_6879),
.Y(n_7378)
);

BUFx2_ASAP7_75t_L g7379 ( 
.A(n_6774),
.Y(n_7379)
);

INVx2_ASAP7_75t_L g7380 ( 
.A(n_6693),
.Y(n_7380)
);

INVx2_ASAP7_75t_L g7381 ( 
.A(n_6694),
.Y(n_7381)
);

INVx4_ASAP7_75t_L g7382 ( 
.A(n_6762),
.Y(n_7382)
);

BUFx3_ASAP7_75t_L g7383 ( 
.A(n_6592),
.Y(n_7383)
);

INVx2_ASAP7_75t_L g7384 ( 
.A(n_6717),
.Y(n_7384)
);

INVx2_ASAP7_75t_SL g7385 ( 
.A(n_7069),
.Y(n_7385)
);

NOR2xp33_ASAP7_75t_L g7386 ( 
.A(n_6745),
.B(n_4071),
.Y(n_7386)
);

INVx2_ASAP7_75t_L g7387 ( 
.A(n_6726),
.Y(n_7387)
);

INVx2_ASAP7_75t_L g7388 ( 
.A(n_6731),
.Y(n_7388)
);

INVx1_ASAP7_75t_L g7389 ( 
.A(n_6883),
.Y(n_7389)
);

AOI22xp33_ASAP7_75t_L g7390 ( 
.A1(n_6995),
.A2(n_4189),
.B1(n_4191),
.B2(n_4187),
.Y(n_7390)
);

NOR2x1p5_ASAP7_75t_L g7391 ( 
.A(n_6828),
.B(n_6831),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_6734),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_6887),
.Y(n_7393)
);

AO22x2_ASAP7_75t_L g7394 ( 
.A1(n_7129),
.A2(n_4198),
.B1(n_4202),
.B2(n_4193),
.Y(n_7394)
);

INVx2_ASAP7_75t_L g7395 ( 
.A(n_6743),
.Y(n_7395)
);

NAND2xp33_ASAP7_75t_L g7396 ( 
.A(n_6832),
.B(n_4073),
.Y(n_7396)
);

BUFx2_ASAP7_75t_L g7397 ( 
.A(n_7070),
.Y(n_7397)
);

CKINVDCx5p33_ASAP7_75t_R g7398 ( 
.A(n_6632),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_6889),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6892),
.Y(n_7400)
);

NAND2xp33_ASAP7_75t_SL g7401 ( 
.A(n_7075),
.B(n_7077),
.Y(n_7401)
);

HB1xp67_ASAP7_75t_L g7402 ( 
.A(n_7023),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_L g7403 ( 
.A(n_7089),
.B(n_4074),
.Y(n_7403)
);

NAND2xp5_ASAP7_75t_L g7404 ( 
.A(n_6701),
.B(n_4075),
.Y(n_7404)
);

NAND2xp5_ASAP7_75t_SL g7405 ( 
.A(n_6858),
.B(n_4076),
.Y(n_7405)
);

CKINVDCx5p33_ASAP7_75t_R g7406 ( 
.A(n_6638),
.Y(n_7406)
);

INVx8_ASAP7_75t_L g7407 ( 
.A(n_6763),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_6893),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_6896),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_6905),
.Y(n_7410)
);

NAND2xp5_ASAP7_75t_L g7411 ( 
.A(n_6897),
.B(n_4078),
.Y(n_7411)
);

NAND2xp5_ASAP7_75t_L g7412 ( 
.A(n_6986),
.B(n_4080),
.Y(n_7412)
);

INVx2_ASAP7_75t_L g7413 ( 
.A(n_6749),
.Y(n_7413)
);

NOR2xp33_ASAP7_75t_L g7414 ( 
.A(n_7080),
.B(n_4083),
.Y(n_7414)
);

AND3x2_ASAP7_75t_L g7415 ( 
.A(n_6979),
.B(n_4206),
.C(n_4203),
.Y(n_7415)
);

INVx2_ASAP7_75t_L g7416 ( 
.A(n_6754),
.Y(n_7416)
);

INVx6_ASAP7_75t_L g7417 ( 
.A(n_6976),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_6757),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_6907),
.Y(n_7419)
);

INVxp67_ASAP7_75t_SL g7420 ( 
.A(n_6595),
.Y(n_7420)
);

OAI22xp33_ASAP7_75t_L g7421 ( 
.A1(n_7101),
.A2(n_4088),
.B1(n_4089),
.B2(n_4086),
.Y(n_7421)
);

AND2x6_ASAP7_75t_L g7422 ( 
.A(n_7001),
.B(n_4207),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6908),
.Y(n_7423)
);

INVx2_ASAP7_75t_SL g7424 ( 
.A(n_7085),
.Y(n_7424)
);

INVx2_ASAP7_75t_L g7425 ( 
.A(n_6770),
.Y(n_7425)
);

CKINVDCx5p33_ASAP7_75t_R g7426 ( 
.A(n_6649),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6911),
.Y(n_7427)
);

INVx2_ASAP7_75t_L g7428 ( 
.A(n_6773),
.Y(n_7428)
);

INVx6_ASAP7_75t_L g7429 ( 
.A(n_6595),
.Y(n_7429)
);

AOI21x1_ASAP7_75t_L g7430 ( 
.A1(n_7079),
.A2(n_4220),
.B(n_4217),
.Y(n_7430)
);

AND3x2_ASAP7_75t_L g7431 ( 
.A(n_6966),
.B(n_7081),
.C(n_7072),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6919),
.Y(n_7432)
);

NAND2xp5_ASAP7_75t_SL g7433 ( 
.A(n_7115),
.B(n_4091),
.Y(n_7433)
);

NAND2xp5_ASAP7_75t_SL g7434 ( 
.A(n_6980),
.B(n_4093),
.Y(n_7434)
);

INVx2_ASAP7_75t_L g7435 ( 
.A(n_6779),
.Y(n_7435)
);

INVxp67_ASAP7_75t_L g7436 ( 
.A(n_6853),
.Y(n_7436)
);

INVx5_ASAP7_75t_L g7437 ( 
.A(n_6574),
.Y(n_7437)
);

AND2x2_ASAP7_75t_L g7438 ( 
.A(n_6967),
.B(n_4094),
.Y(n_7438)
);

INVx2_ASAP7_75t_L g7439 ( 
.A(n_6781),
.Y(n_7439)
);

NOR2xp33_ASAP7_75t_L g7440 ( 
.A(n_7030),
.B(n_4095),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_6922),
.Y(n_7441)
);

INVxp33_ASAP7_75t_SL g7442 ( 
.A(n_6582),
.Y(n_7442)
);

INVx2_ASAP7_75t_L g7443 ( 
.A(n_6810),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_6933),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_6941),
.Y(n_7445)
);

INVx2_ASAP7_75t_L g7446 ( 
.A(n_6817),
.Y(n_7446)
);

INVx5_ASAP7_75t_L g7447 ( 
.A(n_6574),
.Y(n_7447)
);

OAI22xp5_ASAP7_75t_L g7448 ( 
.A1(n_7032),
.A2(n_7039),
.B1(n_6930),
.B2(n_7099),
.Y(n_7448)
);

INVx2_ASAP7_75t_L g7449 ( 
.A(n_6824),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6943),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_6950),
.Y(n_7451)
);

BUFx6f_ASAP7_75t_L g7452 ( 
.A(n_6643),
.Y(n_7452)
);

OAI22xp33_ASAP7_75t_L g7453 ( 
.A1(n_6953),
.A2(n_4098),
.B1(n_4099),
.B2(n_4096),
.Y(n_7453)
);

INVx2_ASAP7_75t_SL g7454 ( 
.A(n_7093),
.Y(n_7454)
);

NAND2xp33_ASAP7_75t_L g7455 ( 
.A(n_6795),
.B(n_4103),
.Y(n_7455)
);

INVx2_ASAP7_75t_L g7456 ( 
.A(n_6827),
.Y(n_7456)
);

INVx2_ASAP7_75t_L g7457 ( 
.A(n_6835),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_6954),
.Y(n_7458)
);

OAI22xp33_ASAP7_75t_SL g7459 ( 
.A1(n_7126),
.A2(n_4226),
.B1(n_4231),
.B2(n_4223),
.Y(n_7459)
);

OR2x2_ASAP7_75t_L g7460 ( 
.A(n_7058),
.B(n_4104),
.Y(n_7460)
);

OR2x2_ASAP7_75t_L g7461 ( 
.A(n_6802),
.B(n_4105),
.Y(n_7461)
);

INVx3_ASAP7_75t_L g7462 ( 
.A(n_7038),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6955),
.Y(n_7463)
);

BUFx3_ASAP7_75t_L g7464 ( 
.A(n_6643),
.Y(n_7464)
);

OR2x2_ASAP7_75t_L g7465 ( 
.A(n_7056),
.B(n_4108),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_6990),
.B(n_4112),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_6961),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6970),
.Y(n_7468)
);

INVx2_ASAP7_75t_L g7469 ( 
.A(n_6843),
.Y(n_7469)
);

BUFx2_ASAP7_75t_L g7470 ( 
.A(n_6993),
.Y(n_7470)
);

BUFx3_ASAP7_75t_L g7471 ( 
.A(n_6699),
.Y(n_7471)
);

INVx2_ASAP7_75t_L g7472 ( 
.A(n_6868),
.Y(n_7472)
);

HB1xp67_ASAP7_75t_L g7473 ( 
.A(n_6898),
.Y(n_7473)
);

INVx2_ASAP7_75t_L g7474 ( 
.A(n_6870),
.Y(n_7474)
);

NAND2xp33_ASAP7_75t_L g7475 ( 
.A(n_7048),
.B(n_4122),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_6973),
.Y(n_7476)
);

A2O1A1Ixp33_ASAP7_75t_L g7477 ( 
.A1(n_6862),
.A2(n_4239),
.B(n_4250),
.C(n_4237),
.Y(n_7477)
);

AOI22xp33_ASAP7_75t_L g7478 ( 
.A1(n_7002),
.A2(n_4260),
.B1(n_4264),
.B2(n_4251),
.Y(n_7478)
);

XNOR2xp5_ASAP7_75t_L g7479 ( 
.A(n_6572),
.B(n_3380),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_6988),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_SL g7481 ( 
.A(n_6992),
.B(n_4124),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_6878),
.Y(n_7482)
);

NOR2xp33_ASAP7_75t_L g7483 ( 
.A(n_6648),
.B(n_4125),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_6881),
.Y(n_7484)
);

INVx2_ASAP7_75t_L g7485 ( 
.A(n_6886),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_SL g7486 ( 
.A(n_6674),
.B(n_4128),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_6901),
.B(n_4134),
.Y(n_7487)
);

NAND2xp5_ASAP7_75t_SL g7488 ( 
.A(n_7106),
.B(n_4137),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_6920),
.Y(n_7489)
);

INVxp33_ASAP7_75t_L g7490 ( 
.A(n_6760),
.Y(n_7490)
);

BUFx10_ASAP7_75t_L g7491 ( 
.A(n_6655),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_6934),
.B(n_4138),
.Y(n_7492)
);

INVx2_ASAP7_75t_SL g7493 ( 
.A(n_6699),
.Y(n_7493)
);

AO22x2_ASAP7_75t_L g7494 ( 
.A1(n_6658),
.A2(n_4285),
.B1(n_4290),
.B2(n_4273),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_6951),
.Y(n_7495)
);

NAND2xp5_ASAP7_75t_L g7496 ( 
.A(n_6968),
.B(n_4139),
.Y(n_7496)
);

OR2x6_ASAP7_75t_L g7497 ( 
.A(n_7053),
.B(n_4291),
.Y(n_7497)
);

INVx2_ASAP7_75t_L g7498 ( 
.A(n_6969),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_6975),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_6984),
.Y(n_7500)
);

NAND2xp5_ASAP7_75t_L g7501 ( 
.A(n_6679),
.B(n_4142),
.Y(n_7501)
);

NAND2xp5_ASAP7_75t_L g7502 ( 
.A(n_6681),
.B(n_4144),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_6685),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_6917),
.Y(n_7504)
);

NAND2xp5_ASAP7_75t_L g7505 ( 
.A(n_6874),
.B(n_4145),
.Y(n_7505)
);

OR2x6_ASAP7_75t_L g7506 ( 
.A(n_7053),
.B(n_4296),
.Y(n_7506)
);

BUFx6f_ASAP7_75t_L g7507 ( 
.A(n_6706),
.Y(n_7507)
);

BUFx6f_ASAP7_75t_L g7508 ( 
.A(n_6706),
.Y(n_7508)
);

INVx2_ASAP7_75t_L g7509 ( 
.A(n_6997),
.Y(n_7509)
);

NAND2xp5_ASAP7_75t_L g7510 ( 
.A(n_6914),
.B(n_4146),
.Y(n_7510)
);

NAND2xp5_ASAP7_75t_L g7511 ( 
.A(n_7004),
.B(n_4148),
.Y(n_7511)
);

NAND2xp5_ASAP7_75t_L g7512 ( 
.A(n_7103),
.B(n_4149),
.Y(n_7512)
);

NAND2xp5_ASAP7_75t_L g7513 ( 
.A(n_7111),
.B(n_4151),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7031),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7036),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_6994),
.Y(n_7516)
);

INVx3_ASAP7_75t_L g7517 ( 
.A(n_7068),
.Y(n_7517)
);

AND2x2_ASAP7_75t_L g7518 ( 
.A(n_6736),
.B(n_4156),
.Y(n_7518)
);

INVx2_ASAP7_75t_L g7519 ( 
.A(n_7005),
.Y(n_7519)
);

INVx2_ASAP7_75t_SL g7520 ( 
.A(n_6732),
.Y(n_7520)
);

XOR2x2_ASAP7_75t_SL g7521 ( 
.A(n_6746),
.B(n_4298),
.Y(n_7521)
);

INVx1_ASAP7_75t_L g7522 ( 
.A(n_7014),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7017),
.Y(n_7523)
);

OR2x2_ASAP7_75t_L g7524 ( 
.A(n_7033),
.B(n_4158),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7019),
.Y(n_7525)
);

INVx2_ASAP7_75t_SL g7526 ( 
.A(n_6732),
.Y(n_7526)
);

NAND2xp5_ASAP7_75t_SL g7527 ( 
.A(n_6991),
.B(n_4159),
.Y(n_7527)
);

INVx2_ASAP7_75t_L g7528 ( 
.A(n_7012),
.Y(n_7528)
);

NAND2xp5_ASAP7_75t_L g7529 ( 
.A(n_6584),
.B(n_4161),
.Y(n_7529)
);

INVx2_ASAP7_75t_L g7530 ( 
.A(n_7018),
.Y(n_7530)
);

NOR2xp33_ASAP7_75t_L g7531 ( 
.A(n_7027),
.B(n_4162),
.Y(n_7531)
);

INVx2_ASAP7_75t_L g7532 ( 
.A(n_7007),
.Y(n_7532)
);

INVx1_ASAP7_75t_L g7533 ( 
.A(n_7021),
.Y(n_7533)
);

OAI22xp33_ASAP7_75t_SL g7534 ( 
.A1(n_7120),
.A2(n_4306),
.B1(n_4308),
.B2(n_4299),
.Y(n_7534)
);

INVx2_ASAP7_75t_L g7535 ( 
.A(n_7025),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7026),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7028),
.Y(n_7537)
);

NOR2xp33_ASAP7_75t_L g7538 ( 
.A(n_6790),
.B(n_4166),
.Y(n_7538)
);

INVx3_ASAP7_75t_L g7539 ( 
.A(n_7068),
.Y(n_7539)
);

NAND2xp33_ASAP7_75t_L g7540 ( 
.A(n_7096),
.B(n_4168),
.Y(n_7540)
);

BUFx6f_ASAP7_75t_L g7541 ( 
.A(n_6778),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7029),
.Y(n_7542)
);

BUFx3_ASAP7_75t_L g7543 ( 
.A(n_6778),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_6755),
.Y(n_7544)
);

NAND2xp5_ASAP7_75t_SL g7545 ( 
.A(n_7113),
.B(n_4171),
.Y(n_7545)
);

CKINVDCx5p33_ASAP7_75t_R g7546 ( 
.A(n_6764),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_6724),
.Y(n_7547)
);

BUFx10_ASAP7_75t_L g7548 ( 
.A(n_6661),
.Y(n_7548)
);

AND3x2_ASAP7_75t_L g7549 ( 
.A(n_7088),
.B(n_4317),
.C(n_4309),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_6814),
.Y(n_7550)
);

INVx3_ASAP7_75t_L g7551 ( 
.A(n_7091),
.Y(n_7551)
);

INVx2_ASAP7_75t_L g7552 ( 
.A(n_7098),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7118),
.Y(n_7553)
);

INVx2_ASAP7_75t_L g7554 ( 
.A(n_7119),
.Y(n_7554)
);

INVx2_ASAP7_75t_L g7555 ( 
.A(n_6830),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_6989),
.B(n_4175),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_6928),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_6935),
.Y(n_7558)
);

BUFx2_ASAP7_75t_L g7559 ( 
.A(n_7003),
.Y(n_7559)
);

BUFx2_ASAP7_75t_L g7560 ( 
.A(n_6768),
.Y(n_7560)
);

NAND3xp33_ASAP7_75t_L g7561 ( 
.A(n_6902),
.B(n_4178),
.C(n_4177),
.Y(n_7561)
);

NOR2xp33_ASAP7_75t_L g7562 ( 
.A(n_6815),
.B(n_4179),
.Y(n_7562)
);

AND2x2_ASAP7_75t_L g7563 ( 
.A(n_7011),
.B(n_4180),
.Y(n_7563)
);

INVx3_ASAP7_75t_L g7564 ( 
.A(n_7091),
.Y(n_7564)
);

NAND2xp5_ASAP7_75t_SL g7565 ( 
.A(n_7113),
.B(n_4184),
.Y(n_7565)
);

INVx1_ASAP7_75t_L g7566 ( 
.A(n_6939),
.Y(n_7566)
);

INVx2_ASAP7_75t_L g7567 ( 
.A(n_7095),
.Y(n_7567)
);

AOI21x1_ASAP7_75t_L g7568 ( 
.A1(n_7128),
.A2(n_4330),
.B(n_4324),
.Y(n_7568)
);

AOI22xp5_ASAP7_75t_L g7569 ( 
.A1(n_7065),
.A2(n_7122),
.B1(n_7041),
.B2(n_6678),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_6957),
.Y(n_7570)
);

NAND2xp5_ASAP7_75t_L g7571 ( 
.A(n_6620),
.B(n_6684),
.Y(n_7571)
);

NAND2xp5_ASAP7_75t_SL g7572 ( 
.A(n_7097),
.B(n_4186),
.Y(n_7572)
);

BUFx6f_ASAP7_75t_L g7573 ( 
.A(n_6793),
.Y(n_7573)
);

AOI22xp33_ASAP7_75t_L g7574 ( 
.A1(n_7116),
.A2(n_4332),
.B1(n_4335),
.B2(n_4331),
.Y(n_7574)
);

BUFx2_ASAP7_75t_L g7575 ( 
.A(n_6816),
.Y(n_7575)
);

CKINVDCx11_ASAP7_75t_R g7576 ( 
.A(n_6799),
.Y(n_7576)
);

BUFx10_ASAP7_75t_L g7577 ( 
.A(n_6671),
.Y(n_7577)
);

INVx2_ASAP7_75t_SL g7578 ( 
.A(n_6793),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_6962),
.Y(n_7579)
);

INVx2_ASAP7_75t_L g7580 ( 
.A(n_7094),
.Y(n_7580)
);

NAND2xp5_ASAP7_75t_L g7581 ( 
.A(n_6687),
.B(n_4188),
.Y(n_7581)
);

AOI22xp5_ASAP7_75t_L g7582 ( 
.A1(n_6690),
.A2(n_4196),
.B1(n_4199),
.B2(n_4194),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_6971),
.Y(n_7583)
);

NOR2xp33_ASAP7_75t_L g7584 ( 
.A(n_6640),
.B(n_4201),
.Y(n_7584)
);

NAND2xp5_ASAP7_75t_L g7585 ( 
.A(n_6696),
.B(n_4204),
.Y(n_7585)
);

INVxp33_ASAP7_75t_L g7586 ( 
.A(n_7013),
.Y(n_7586)
);

BUFx3_ASAP7_75t_L g7587 ( 
.A(n_6841),
.Y(n_7587)
);

AO22x2_ASAP7_75t_L g7588 ( 
.A1(n_7124),
.A2(n_4347),
.B1(n_4348),
.B2(n_4339),
.Y(n_7588)
);

INVx2_ASAP7_75t_L g7589 ( 
.A(n_7006),
.Y(n_7589)
);

NOR2xp33_ASAP7_75t_L g7590 ( 
.A(n_6765),
.B(n_4208),
.Y(n_7590)
);

INVx2_ASAP7_75t_L g7591 ( 
.A(n_6996),
.Y(n_7591)
);

BUFx3_ASAP7_75t_L g7592 ( 
.A(n_6841),
.Y(n_7592)
);

NOR2xp33_ASAP7_75t_R g7593 ( 
.A(n_6613),
.B(n_6913),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_6974),
.Y(n_7594)
);

INVx2_ASAP7_75t_L g7595 ( 
.A(n_7092),
.Y(n_7595)
);

OR2x6_ASAP7_75t_L g7596 ( 
.A(n_6585),
.B(n_4349),
.Y(n_7596)
);

INVx2_ASAP7_75t_L g7597 ( 
.A(n_6753),
.Y(n_7597)
);

INVx2_ASAP7_75t_L g7598 ( 
.A(n_7052),
.Y(n_7598)
);

CKINVDCx5p33_ASAP7_75t_R g7599 ( 
.A(n_6777),
.Y(n_7599)
);

AND2x2_ASAP7_75t_L g7600 ( 
.A(n_7067),
.B(n_4209),
.Y(n_7600)
);

INVx2_ASAP7_75t_SL g7601 ( 
.A(n_6860),
.Y(n_7601)
);

NAND2xp5_ASAP7_75t_L g7602 ( 
.A(n_7102),
.B(n_4211),
.Y(n_7602)
);

AND2x2_ASAP7_75t_L g7603 ( 
.A(n_7105),
.B(n_4214),
.Y(n_7603)
);

INVx2_ASAP7_75t_L g7604 ( 
.A(n_7055),
.Y(n_7604)
);

BUFx6f_ASAP7_75t_L g7605 ( 
.A(n_6860),
.Y(n_7605)
);

INVx2_ASAP7_75t_L g7606 ( 
.A(n_7061),
.Y(n_7606)
);

INVx3_ASAP7_75t_L g7607 ( 
.A(n_6865),
.Y(n_7607)
);

CKINVDCx5p33_ASAP7_75t_R g7608 ( 
.A(n_6780),
.Y(n_7608)
);

HB1xp67_ASAP7_75t_L g7609 ( 
.A(n_7107),
.Y(n_7609)
);

INVx2_ASAP7_75t_L g7610 ( 
.A(n_7062),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_7064),
.Y(n_7611)
);

AOI22xp33_ASAP7_75t_L g7612 ( 
.A1(n_7121),
.A2(n_4357),
.B1(n_4361),
.B2(n_4354),
.Y(n_7612)
);

OR2x2_ASAP7_75t_L g7613 ( 
.A(n_6857),
.B(n_4219),
.Y(n_7613)
);

OAI22xp33_ASAP7_75t_L g7614 ( 
.A1(n_6981),
.A2(n_4225),
.B1(n_4227),
.B2(n_4222),
.Y(n_7614)
);

INVx2_ASAP7_75t_L g7615 ( 
.A(n_7110),
.Y(n_7615)
);

NAND2xp5_ASAP7_75t_SL g7616 ( 
.A(n_7112),
.B(n_4229),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6982),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_6998),
.Y(n_7618)
);

NOR2xp33_ASAP7_75t_L g7619 ( 
.A(n_6782),
.B(n_4230),
.Y(n_7619)
);

AO21x2_ASAP7_75t_L g7620 ( 
.A1(n_7016),
.A2(n_4368),
.B(n_4362),
.Y(n_7620)
);

AOI22xp33_ASAP7_75t_L g7621 ( 
.A1(n_6983),
.A2(n_4378),
.B1(n_4379),
.B2(n_4369),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7054),
.Y(n_7622)
);

INVx3_ASAP7_75t_L g7623 ( 
.A(n_6872),
.Y(n_7623)
);

NAND2xp5_ASAP7_75t_SL g7624 ( 
.A(n_6758),
.B(n_4232),
.Y(n_7624)
);

INVx2_ASAP7_75t_L g7625 ( 
.A(n_6895),
.Y(n_7625)
);

BUFx6f_ASAP7_75t_L g7626 ( 
.A(n_6668),
.Y(n_7626)
);

OR2x2_ASAP7_75t_L g7627 ( 
.A(n_6859),
.B(n_4233),
.Y(n_7627)
);

BUFx6f_ASAP7_75t_L g7628 ( 
.A(n_6927),
.Y(n_7628)
);

BUFx2_ASAP7_75t_L g7629 ( 
.A(n_6787),
.Y(n_7629)
);

INVx2_ASAP7_75t_L g7630 ( 
.A(n_6912),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_6945),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_6884),
.Y(n_7632)
);

INVx1_ASAP7_75t_SL g7633 ( 
.A(n_6788),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_6904),
.Y(n_7634)
);

AND3x2_ASAP7_75t_L g7635 ( 
.A(n_6851),
.B(n_4381),
.C(n_4380),
.Y(n_7635)
);

INVx2_ASAP7_75t_L g7636 ( 
.A(n_6918),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_6936),
.Y(n_7637)
);

INVx3_ASAP7_75t_L g7638 ( 
.A(n_6948),
.Y(n_7638)
);

INVx3_ASAP7_75t_L g7639 ( 
.A(n_6959),
.Y(n_7639)
);

INVx5_ASAP7_75t_L g7640 ( 
.A(n_7100),
.Y(n_7640)
);

INVx2_ASAP7_75t_L g7641 ( 
.A(n_7042),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_L g7642 ( 
.A(n_7096),
.B(n_4238),
.Y(n_7642)
);

INVx4_ASAP7_75t_L g7643 ( 
.A(n_6785),
.Y(n_7643)
);

BUFx2_ASAP7_75t_L g7644 ( 
.A(n_6864),
.Y(n_7644)
);

INVx3_ASAP7_75t_L g7645 ( 
.A(n_7090),
.Y(n_7645)
);

INVx4_ASAP7_75t_L g7646 ( 
.A(n_6593),
.Y(n_7646)
);

INVx2_ASAP7_75t_SL g7647 ( 
.A(n_7037),
.Y(n_7647)
);

INVx1_ASAP7_75t_SL g7648 ( 
.A(n_6867),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_6932),
.Y(n_7649)
);

AND2x2_ASAP7_75t_L g7650 ( 
.A(n_6728),
.B(n_4240),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_6646),
.Y(n_7651)
);

INVx2_ASAP7_75t_L g7652 ( 
.A(n_6672),
.Y(n_7652)
);

INVx2_ASAP7_75t_L g7653 ( 
.A(n_6723),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_6738),
.Y(n_7654)
);

BUFx3_ASAP7_75t_L g7655 ( 
.A(n_6604),
.Y(n_7655)
);

BUFx2_ASAP7_75t_L g7656 ( 
.A(n_6882),
.Y(n_7656)
);

INVx1_ASAP7_75t_L g7657 ( 
.A(n_6771),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_6807),
.Y(n_7658)
);

INVx2_ASAP7_75t_L g7659 ( 
.A(n_6825),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_6847),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_6890),
.Y(n_7661)
);

INVx2_ASAP7_75t_L g7662 ( 
.A(n_7096),
.Y(n_7662)
);

INVx3_ASAP7_75t_L g7663 ( 
.A(n_6909),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7104),
.Y(n_7664)
);

NAND2xp5_ASAP7_75t_L g7665 ( 
.A(n_7104),
.B(n_4241),
.Y(n_7665)
);

BUFx3_ASAP7_75t_L g7666 ( 
.A(n_6635),
.Y(n_7666)
);

NAND3xp33_ASAP7_75t_L g7667 ( 
.A(n_7074),
.B(n_4245),
.C(n_4244),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7104),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_6900),
.Y(n_7669)
);

INVx4_ASAP7_75t_L g7670 ( 
.A(n_6675),
.Y(n_7670)
);

INVx4_ASAP7_75t_L g7671 ( 
.A(n_6682),
.Y(n_7671)
);

INVx2_ASAP7_75t_L g7672 ( 
.A(n_7076),
.Y(n_7672)
);

NAND2xp5_ASAP7_75t_L g7673 ( 
.A(n_6645),
.B(n_6673),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_6921),
.B(n_4246),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7020),
.Y(n_7675)
);

INVx2_ASAP7_75t_L g7676 ( 
.A(n_6947),
.Y(n_7676)
);

NAND2xp5_ASAP7_75t_L g7677 ( 
.A(n_7022),
.B(n_4248),
.Y(n_7677)
);

NAND2xp5_ASAP7_75t_L g7678 ( 
.A(n_7114),
.B(n_4252),
.Y(n_7678)
);

INVx2_ASAP7_75t_L g7679 ( 
.A(n_6910),
.Y(n_7679)
);

INVx2_ASAP7_75t_L g7680 ( 
.A(n_6894),
.Y(n_7680)
);

INVx2_ASAP7_75t_L g7681 ( 
.A(n_6899),
.Y(n_7681)
);

INVx4_ASAP7_75t_L g7682 ( 
.A(n_6683),
.Y(n_7682)
);

INVx2_ASAP7_75t_L g7683 ( 
.A(n_7109),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7132),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7148),
.Y(n_7685)
);

INVx1_ASAP7_75t_L g7686 ( 
.A(n_7161),
.Y(n_7686)
);

INVx1_ASAP7_75t_L g7687 ( 
.A(n_7180),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7188),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_7193),
.Y(n_7689)
);

NOR2xp67_ASAP7_75t_L g7690 ( 
.A(n_7235),
.B(n_6697),
.Y(n_7690)
);

HB1xp67_ASAP7_75t_L g7691 ( 
.A(n_7208),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_7194),
.Y(n_7692)
);

AND2x2_ASAP7_75t_SL g7693 ( 
.A(n_7270),
.B(n_6601),
.Y(n_7693)
);

NAND2xp5_ASAP7_75t_L g7694 ( 
.A(n_7304),
.B(n_6660),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7552),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7196),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7199),
.Y(n_7697)
);

INVx2_ASAP7_75t_L g7698 ( 
.A(n_7553),
.Y(n_7698)
);

CKINVDCx20_ASAP7_75t_R g7699 ( 
.A(n_7179),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7201),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_7202),
.Y(n_7701)
);

INVx1_ASAP7_75t_L g7702 ( 
.A(n_7204),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7207),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7210),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7213),
.Y(n_7705)
);

AND2x4_ASAP7_75t_L g7706 ( 
.A(n_7170),
.B(n_6641),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7217),
.Y(n_7707)
);

CKINVDCx20_ASAP7_75t_R g7708 ( 
.A(n_7189),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_7223),
.Y(n_7709)
);

INVxp33_ASAP7_75t_L g7710 ( 
.A(n_7473),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7226),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7227),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7228),
.Y(n_7713)
);

INVx4_ASAP7_75t_L g7714 ( 
.A(n_7185),
.Y(n_7714)
);

AND2x2_ASAP7_75t_L g7715 ( 
.A(n_7215),
.B(n_7440),
.Y(n_7715)
);

AND2x4_ASAP7_75t_L g7716 ( 
.A(n_7175),
.B(n_6709),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7237),
.Y(n_7717)
);

INVx1_ASAP7_75t_L g7718 ( 
.A(n_7250),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_7251),
.Y(n_7719)
);

INVx2_ASAP7_75t_SL g7720 ( 
.A(n_7429),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_7255),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_7256),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_7323),
.B(n_7043),
.Y(n_7723)
);

NOR2xp33_ASAP7_75t_L g7724 ( 
.A(n_7165),
.B(n_7000),
.Y(n_7724)
);

NOR2xp33_ASAP7_75t_SL g7725 ( 
.A(n_7146),
.B(n_6698),
.Y(n_7725)
);

AND2x4_ASAP7_75t_L g7726 ( 
.A(n_7218),
.B(n_6702),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_7271),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7272),
.Y(n_7728)
);

AND2x2_ASAP7_75t_L g7729 ( 
.A(n_7414),
.B(n_6705),
.Y(n_7729)
);

INVx1_ASAP7_75t_L g7730 ( 
.A(n_7283),
.Y(n_7730)
);

NOR2xp33_ASAP7_75t_L g7731 ( 
.A(n_7156),
.B(n_6707),
.Y(n_7731)
);

CKINVDCx20_ASAP7_75t_R g7732 ( 
.A(n_7576),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7287),
.Y(n_7733)
);

NOR2xp33_ASAP7_75t_SL g7734 ( 
.A(n_7154),
.B(n_6704),
.Y(n_7734)
);

INVx1_ASAP7_75t_L g7735 ( 
.A(n_7298),
.Y(n_7735)
);

INVx1_ASAP7_75t_SL g7736 ( 
.A(n_7241),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_7303),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7305),
.Y(n_7738)
);

AND2x2_ASAP7_75t_L g7739 ( 
.A(n_7220),
.B(n_7047),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_7311),
.Y(n_7740)
);

CKINVDCx20_ASAP7_75t_R g7741 ( 
.A(n_7249),
.Y(n_7741)
);

BUFx6f_ASAP7_75t_L g7742 ( 
.A(n_7177),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_7314),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7320),
.Y(n_7744)
);

AND2x4_ASAP7_75t_L g7745 ( 
.A(n_7236),
.B(n_7655),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_SL g7746 ( 
.A(n_7309),
.B(n_6834),
.Y(n_7746)
);

INVx2_ASAP7_75t_L g7747 ( 
.A(n_7554),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7328),
.Y(n_7748)
);

NOR2x1p5_ASAP7_75t_L g7749 ( 
.A(n_7258),
.B(n_6956),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7341),
.Y(n_7750)
);

INVxp33_ASAP7_75t_L g7751 ( 
.A(n_7379),
.Y(n_7751)
);

BUFx3_ASAP7_75t_L g7752 ( 
.A(n_7185),
.Y(n_7752)
);

INVx1_ASAP7_75t_L g7753 ( 
.A(n_7342),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_7348),
.Y(n_7754)
);

NOR2xp33_ASAP7_75t_L g7755 ( 
.A(n_7150),
.B(n_7377),
.Y(n_7755)
);

INVx1_ASAP7_75t_L g7756 ( 
.A(n_7350),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7352),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_7354),
.Y(n_7758)
);

AOI21xp5_ASAP7_75t_L g7759 ( 
.A1(n_7673),
.A2(n_4393),
.B(n_4386),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_7355),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7357),
.Y(n_7761)
);

INVx1_ASAP7_75t_L g7762 ( 
.A(n_7359),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7219),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7224),
.Y(n_7764)
);

INVx2_ASAP7_75t_L g7765 ( 
.A(n_7231),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7233),
.Y(n_7766)
);

NAND2x1p5_ASAP7_75t_L g7767 ( 
.A(n_7245),
.B(n_6644),
.Y(n_7767)
);

AND2x2_ASAP7_75t_L g7768 ( 
.A(n_7240),
.B(n_6915),
.Y(n_7768)
);

OR2x2_ASAP7_75t_L g7769 ( 
.A(n_7678),
.B(n_4256),
.Y(n_7769)
);

OAI21xp5_ASAP7_75t_L g7770 ( 
.A1(n_7571),
.A2(n_4399),
.B(n_4396),
.Y(n_7770)
);

CKINVDCx5p33_ASAP7_75t_R g7771 ( 
.A(n_7297),
.Y(n_7771)
);

INVxp33_ASAP7_75t_L g7772 ( 
.A(n_7153),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7239),
.Y(n_7773)
);

INVx2_ASAP7_75t_L g7774 ( 
.A(n_7243),
.Y(n_7774)
);

NOR2xp67_ASAP7_75t_L g7775 ( 
.A(n_7319),
.B(n_3383),
.Y(n_7775)
);

CKINVDCx20_ASAP7_75t_R g7776 ( 
.A(n_7331),
.Y(n_7776)
);

INVx1_ASAP7_75t_L g7777 ( 
.A(n_7244),
.Y(n_7777)
);

CKINVDCx20_ASAP7_75t_R g7778 ( 
.A(n_7336),
.Y(n_7778)
);

CKINVDCx20_ASAP7_75t_R g7779 ( 
.A(n_7398),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7247),
.Y(n_7780)
);

AOI21x1_ASAP7_75t_L g7781 ( 
.A1(n_7547),
.A2(n_4404),
.B(n_4403),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7252),
.Y(n_7782)
);

INVx2_ASAP7_75t_L g7783 ( 
.A(n_7257),
.Y(n_7783)
);

INVx2_ASAP7_75t_L g7784 ( 
.A(n_7261),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7269),
.Y(n_7785)
);

INVx2_ASAP7_75t_L g7786 ( 
.A(n_7289),
.Y(n_7786)
);

XOR2xp5_ASAP7_75t_L g7787 ( 
.A(n_7442),
.B(n_6621),
.Y(n_7787)
);

INVx2_ASAP7_75t_L g7788 ( 
.A(n_7296),
.Y(n_7788)
);

INVx1_ASAP7_75t_L g7789 ( 
.A(n_7312),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7316),
.Y(n_7790)
);

OR2x2_ASAP7_75t_L g7791 ( 
.A(n_7200),
.B(n_4257),
.Y(n_7791)
);

INVx2_ASAP7_75t_L g7792 ( 
.A(n_7317),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_7326),
.Y(n_7793)
);

NOR2xp33_ASAP7_75t_L g7794 ( 
.A(n_7531),
.B(n_6629),
.Y(n_7794)
);

NOR2xp33_ASAP7_75t_L g7795 ( 
.A(n_7276),
.B(n_6801),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7327),
.Y(n_7796)
);

CKINVDCx5p33_ASAP7_75t_R g7797 ( 
.A(n_7406),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7330),
.Y(n_7798)
);

NOR2xp33_ASAP7_75t_L g7799 ( 
.A(n_7361),
.B(n_6804),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_7332),
.Y(n_7800)
);

INVx1_ASAP7_75t_L g7801 ( 
.A(n_7333),
.Y(n_7801)
);

CKINVDCx5p33_ASAP7_75t_R g7802 ( 
.A(n_7426),
.Y(n_7802)
);

INVx1_ASAP7_75t_L g7803 ( 
.A(n_7338),
.Y(n_7803)
);

NAND2xp5_ASAP7_75t_L g7804 ( 
.A(n_7159),
.B(n_7164),
.Y(n_7804)
);

INVx1_ASAP7_75t_L g7805 ( 
.A(n_7339),
.Y(n_7805)
);

INVxp67_ASAP7_75t_L g7806 ( 
.A(n_7402),
.Y(n_7806)
);

INVx2_ASAP7_75t_L g7807 ( 
.A(n_7344),
.Y(n_7807)
);

INVx1_ASAP7_75t_L g7808 ( 
.A(n_7356),
.Y(n_7808)
);

NAND2xp5_ASAP7_75t_SL g7809 ( 
.A(n_7569),
.B(n_4258),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7365),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_7366),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7375),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7378),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_7389),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7393),
.Y(n_7815)
);

INVxp67_ASAP7_75t_SL g7816 ( 
.A(n_7609),
.Y(n_7816)
);

NOR2xp33_ASAP7_75t_L g7817 ( 
.A(n_7364),
.B(n_4259),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7399),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_7400),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7408),
.Y(n_7820)
);

INVx1_ASAP7_75t_L g7821 ( 
.A(n_7409),
.Y(n_7821)
);

AND2x2_ASAP7_75t_L g7822 ( 
.A(n_7315),
.B(n_4261),
.Y(n_7822)
);

NOR2xp33_ASAP7_75t_SL g7823 ( 
.A(n_7546),
.B(n_4262),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_7410),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_7419),
.Y(n_7825)
);

INVx1_ASAP7_75t_L g7826 ( 
.A(n_7423),
.Y(n_7826)
);

INVx2_ASAP7_75t_L g7827 ( 
.A(n_7532),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_7427),
.Y(n_7828)
);

AND2x2_ASAP7_75t_L g7829 ( 
.A(n_7556),
.B(n_4266),
.Y(n_7829)
);

INVx2_ASAP7_75t_L g7830 ( 
.A(n_7595),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7432),
.Y(n_7831)
);

NOR2xp33_ASAP7_75t_L g7832 ( 
.A(n_7184),
.B(n_4267),
.Y(n_7832)
);

NOR2xp33_ASAP7_75t_L g7833 ( 
.A(n_7345),
.B(n_7586),
.Y(n_7833)
);

INVxp67_ASAP7_75t_SL g7834 ( 
.A(n_7178),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7441),
.Y(n_7835)
);

INVx1_ASAP7_75t_L g7836 ( 
.A(n_7444),
.Y(n_7836)
);

INVx1_ASAP7_75t_SL g7837 ( 
.A(n_7293),
.Y(n_7837)
);

CKINVDCx11_ASAP7_75t_R g7838 ( 
.A(n_7491),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7445),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7450),
.Y(n_7840)
);

INVx2_ASAP7_75t_L g7841 ( 
.A(n_7130),
.Y(n_7841)
);

INVx2_ASAP7_75t_L g7842 ( 
.A(n_7133),
.Y(n_7842)
);

INVx2_ASAP7_75t_L g7843 ( 
.A(n_7136),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_7451),
.Y(n_7844)
);

INVxp67_ASAP7_75t_SL g7845 ( 
.A(n_7171),
.Y(n_7845)
);

INVx1_ASAP7_75t_L g7846 ( 
.A(n_7458),
.Y(n_7846)
);

XOR2xp5_ASAP7_75t_L g7847 ( 
.A(n_7599),
.B(n_3384),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7463),
.Y(n_7848)
);

AND2x2_ASAP7_75t_L g7849 ( 
.A(n_7563),
.B(n_4268),
.Y(n_7849)
);

NOR2xp33_ASAP7_75t_L g7850 ( 
.A(n_7308),
.B(n_4270),
.Y(n_7850)
);

NOR2xp33_ASAP7_75t_L g7851 ( 
.A(n_7313),
.B(n_4271),
.Y(n_7851)
);

INVx2_ASAP7_75t_L g7852 ( 
.A(n_7137),
.Y(n_7852)
);

AND2x2_ASAP7_75t_L g7853 ( 
.A(n_7438),
.B(n_4274),
.Y(n_7853)
);

INVx2_ASAP7_75t_L g7854 ( 
.A(n_7138),
.Y(n_7854)
);

NOR2xp33_ASAP7_75t_SL g7855 ( 
.A(n_7608),
.B(n_7670),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7467),
.Y(n_7856)
);

INVxp67_ASAP7_75t_SL g7857 ( 
.A(n_7216),
.Y(n_7857)
);

NOR2xp33_ASAP7_75t_L g7858 ( 
.A(n_7557),
.B(n_4277),
.Y(n_7858)
);

CKINVDCx5p33_ASAP7_75t_R g7859 ( 
.A(n_7151),
.Y(n_7859)
);

INVx1_ASAP7_75t_L g7860 ( 
.A(n_7468),
.Y(n_7860)
);

NAND2xp5_ASAP7_75t_L g7861 ( 
.A(n_7558),
.B(n_4279),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_7476),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_7480),
.Y(n_7863)
);

NOR2xp33_ASAP7_75t_L g7864 ( 
.A(n_7566),
.B(n_4280),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7482),
.Y(n_7865)
);

BUFx3_ASAP7_75t_L g7866 ( 
.A(n_7275),
.Y(n_7866)
);

XNOR2xp5_ASAP7_75t_L g7867 ( 
.A(n_7349),
.B(n_7292),
.Y(n_7867)
);

INVx1_ASAP7_75t_L g7868 ( 
.A(n_7484),
.Y(n_7868)
);

AND2x2_ASAP7_75t_L g7869 ( 
.A(n_7343),
.B(n_4281),
.Y(n_7869)
);

XOR2xp5_ASAP7_75t_L g7870 ( 
.A(n_7629),
.B(n_3387),
.Y(n_7870)
);

INVx4_ASAP7_75t_L g7871 ( 
.A(n_7275),
.Y(n_7871)
);

INVxp67_ASAP7_75t_SL g7872 ( 
.A(n_7234),
.Y(n_7872)
);

NAND2xp5_ASAP7_75t_L g7873 ( 
.A(n_7570),
.B(n_4282),
.Y(n_7873)
);

CKINVDCx5p33_ASAP7_75t_R g7874 ( 
.A(n_7174),
.Y(n_7874)
);

AND2x2_ASAP7_75t_SL g7875 ( 
.A(n_7281),
.B(n_4407),
.Y(n_7875)
);

OR2x2_ASAP7_75t_L g7876 ( 
.A(n_7676),
.B(n_4283),
.Y(n_7876)
);

CKINVDCx20_ASAP7_75t_R g7877 ( 
.A(n_7407),
.Y(n_7877)
);

INVx2_ASAP7_75t_L g7878 ( 
.A(n_7139),
.Y(n_7878)
);

CKINVDCx20_ASAP7_75t_R g7879 ( 
.A(n_7407),
.Y(n_7879)
);

AND2x4_ASAP7_75t_L g7880 ( 
.A(n_7385),
.B(n_7424),
.Y(n_7880)
);

INVxp33_ASAP7_75t_L g7881 ( 
.A(n_7263),
.Y(n_7881)
);

NOR2xp33_ASAP7_75t_L g7882 ( 
.A(n_7579),
.B(n_4284),
.Y(n_7882)
);

NOR2xp67_ASAP7_75t_L g7883 ( 
.A(n_7221),
.B(n_3391),
.Y(n_7883)
);

BUFx3_ASAP7_75t_L g7884 ( 
.A(n_7268),
.Y(n_7884)
);

NOR2xp33_ASAP7_75t_L g7885 ( 
.A(n_7583),
.B(n_4286),
.Y(n_7885)
);

CKINVDCx20_ASAP7_75t_R g7886 ( 
.A(n_7593),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_7489),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_7495),
.Y(n_7888)
);

NAND2xp5_ASAP7_75t_L g7889 ( 
.A(n_7209),
.B(n_4287),
.Y(n_7889)
);

AND2x2_ASAP7_75t_L g7890 ( 
.A(n_7353),
.B(n_7363),
.Y(n_7890)
);

NAND2x1p5_ASAP7_75t_L g7891 ( 
.A(n_7643),
.B(n_7360),
.Y(n_7891)
);

INVxp67_ASAP7_75t_L g7892 ( 
.A(n_7259),
.Y(n_7892)
);

INVx1_ASAP7_75t_L g7893 ( 
.A(n_7499),
.Y(n_7893)
);

AND2x2_ASAP7_75t_L g7894 ( 
.A(n_7518),
.B(n_4288),
.Y(n_7894)
);

NOR2xp33_ASAP7_75t_L g7895 ( 
.A(n_7412),
.B(n_4293),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_7500),
.Y(n_7896)
);

INVx1_ASAP7_75t_L g7897 ( 
.A(n_7503),
.Y(n_7897)
);

AND2x4_ASAP7_75t_L g7898 ( 
.A(n_7454),
.B(n_4408),
.Y(n_7898)
);

OAI21xp5_ASAP7_75t_L g7899 ( 
.A1(n_7615),
.A2(n_4416),
.B(n_4415),
.Y(n_7899)
);

INVx2_ASAP7_75t_L g7900 ( 
.A(n_7140),
.Y(n_7900)
);

AND2x2_ASAP7_75t_L g7901 ( 
.A(n_7675),
.B(n_4294),
.Y(n_7901)
);

CKINVDCx5p33_ASAP7_75t_R g7902 ( 
.A(n_7246),
.Y(n_7902)
);

AND2x2_ASAP7_75t_L g7903 ( 
.A(n_7483),
.B(n_4295),
.Y(n_7903)
);

NAND2xp33_ASAP7_75t_R g7904 ( 
.A(n_7644),
.B(n_3392),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7142),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7147),
.Y(n_7906)
);

INVx1_ASAP7_75t_L g7907 ( 
.A(n_7149),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7163),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_7182),
.Y(n_7909)
);

BUFx6f_ASAP7_75t_L g7910 ( 
.A(n_7177),
.Y(n_7910)
);

INVx2_ASAP7_75t_L g7911 ( 
.A(n_7183),
.Y(n_7911)
);

INVx1_ASAP7_75t_L g7912 ( 
.A(n_7186),
.Y(n_7912)
);

INVx2_ASAP7_75t_L g7913 ( 
.A(n_7203),
.Y(n_7913)
);

INVx1_ASAP7_75t_L g7914 ( 
.A(n_7206),
.Y(n_7914)
);

AND2x2_ASAP7_75t_L g7915 ( 
.A(n_7600),
.B(n_4300),
.Y(n_7915)
);

NOR2xp33_ASAP7_75t_L g7916 ( 
.A(n_7325),
.B(n_4301),
.Y(n_7916)
);

AND2x2_ASAP7_75t_L g7917 ( 
.A(n_7603),
.B(n_4302),
.Y(n_7917)
);

NOR2xp33_ASAP7_75t_L g7918 ( 
.A(n_7448),
.B(n_4303),
.Y(n_7918)
);

OAI21xp5_ASAP7_75t_L g7919 ( 
.A1(n_7510),
.A2(n_4427),
.B(n_4418),
.Y(n_7919)
);

CKINVDCx20_ASAP7_75t_R g7920 ( 
.A(n_7656),
.Y(n_7920)
);

INVx1_ASAP7_75t_L g7921 ( 
.A(n_7211),
.Y(n_7921)
);

INVxp67_ASAP7_75t_L g7922 ( 
.A(n_7279),
.Y(n_7922)
);

CKINVDCx5p33_ASAP7_75t_R g7923 ( 
.A(n_7322),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7212),
.Y(n_7924)
);

INVx1_ASAP7_75t_L g7925 ( 
.A(n_7380),
.Y(n_7925)
);

AND2x2_ASAP7_75t_L g7926 ( 
.A(n_7436),
.B(n_4304),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7381),
.Y(n_7927)
);

INVx1_ASAP7_75t_L g7928 ( 
.A(n_7384),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_7387),
.Y(n_7929)
);

NAND2xp33_ASAP7_75t_R g7930 ( 
.A(n_7470),
.B(n_3393),
.Y(n_7930)
);

AND2x4_ASAP7_75t_L g7931 ( 
.A(n_7371),
.B(n_4432),
.Y(n_7931)
);

AND2x2_ASAP7_75t_L g7932 ( 
.A(n_7590),
.B(n_4310),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_7388),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_7392),
.Y(n_7934)
);

NOR2xp33_ASAP7_75t_L g7935 ( 
.A(n_7619),
.B(n_4312),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_7395),
.Y(n_7936)
);

CKINVDCx16_ASAP7_75t_R g7937 ( 
.A(n_7152),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7413),
.Y(n_7938)
);

INVx1_ASAP7_75t_SL g7939 ( 
.A(n_7559),
.Y(n_7939)
);

XOR2xp5_ASAP7_75t_L g7940 ( 
.A(n_7479),
.B(n_3394),
.Y(n_7940)
);

AND2x2_ASAP7_75t_L g7941 ( 
.A(n_7254),
.B(n_4313),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_7416),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7418),
.Y(n_7943)
);

INVxp33_ASAP7_75t_L g7944 ( 
.A(n_7397),
.Y(n_7944)
);

INVx1_ASAP7_75t_L g7945 ( 
.A(n_7425),
.Y(n_7945)
);

INVx1_ASAP7_75t_L g7946 ( 
.A(n_7428),
.Y(n_7946)
);

XOR2x2_ASAP7_75t_L g7947 ( 
.A(n_7521),
.B(n_6),
.Y(n_7947)
);

INVx1_ASAP7_75t_L g7948 ( 
.A(n_7435),
.Y(n_7948)
);

XNOR2xp5_ASAP7_75t_L g7949 ( 
.A(n_7633),
.B(n_3395),
.Y(n_7949)
);

BUFx6f_ASAP7_75t_L g7950 ( 
.A(n_7288),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7439),
.Y(n_7951)
);

INVx2_ASAP7_75t_L g7952 ( 
.A(n_7443),
.Y(n_7952)
);

INVx2_ASAP7_75t_L g7953 ( 
.A(n_7446),
.Y(n_7953)
);

INVx1_ASAP7_75t_L g7954 ( 
.A(n_7449),
.Y(n_7954)
);

INVx1_ASAP7_75t_L g7955 ( 
.A(n_7456),
.Y(n_7955)
);

AND2x2_ASAP7_75t_L g7956 ( 
.A(n_7260),
.B(n_4314),
.Y(n_7956)
);

INVx1_ASAP7_75t_SL g7957 ( 
.A(n_7648),
.Y(n_7957)
);

AND2x2_ASAP7_75t_L g7958 ( 
.A(n_7190),
.B(n_4316),
.Y(n_7958)
);

INVx1_ASAP7_75t_L g7959 ( 
.A(n_7457),
.Y(n_7959)
);

INVx1_ASAP7_75t_L g7960 ( 
.A(n_7469),
.Y(n_7960)
);

NAND2xp33_ASAP7_75t_R g7961 ( 
.A(n_7560),
.B(n_3397),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_7472),
.Y(n_7962)
);

OR2x2_ASAP7_75t_L g7963 ( 
.A(n_7683),
.B(n_4318),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7474),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7485),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_7498),
.Y(n_7966)
);

INVxp67_ASAP7_75t_L g7967 ( 
.A(n_7280),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_7514),
.Y(n_7968)
);

INVx1_ASAP7_75t_L g7969 ( 
.A(n_7515),
.Y(n_7969)
);

XOR2xp5_ASAP7_75t_L g7970 ( 
.A(n_7490),
.B(n_3399),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_7509),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_7522),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_7523),
.Y(n_7973)
);

INVx2_ASAP7_75t_SL g7974 ( 
.A(n_7288),
.Y(n_7974)
);

XOR2xp5_ASAP7_75t_L g7975 ( 
.A(n_7666),
.B(n_3400),
.Y(n_7975)
);

AND2x2_ASAP7_75t_L g7976 ( 
.A(n_7650),
.B(n_4319),
.Y(n_7976)
);

CKINVDCx20_ASAP7_75t_R g7977 ( 
.A(n_7144),
.Y(n_7977)
);

AND2x2_ASAP7_75t_L g7978 ( 
.A(n_7135),
.B(n_7386),
.Y(n_7978)
);

INVx2_ASAP7_75t_L g7979 ( 
.A(n_7567),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7525),
.Y(n_7980)
);

INVx1_ASAP7_75t_L g7981 ( 
.A(n_7533),
.Y(n_7981)
);

AND2x6_ASAP7_75t_L g7982 ( 
.A(n_7664),
.B(n_4434),
.Y(n_7982)
);

INVx1_ASAP7_75t_L g7983 ( 
.A(n_7536),
.Y(n_7983)
);

INVx1_ASAP7_75t_L g7984 ( 
.A(n_7537),
.Y(n_7984)
);

INVx1_ASAP7_75t_L g7985 ( 
.A(n_7542),
.Y(n_7985)
);

NOR2xp33_ASAP7_75t_L g7986 ( 
.A(n_7460),
.B(n_7367),
.Y(n_7986)
);

AND2x4_ASAP7_75t_L g7987 ( 
.A(n_7229),
.B(n_4435),
.Y(n_7987)
);

CKINVDCx16_ASAP7_75t_R g7988 ( 
.A(n_7141),
.Y(n_7988)
);

INVx2_ASAP7_75t_L g7989 ( 
.A(n_7580),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7535),
.Y(n_7990)
);

NOR2xp33_ASAP7_75t_L g7991 ( 
.A(n_7461),
.B(n_4320),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7516),
.Y(n_7992)
);

AND2x2_ASAP7_75t_L g7993 ( 
.A(n_7679),
.B(n_4321),
.Y(n_7993)
);

XOR2x2_ASAP7_75t_L g7994 ( 
.A(n_7242),
.B(n_7),
.Y(n_7994)
);

INVxp33_ASAP7_75t_L g7995 ( 
.A(n_7672),
.Y(n_7995)
);

NOR2xp67_ASAP7_75t_L g7996 ( 
.A(n_7221),
.B(n_3402),
.Y(n_7996)
);

INVx1_ASAP7_75t_L g7997 ( 
.A(n_7504),
.Y(n_7997)
);

NAND2xp33_ASAP7_75t_SL g7998 ( 
.A(n_7391),
.B(n_4323),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_7519),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_7528),
.Y(n_8000)
);

INVx2_ASAP7_75t_L g8001 ( 
.A(n_7530),
.Y(n_8001)
);

NOR2xp33_ASAP7_75t_L g8002 ( 
.A(n_7334),
.B(n_4325),
.Y(n_8002)
);

NOR2xp33_ASAP7_75t_L g8003 ( 
.A(n_7346),
.B(n_4327),
.Y(n_8003)
);

INVx2_ASAP7_75t_L g8004 ( 
.A(n_7591),
.Y(n_8004)
);

AND2x4_ASAP7_75t_L g8005 ( 
.A(n_7232),
.B(n_7640),
.Y(n_8005)
);

NAND2xp5_ASAP7_75t_L g8006 ( 
.A(n_7369),
.B(n_4329),
.Y(n_8006)
);

INVx1_ASAP7_75t_L g8007 ( 
.A(n_7598),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_7604),
.Y(n_8008)
);

NOR2x1p5_ASAP7_75t_L g8009 ( 
.A(n_7626),
.B(n_4337),
.Y(n_8009)
);

NOR2xp33_ASAP7_75t_L g8010 ( 
.A(n_7455),
.B(n_7411),
.Y(n_8010)
);

CKINVDCx20_ASAP7_75t_R g8011 ( 
.A(n_7575),
.Y(n_8011)
);

NAND2x1p5_ASAP7_75t_L g8012 ( 
.A(n_7382),
.B(n_4440),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_7606),
.Y(n_8013)
);

INVx1_ASAP7_75t_L g8014 ( 
.A(n_7610),
.Y(n_8014)
);

INVx1_ASAP7_75t_L g8015 ( 
.A(n_7611),
.Y(n_8015)
);

CKINVDCx5p33_ASAP7_75t_R g8016 ( 
.A(n_7548),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7373),
.B(n_4338),
.Y(n_8017)
);

XNOR2x2_ASAP7_75t_L g8018 ( 
.A(n_7394),
.B(n_4444),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7487),
.Y(n_8019)
);

NOR2xp33_ASAP7_75t_L g8020 ( 
.A(n_7613),
.B(n_4341),
.Y(n_8020)
);

INVx2_ASAP7_75t_L g8021 ( 
.A(n_7172),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7492),
.Y(n_8022)
);

INVx2_ASAP7_75t_SL g8023 ( 
.A(n_7452),
.Y(n_8023)
);

NOR2xp33_ASAP7_75t_L g8024 ( 
.A(n_7627),
.B(n_4344),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7496),
.Y(n_8025)
);

AND2x2_ASAP7_75t_SL g8026 ( 
.A(n_7621),
.B(n_4446),
.Y(n_8026)
);

BUFx6f_ASAP7_75t_L g8027 ( 
.A(n_7452),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7663),
.B(n_4346),
.Y(n_8028)
);

CKINVDCx16_ASAP7_75t_R g8029 ( 
.A(n_7577),
.Y(n_8029)
);

NOR2xp33_ASAP7_75t_SL g8030 ( 
.A(n_7671),
.B(n_4350),
.Y(n_8030)
);

INVx1_ASAP7_75t_L g8031 ( 
.A(n_7501),
.Y(n_8031)
);

INVx2_ASAP7_75t_L g8032 ( 
.A(n_7430),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_7502),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7225),
.Y(n_8034)
);

INVx1_ASAP7_75t_SL g8035 ( 
.A(n_7324),
.Y(n_8035)
);

INVx1_ASAP7_75t_L g8036 ( 
.A(n_7466),
.Y(n_8036)
);

BUFx8_ASAP7_75t_L g8037 ( 
.A(n_7626),
.Y(n_8037)
);

AND2x2_ASAP7_75t_L g8038 ( 
.A(n_7404),
.B(n_4352),
.Y(n_8038)
);

INVx1_ASAP7_75t_L g8039 ( 
.A(n_7505),
.Y(n_8039)
);

NAND2xp5_ASAP7_75t_L g8040 ( 
.A(n_7374),
.B(n_4353),
.Y(n_8040)
);

INVx1_ASAP7_75t_L g8041 ( 
.A(n_7512),
.Y(n_8041)
);

INVx1_ASAP7_75t_L g8042 ( 
.A(n_7513),
.Y(n_8042)
);

INVx1_ASAP7_75t_SL g8043 ( 
.A(n_7337),
.Y(n_8043)
);

INVx1_ASAP7_75t_L g8044 ( 
.A(n_7544),
.Y(n_8044)
);

INVxp67_ASAP7_75t_SL g8045 ( 
.A(n_7507),
.Y(n_8045)
);

INVx1_ASAP7_75t_L g8046 ( 
.A(n_7550),
.Y(n_8046)
);

INVxp67_ASAP7_75t_L g8047 ( 
.A(n_7230),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7568),
.Y(n_8048)
);

NAND2x1p5_ASAP7_75t_L g8049 ( 
.A(n_7628),
.B(n_4453),
.Y(n_8049)
);

AND2x2_ASAP7_75t_L g8050 ( 
.A(n_7524),
.B(n_4363),
.Y(n_8050)
);

NOR2xp33_ASAP7_75t_L g8051 ( 
.A(n_7529),
.B(n_7581),
.Y(n_8051)
);

INVxp33_ASAP7_75t_SL g8052 ( 
.A(n_7674),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_7187),
.Y(n_8053)
);

INVx2_ASAP7_75t_L g8054 ( 
.A(n_7597),
.Y(n_8054)
);

AND2x4_ASAP7_75t_L g8055 ( 
.A(n_7640),
.B(n_4454),
.Y(n_8055)
);

AND2x2_ASAP7_75t_L g8056 ( 
.A(n_7306),
.B(n_4364),
.Y(n_8056)
);

AND2x2_ASAP7_75t_L g8057 ( 
.A(n_7310),
.B(n_4365),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_7198),
.Y(n_8058)
);

OAI21xp5_ASAP7_75t_L g8059 ( 
.A1(n_7403),
.A2(n_4462),
.B(n_4458),
.Y(n_8059)
);

NOR2xp33_ASAP7_75t_L g8060 ( 
.A(n_7585),
.B(n_4366),
.Y(n_8060)
);

INVxp33_ASAP7_75t_L g8061 ( 
.A(n_7465),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_L g8062 ( 
.A(n_7262),
.B(n_4367),
.Y(n_8062)
);

INVx1_ASAP7_75t_L g8063 ( 
.A(n_7264),
.Y(n_8063)
);

BUFx6f_ASAP7_75t_L g8064 ( 
.A(n_7507),
.Y(n_8064)
);

AND2x2_ASAP7_75t_L g8065 ( 
.A(n_7267),
.B(n_4372),
.Y(n_8065)
);

AND2x2_ASAP7_75t_L g8066 ( 
.A(n_7301),
.B(n_4373),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7160),
.Y(n_8067)
);

AND2x2_ASAP7_75t_L g8068 ( 
.A(n_7625),
.B(n_4374),
.Y(n_8068)
);

NOR2xp33_ASAP7_75t_L g8069 ( 
.A(n_7168),
.B(n_4375),
.Y(n_8069)
);

INVx1_ASAP7_75t_L g8070 ( 
.A(n_7651),
.Y(n_8070)
);

AOI21xp5_ASAP7_75t_L g8071 ( 
.A1(n_7618),
.A2(n_4466),
.B(n_4465),
.Y(n_8071)
);

CKINVDCx5p33_ASAP7_75t_R g8072 ( 
.A(n_7291),
.Y(n_8072)
);

INVx1_ASAP7_75t_L g8073 ( 
.A(n_7654),
.Y(n_8073)
);

INVx1_ASAP7_75t_L g8074 ( 
.A(n_7657),
.Y(n_8074)
);

INVx2_ASAP7_75t_L g8075 ( 
.A(n_7589),
.Y(n_8075)
);

INVx1_ASAP7_75t_L g8076 ( 
.A(n_7658),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7660),
.Y(n_8077)
);

CKINVDCx20_ASAP7_75t_R g8078 ( 
.A(n_7401),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7632),
.Y(n_8079)
);

INVx1_ASAP7_75t_L g8080 ( 
.A(n_7634),
.Y(n_8080)
);

AND2x2_ASAP7_75t_L g8081 ( 
.A(n_7630),
.B(n_4376),
.Y(n_8081)
);

AND2x4_ASAP7_75t_L g8082 ( 
.A(n_7646),
.B(n_4470),
.Y(n_8082)
);

BUFx8_ASAP7_75t_L g8083 ( 
.A(n_7628),
.Y(n_8083)
);

AND2x4_ASAP7_75t_L g8084 ( 
.A(n_7647),
.B(n_4471),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_7637),
.Y(n_8085)
);

AND2x2_ASAP7_75t_L g8086 ( 
.A(n_7555),
.B(n_4382),
.Y(n_8086)
);

AND2x2_ASAP7_75t_L g8087 ( 
.A(n_7584),
.B(n_4384),
.Y(n_8087)
);

NOR2xp33_ASAP7_75t_L g8088 ( 
.A(n_7661),
.B(n_4388),
.Y(n_8088)
);

NOR2xp33_ASAP7_75t_L g8089 ( 
.A(n_7421),
.B(n_4389),
.Y(n_8089)
);

XOR2xp5_ASAP7_75t_L g8090 ( 
.A(n_7561),
.B(n_3404),
.Y(n_8090)
);

NOR2xp67_ASAP7_75t_L g8091 ( 
.A(n_7291),
.B(n_3405),
.Y(n_8091)
);

HB1xp67_ASAP7_75t_L g8092 ( 
.A(n_7508),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_7652),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_7653),
.Y(n_8094)
);

XOR2xp5_ASAP7_75t_L g8095 ( 
.A(n_7667),
.B(n_3406),
.Y(n_8095)
);

INVx1_ASAP7_75t_SL g8096 ( 
.A(n_7376),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_7659),
.Y(n_8097)
);

NOR2xp33_ASAP7_75t_L g8098 ( 
.A(n_7453),
.B(n_7278),
.Y(n_8098)
);

INVx2_ASAP7_75t_L g8099 ( 
.A(n_7636),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_7641),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_L g8101 ( 
.A(n_7538),
.B(n_4390),
.Y(n_8101)
);

BUFx8_ASAP7_75t_L g8102 ( 
.A(n_7508),
.Y(n_8102)
);

INVx2_ASAP7_75t_L g8103 ( 
.A(n_7620),
.Y(n_8103)
);

INVx1_ASAP7_75t_L g8104 ( 
.A(n_7594),
.Y(n_8104)
);

XOR2xp5_ASAP7_75t_L g8105 ( 
.A(n_7494),
.B(n_3408),
.Y(n_8105)
);

NOR2xp33_ASAP7_75t_L g8106 ( 
.A(n_7286),
.B(n_4391),
.Y(n_8106)
);

NAND2xp5_ASAP7_75t_SL g8107 ( 
.A(n_7294),
.B(n_4394),
.Y(n_8107)
);

NOR2xp33_ASAP7_75t_L g8108 ( 
.A(n_7290),
.B(n_4395),
.Y(n_8108)
);

INVx1_ASAP7_75t_L g8109 ( 
.A(n_7617),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_7511),
.Y(n_8110)
);

INVxp33_ASAP7_75t_L g8111 ( 
.A(n_7541),
.Y(n_8111)
);

BUFx6f_ASAP7_75t_L g8112 ( 
.A(n_7541),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7631),
.Y(n_8113)
);

AND2x4_ASAP7_75t_L g8114 ( 
.A(n_7131),
.B(n_4477),
.Y(n_8114)
);

INVx1_ASAP7_75t_SL g8115 ( 
.A(n_7383),
.Y(n_8115)
);

INVx4_ASAP7_75t_SL g8116 ( 
.A(n_7166),
.Y(n_8116)
);

CKINVDCx5p33_ASAP7_75t_R g8117 ( 
.A(n_7145),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7588),
.Y(n_8118)
);

NAND2xp5_ASAP7_75t_L g8119 ( 
.A(n_7562),
.B(n_4398),
.Y(n_8119)
);

AND2x2_ASAP7_75t_L g8120 ( 
.A(n_7574),
.B(n_4400),
.Y(n_8120)
);

AND2x2_ASAP7_75t_L g8121 ( 
.A(n_7612),
.B(n_4402),
.Y(n_8121)
);

INVx2_ASAP7_75t_L g8122 ( 
.A(n_7669),
.Y(n_8122)
);

AND2x2_ASAP7_75t_L g8123 ( 
.A(n_7300),
.B(n_4405),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_7477),
.Y(n_8124)
);

NOR2xp33_ASAP7_75t_L g8125 ( 
.A(n_7318),
.B(n_4406),
.Y(n_8125)
);

INVxp33_ASAP7_75t_L g8126 ( 
.A(n_7573),
.Y(n_8126)
);

NOR2xp33_ASAP7_75t_L g8127 ( 
.A(n_7358),
.B(n_4409),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_7649),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_7622),
.Y(n_8129)
);

INVx1_ASAP7_75t_L g8130 ( 
.A(n_7176),
.Y(n_8130)
);

CKINVDCx20_ASAP7_75t_R g8131 ( 
.A(n_7682),
.Y(n_8131)
);

INVx1_ASAP7_75t_L g8132 ( 
.A(n_7176),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_7176),
.Y(n_8133)
);

NOR2xp33_ASAP7_75t_L g8134 ( 
.A(n_7191),
.B(n_4410),
.Y(n_8134)
);

AND2x2_ASAP7_75t_L g8135 ( 
.A(n_7155),
.B(n_4411),
.Y(n_8135)
);

INVx2_ASAP7_75t_SL g8136 ( 
.A(n_7573),
.Y(n_8136)
);

OAI21xp5_ASAP7_75t_L g8137 ( 
.A1(n_7134),
.A2(n_4485),
.B(n_4481),
.Y(n_8137)
);

CKINVDCx5p33_ASAP7_75t_R g8138 ( 
.A(n_7145),
.Y(n_8138)
);

INVx1_ASAP7_75t_L g8139 ( 
.A(n_7422),
.Y(n_8139)
);

INVx3_ASAP7_75t_L g8140 ( 
.A(n_7605),
.Y(n_8140)
);

INVx2_ASAP7_75t_L g8141 ( 
.A(n_7607),
.Y(n_8141)
);

NOR2xp33_ASAP7_75t_L g8142 ( 
.A(n_7205),
.B(n_4412),
.Y(n_8142)
);

INVxp33_ASAP7_75t_L g8143 ( 
.A(n_7605),
.Y(n_8143)
);

NOR2xp33_ASAP7_75t_L g8144 ( 
.A(n_7214),
.B(n_4414),
.Y(n_8144)
);

INVxp33_ASAP7_75t_L g8145 ( 
.A(n_7677),
.Y(n_8145)
);

AOI21x1_ASAP7_75t_L g8146 ( 
.A1(n_7434),
.A2(n_4489),
.B(n_4486),
.Y(n_8146)
);

CKINVDCx20_ASAP7_75t_R g8147 ( 
.A(n_7173),
.Y(n_8147)
);

CKINVDCx20_ASAP7_75t_R g8148 ( 
.A(n_7417),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7422),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_7422),
.Y(n_8150)
);

INVx2_ASAP7_75t_L g8151 ( 
.A(n_7623),
.Y(n_8151)
);

XOR2x2_ASAP7_75t_L g8152 ( 
.A(n_7433),
.B(n_7),
.Y(n_8152)
);

INVx1_ASAP7_75t_L g8153 ( 
.A(n_7602),
.Y(n_8153)
);

INVx1_ASAP7_75t_L g8154 ( 
.A(n_7638),
.Y(n_8154)
);

INVx1_ASAP7_75t_L g8155 ( 
.A(n_7639),
.Y(n_8155)
);

AOI21xp5_ASAP7_75t_L g8156 ( 
.A1(n_7572),
.A2(n_4501),
.B(n_4492),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7645),
.Y(n_8157)
);

INVx2_ASAP7_75t_L g8158 ( 
.A(n_7162),
.Y(n_8158)
);

XOR2xp5_ASAP7_75t_L g8159 ( 
.A(n_7680),
.B(n_3409),
.Y(n_8159)
);

INVx1_ASAP7_75t_L g8160 ( 
.A(n_7347),
.Y(n_8160)
);

INVx1_ASAP7_75t_L g8161 ( 
.A(n_7481),
.Y(n_8161)
);

BUFx6f_ASAP7_75t_SL g8162 ( 
.A(n_7464),
.Y(n_8162)
);

INVx1_ASAP7_75t_L g8163 ( 
.A(n_7299),
.Y(n_8163)
);

INVx1_ASAP7_75t_L g8164 ( 
.A(n_7362),
.Y(n_8164)
);

INVx1_ASAP7_75t_L g8165 ( 
.A(n_7420),
.Y(n_8165)
);

INVx1_ASAP7_75t_L g8166 ( 
.A(n_7169),
.Y(n_8166)
);

INVx2_ASAP7_75t_L g8167 ( 
.A(n_7192),
.Y(n_8167)
);

AND2x2_ASAP7_75t_L g8168 ( 
.A(n_7248),
.B(n_4417),
.Y(n_8168)
);

INVxp67_ASAP7_75t_SL g8169 ( 
.A(n_7471),
.Y(n_8169)
);

AND2x4_ASAP7_75t_L g8170 ( 
.A(n_7197),
.B(n_4508),
.Y(n_8170)
);

OAI21xp5_ASAP7_75t_L g8171 ( 
.A1(n_7277),
.A2(n_4514),
.B(n_4510),
.Y(n_8171)
);

XOR2xp5_ASAP7_75t_L g8172 ( 
.A(n_7681),
.B(n_3410),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7222),
.Y(n_8173)
);

NAND2xp5_ASAP7_75t_L g8174 ( 
.A(n_7390),
.B(n_7478),
.Y(n_8174)
);

NOR2xp33_ASAP7_75t_SL g8175 ( 
.A(n_7294),
.B(n_4420),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_7253),
.Y(n_8176)
);

AND2x4_ASAP7_75t_L g8177 ( 
.A(n_7265),
.B(n_7273),
.Y(n_8177)
);

INVx2_ASAP7_75t_L g8178 ( 
.A(n_7284),
.Y(n_8178)
);

INVx1_ASAP7_75t_L g8179 ( 
.A(n_7285),
.Y(n_8179)
);

INVx1_ASAP7_75t_L g8180 ( 
.A(n_7321),
.Y(n_8180)
);

CKINVDCx5p33_ASAP7_75t_R g8181 ( 
.A(n_7195),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7335),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7462),
.Y(n_8183)
);

XOR2xp5_ASAP7_75t_L g8184 ( 
.A(n_7351),
.B(n_3411),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7517),
.Y(n_8185)
);

INVxp67_ASAP7_75t_SL g8186 ( 
.A(n_7543),
.Y(n_8186)
);

INVx1_ASAP7_75t_L g8187 ( 
.A(n_7539),
.Y(n_8187)
);

XOR2xp5_ASAP7_75t_L g8188 ( 
.A(n_7582),
.B(n_3412),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_7551),
.Y(n_8189)
);

INVx4_ASAP7_75t_SL g8190 ( 
.A(n_7587),
.Y(n_8190)
);

AND2x2_ASAP7_75t_L g8191 ( 
.A(n_7274),
.B(n_4423),
.Y(n_8191)
);

NOR2xp33_ASAP7_75t_L g8192 ( 
.A(n_7158),
.B(n_4424),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7564),
.Y(n_8193)
);

AND2x2_ASAP7_75t_L g8194 ( 
.A(n_7715),
.B(n_7486),
.Y(n_8194)
);

NAND2xp5_ASAP7_75t_L g8195 ( 
.A(n_7755),
.B(n_7181),
.Y(n_8195)
);

AOI22xp33_ASAP7_75t_L g8196 ( 
.A1(n_7724),
.A2(n_7167),
.B1(n_7143),
.B2(n_7614),
.Y(n_8196)
);

NAND2xp5_ASAP7_75t_L g8197 ( 
.A(n_8051),
.B(n_7266),
.Y(n_8197)
);

INVx2_ASAP7_75t_SL g8198 ( 
.A(n_8102),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7684),
.Y(n_8199)
);

NAND2xp5_ASAP7_75t_L g8200 ( 
.A(n_7804),
.B(n_7534),
.Y(n_8200)
);

INVx2_ASAP7_75t_L g8201 ( 
.A(n_7685),
.Y(n_8201)
);

INVx2_ASAP7_75t_SL g8202 ( 
.A(n_7742),
.Y(n_8202)
);

AND2x2_ASAP7_75t_L g8203 ( 
.A(n_7723),
.B(n_7302),
.Y(n_8203)
);

AOI22xp5_ASAP7_75t_L g8204 ( 
.A1(n_7817),
.A2(n_7238),
.B1(n_7396),
.B2(n_7295),
.Y(n_8204)
);

BUFx6f_ASAP7_75t_L g8205 ( 
.A(n_7742),
.Y(n_8205)
);

NAND2xp5_ASAP7_75t_SL g8206 ( 
.A(n_7875),
.B(n_7437),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7686),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_7687),
.Y(n_8208)
);

NAND2xp5_ASAP7_75t_SL g8209 ( 
.A(n_7694),
.B(n_7986),
.Y(n_8209)
);

NAND2xp33_ASAP7_75t_L g8210 ( 
.A(n_8053),
.B(n_7662),
.Y(n_8210)
);

NAND2xp5_ASAP7_75t_L g8211 ( 
.A(n_8058),
.B(n_7527),
.Y(n_8211)
);

INVxp67_ASAP7_75t_L g8212 ( 
.A(n_7691),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_8063),
.B(n_7642),
.Y(n_8213)
);

NOR2xp33_ASAP7_75t_L g8214 ( 
.A(n_7881),
.B(n_7372),
.Y(n_8214)
);

NAND2xp5_ASAP7_75t_L g8215 ( 
.A(n_8010),
.B(n_7665),
.Y(n_8215)
);

INVx1_ASAP7_75t_SL g8216 ( 
.A(n_7736),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_L g8217 ( 
.A(n_7997),
.B(n_7668),
.Y(n_8217)
);

NOR2xp33_ASAP7_75t_L g8218 ( 
.A(n_7772),
.B(n_7545),
.Y(n_8218)
);

INVx2_ASAP7_75t_L g8219 ( 
.A(n_7688),
.Y(n_8219)
);

OAI22xp5_ASAP7_75t_SL g8220 ( 
.A1(n_7693),
.A2(n_7506),
.B1(n_7497),
.B2(n_7596),
.Y(n_8220)
);

OA22x2_ASAP7_75t_L g8221 ( 
.A1(n_8118),
.A2(n_7157),
.B1(n_7368),
.B2(n_7329),
.Y(n_8221)
);

INVx2_ASAP7_75t_L g8222 ( 
.A(n_7689),
.Y(n_8222)
);

AND2x4_ASAP7_75t_L g8223 ( 
.A(n_7745),
.B(n_7592),
.Y(n_8223)
);

OR2x6_ASAP7_75t_L g8224 ( 
.A(n_7714),
.B(n_7282),
.Y(n_8224)
);

INVx3_ASAP7_75t_L g8225 ( 
.A(n_7884),
.Y(n_8225)
);

OAI22xp33_ASAP7_75t_L g8226 ( 
.A1(n_8101),
.A2(n_7447),
.B1(n_7437),
.B2(n_7497),
.Y(n_8226)
);

BUFx2_ASAP7_75t_SL g8227 ( 
.A(n_7741),
.Y(n_8227)
);

INVx2_ASAP7_75t_SL g8228 ( 
.A(n_7910),
.Y(n_8228)
);

OAI22xp5_ASAP7_75t_L g8229 ( 
.A1(n_8110),
.A2(n_7616),
.B1(n_7624),
.B2(n_7488),
.Y(n_8229)
);

OAI22xp33_ASAP7_75t_L g8230 ( 
.A1(n_8119),
.A2(n_7447),
.B1(n_7506),
.B2(n_7596),
.Y(n_8230)
);

NAND2xp33_ASAP7_75t_L g8231 ( 
.A(n_7771),
.B(n_7307),
.Y(n_8231)
);

OAI22xp5_ASAP7_75t_L g8232 ( 
.A1(n_8098),
.A2(n_7565),
.B1(n_7370),
.B2(n_7493),
.Y(n_8232)
);

INVx2_ASAP7_75t_L g8233 ( 
.A(n_7692),
.Y(n_8233)
);

NOR2xp33_ASAP7_75t_SL g8234 ( 
.A(n_7797),
.B(n_7802),
.Y(n_8234)
);

NAND2xp5_ASAP7_75t_SL g8235 ( 
.A(n_7833),
.B(n_7459),
.Y(n_8235)
);

BUFx6f_ASAP7_75t_L g8236 ( 
.A(n_7910),
.Y(n_8236)
);

NAND2xp5_ASAP7_75t_L g8237 ( 
.A(n_7895),
.B(n_8041),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7696),
.Y(n_8238)
);

INVx2_ASAP7_75t_L g8239 ( 
.A(n_7697),
.Y(n_8239)
);

NAND2xp5_ASAP7_75t_L g8240 ( 
.A(n_8042),
.B(n_8002),
.Y(n_8240)
);

AOI22xp33_ASAP7_75t_L g8241 ( 
.A1(n_8089),
.A2(n_7540),
.B1(n_7405),
.B2(n_7475),
.Y(n_8241)
);

INVx1_ASAP7_75t_L g8242 ( 
.A(n_7700),
.Y(n_8242)
);

NOR2xp33_ASAP7_75t_L g8243 ( 
.A(n_8052),
.B(n_7340),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7701),
.Y(n_8244)
);

INVxp67_ASAP7_75t_SL g8245 ( 
.A(n_7892),
.Y(n_8245)
);

INVx2_ASAP7_75t_L g8246 ( 
.A(n_7702),
.Y(n_8246)
);

INVx2_ASAP7_75t_L g8247 ( 
.A(n_7703),
.Y(n_8247)
);

NAND2xp5_ASAP7_75t_L g8248 ( 
.A(n_8003),
.B(n_7431),
.Y(n_8248)
);

NAND2xp5_ASAP7_75t_L g8249 ( 
.A(n_8060),
.B(n_7520),
.Y(n_8249)
);

NAND2xp5_ASAP7_75t_L g8250 ( 
.A(n_8036),
.B(n_7526),
.Y(n_8250)
);

NAND2xp5_ASAP7_75t_L g8251 ( 
.A(n_8039),
.B(n_7578),
.Y(n_8251)
);

O2A1O1Ixp33_ASAP7_75t_L g8252 ( 
.A1(n_8059),
.A2(n_7601),
.B(n_4526),
.C(n_4531),
.Y(n_8252)
);

NAND2xp5_ASAP7_75t_SL g8253 ( 
.A(n_7978),
.B(n_4425),
.Y(n_8253)
);

NAND2xp5_ASAP7_75t_L g8254 ( 
.A(n_8019),
.B(n_7549),
.Y(n_8254)
);

OR2x2_ASAP7_75t_L g8255 ( 
.A(n_7939),
.B(n_4426),
.Y(n_8255)
);

INVx1_ASAP7_75t_L g8256 ( 
.A(n_7704),
.Y(n_8256)
);

NAND2x1_ASAP7_75t_L g8257 ( 
.A(n_7695),
.B(n_4517),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7705),
.Y(n_8258)
);

A2O1A1Ixp33_ASAP7_75t_L g8259 ( 
.A1(n_7770),
.A2(n_7919),
.B(n_7850),
.C(n_7851),
.Y(n_8259)
);

NOR2xp33_ASAP7_75t_L g8260 ( 
.A(n_7935),
.B(n_7415),
.Y(n_8260)
);

NAND2xp5_ASAP7_75t_SL g8261 ( 
.A(n_8181),
.B(n_4428),
.Y(n_8261)
);

BUFx3_ASAP7_75t_L g8262 ( 
.A(n_8083),
.Y(n_8262)
);

OAI21xp33_ASAP7_75t_L g8263 ( 
.A1(n_8127),
.A2(n_4430),
.B(n_4429),
.Y(n_8263)
);

NAND2xp5_ASAP7_75t_L g8264 ( 
.A(n_8022),
.B(n_8025),
.Y(n_8264)
);

INVx2_ASAP7_75t_SL g8265 ( 
.A(n_7950),
.Y(n_8265)
);

AOI22xp5_ASAP7_75t_L g8266 ( 
.A1(n_7731),
.A2(n_7635),
.B1(n_4437),
.B2(n_4438),
.Y(n_8266)
);

NOR2xp33_ASAP7_75t_SL g8267 ( 
.A(n_7725),
.B(n_4431),
.Y(n_8267)
);

BUFx3_ASAP7_75t_L g8268 ( 
.A(n_8037),
.Y(n_8268)
);

NAND2xp5_ASAP7_75t_L g8269 ( 
.A(n_8031),
.B(n_4543),
.Y(n_8269)
);

NOR2xp33_ASAP7_75t_L g8270 ( 
.A(n_7889),
.B(n_4445),
.Y(n_8270)
);

NAND2xp5_ASAP7_75t_L g8271 ( 
.A(n_8033),
.B(n_4544),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_7958),
.B(n_4548),
.Y(n_8272)
);

NOR2xp33_ASAP7_75t_L g8273 ( 
.A(n_8153),
.B(n_4452),
.Y(n_8273)
);

INVx1_ASAP7_75t_L g8274 ( 
.A(n_7707),
.Y(n_8274)
);

NAND2xp5_ASAP7_75t_L g8275 ( 
.A(n_8038),
.B(n_4558),
.Y(n_8275)
);

NOR2xp33_ASAP7_75t_L g8276 ( 
.A(n_7995),
.B(n_4455),
.Y(n_8276)
);

NOR2xp33_ASAP7_75t_L g8277 ( 
.A(n_7751),
.B(n_8145),
.Y(n_8277)
);

O2A1O1Ixp33_ASAP7_75t_L g8278 ( 
.A1(n_7918),
.A2(n_4563),
.B(n_4570),
.C(n_4561),
.Y(n_8278)
);

NAND2xp5_ASAP7_75t_L g8279 ( 
.A(n_7890),
.B(n_8087),
.Y(n_8279)
);

NAND2xp5_ASAP7_75t_L g8280 ( 
.A(n_8056),
.B(n_4573),
.Y(n_8280)
);

INVx2_ASAP7_75t_SL g8281 ( 
.A(n_7950),
.Y(n_8281)
);

NAND2xp5_ASAP7_75t_L g8282 ( 
.A(n_8057),
.B(n_4584),
.Y(n_8282)
);

OAI221xp5_ASAP7_75t_L g8283 ( 
.A1(n_8134),
.A2(n_4594),
.B1(n_4596),
.B2(n_4592),
.C(n_4585),
.Y(n_8283)
);

NAND2xp5_ASAP7_75t_L g8284 ( 
.A(n_8065),
.B(n_4598),
.Y(n_8284)
);

AND2x2_ASAP7_75t_L g8285 ( 
.A(n_7976),
.B(n_4456),
.Y(n_8285)
);

NOR2xp33_ASAP7_75t_L g8286 ( 
.A(n_7729),
.B(n_4457),
.Y(n_8286)
);

INVx1_ASAP7_75t_L g8287 ( 
.A(n_7709),
.Y(n_8287)
);

NAND2xp5_ASAP7_75t_L g8288 ( 
.A(n_8066),
.B(n_4602),
.Y(n_8288)
);

INVx1_ASAP7_75t_L g8289 ( 
.A(n_7711),
.Y(n_8289)
);

NAND2xp5_ASAP7_75t_SL g8290 ( 
.A(n_7855),
.B(n_4460),
.Y(n_8290)
);

INVxp67_ASAP7_75t_L g8291 ( 
.A(n_7816),
.Y(n_8291)
);

NAND2xp5_ASAP7_75t_L g8292 ( 
.A(n_7858),
.B(n_4603),
.Y(n_8292)
);

INVx2_ASAP7_75t_SL g8293 ( 
.A(n_8027),
.Y(n_8293)
);

INVx2_ASAP7_75t_L g8294 ( 
.A(n_7712),
.Y(n_8294)
);

NOR2xp33_ASAP7_75t_L g8295 ( 
.A(n_8061),
.B(n_4461),
.Y(n_8295)
);

INVx1_ASAP7_75t_L g8296 ( 
.A(n_7713),
.Y(n_8296)
);

NAND2xp5_ASAP7_75t_L g8297 ( 
.A(n_7864),
.B(n_4605),
.Y(n_8297)
);

NOR2x1p5_ASAP7_75t_L g8298 ( 
.A(n_7752),
.B(n_4463),
.Y(n_8298)
);

AND2x2_ASAP7_75t_L g8299 ( 
.A(n_7829),
.B(n_4467),
.Y(n_8299)
);

NOR3xp33_ASAP7_75t_L g8300 ( 
.A(n_7991),
.B(n_8069),
.C(n_8024),
.Y(n_8300)
);

HB1xp67_ASAP7_75t_L g8301 ( 
.A(n_7806),
.Y(n_8301)
);

AND2x2_ASAP7_75t_SL g8302 ( 
.A(n_7734),
.B(n_4607),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7717),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_L g8304 ( 
.A(n_7882),
.B(n_4608),
.Y(n_8304)
);

NAND2xp5_ASAP7_75t_L g8305 ( 
.A(n_7885),
.B(n_4610),
.Y(n_8305)
);

AOI22xp5_ASAP7_75t_L g8306 ( 
.A1(n_7799),
.A2(n_4476),
.B1(n_4478),
.B2(n_4468),
.Y(n_8306)
);

INVx2_ASAP7_75t_L g8307 ( 
.A(n_7718),
.Y(n_8307)
);

AOI22xp33_ASAP7_75t_L g8308 ( 
.A1(n_8026),
.A2(n_4619),
.B1(n_4622),
.B2(n_4617),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_7849),
.B(n_4479),
.Y(n_8309)
);

NAND2xp5_ASAP7_75t_L g8310 ( 
.A(n_7903),
.B(n_7941),
.Y(n_8310)
);

INVx2_ASAP7_75t_L g8311 ( 
.A(n_7719),
.Y(n_8311)
);

AOI22xp5_ASAP7_75t_L g8312 ( 
.A1(n_7794),
.A2(n_4482),
.B1(n_4483),
.B2(n_4480),
.Y(n_8312)
);

INVx2_ASAP7_75t_L g8313 ( 
.A(n_7721),
.Y(n_8313)
);

INVx3_ASAP7_75t_L g8314 ( 
.A(n_7871),
.Y(n_8314)
);

BUFx12f_ASAP7_75t_SL g8315 ( 
.A(n_8027),
.Y(n_8315)
);

INVxp33_ASAP7_75t_L g8316 ( 
.A(n_7867),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7722),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_7727),
.Y(n_8318)
);

NOR2xp33_ASAP7_75t_L g8319 ( 
.A(n_7967),
.B(n_4488),
.Y(n_8319)
);

NAND2xp5_ASAP7_75t_L g8320 ( 
.A(n_7956),
.B(n_4629),
.Y(n_8320)
);

AOI22xp5_ASAP7_75t_L g8321 ( 
.A1(n_8020),
.A2(n_4494),
.B1(n_4495),
.B2(n_4493),
.Y(n_8321)
);

O2A1O1Ixp33_ASAP7_75t_L g8322 ( 
.A1(n_7809),
.A2(n_4636),
.B(n_4642),
.C(n_4635),
.Y(n_8322)
);

AND2x2_ASAP7_75t_L g8323 ( 
.A(n_7894),
.B(n_4496),
.Y(n_8323)
);

NAND2xp5_ASAP7_75t_L g8324 ( 
.A(n_7932),
.B(n_4652),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_7728),
.Y(n_8325)
);

A2O1A1Ixp33_ASAP7_75t_L g8326 ( 
.A1(n_8192),
.A2(n_4657),
.B(n_4659),
.C(n_4654),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_7730),
.Y(n_8327)
);

INVx2_ASAP7_75t_L g8328 ( 
.A(n_7733),
.Y(n_8328)
);

INVx2_ASAP7_75t_L g8329 ( 
.A(n_7735),
.Y(n_8329)
);

NOR2xp33_ASAP7_75t_L g8330 ( 
.A(n_7944),
.B(n_4498),
.Y(n_8330)
);

INVx2_ASAP7_75t_L g8331 ( 
.A(n_7737),
.Y(n_8331)
);

AOI22xp33_ASAP7_75t_L g8332 ( 
.A1(n_8135),
.A2(n_4669),
.B1(n_4670),
.B2(n_4667),
.Y(n_8332)
);

NOR2xp33_ASAP7_75t_L g8333 ( 
.A(n_7957),
.B(n_4499),
.Y(n_8333)
);

OAI221xp5_ASAP7_75t_L g8334 ( 
.A1(n_8142),
.A2(n_4678),
.B1(n_4687),
.B2(n_4677),
.C(n_4676),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7738),
.Y(n_8335)
);

AND2x2_ASAP7_75t_L g8336 ( 
.A(n_7822),
.B(n_7853),
.Y(n_8336)
);

INVx3_ASAP7_75t_L g8337 ( 
.A(n_7866),
.Y(n_8337)
);

OR2x6_ASAP7_75t_L g8338 ( 
.A(n_7891),
.B(n_4688),
.Y(n_8338)
);

AND2x2_ASAP7_75t_L g8339 ( 
.A(n_7869),
.B(n_4500),
.Y(n_8339)
);

AOI21xp5_ASAP7_75t_L g8340 ( 
.A1(n_8174),
.A2(n_4702),
.B(n_4694),
.Y(n_8340)
);

NAND2xp5_ASAP7_75t_L g8341 ( 
.A(n_8006),
.B(n_4704),
.Y(n_8341)
);

AOI22xp5_ASAP7_75t_L g8342 ( 
.A1(n_7768),
.A2(n_4505),
.B1(n_4506),
.B2(n_4503),
.Y(n_8342)
);

INVx1_ASAP7_75t_L g8343 ( 
.A(n_7740),
.Y(n_8343)
);

O2A1O1Ixp5_ASAP7_75t_L g8344 ( 
.A1(n_7899),
.A2(n_4711),
.B(n_4716),
.C(n_4706),
.Y(n_8344)
);

HB1xp67_ASAP7_75t_L g8345 ( 
.A(n_8190),
.Y(n_8345)
);

INVxp67_ASAP7_75t_L g8346 ( 
.A(n_8092),
.Y(n_8346)
);

INVx4_ASAP7_75t_L g8347 ( 
.A(n_8190),
.Y(n_8347)
);

INVx8_ASAP7_75t_L g8348 ( 
.A(n_8162),
.Y(n_8348)
);

INVx2_ASAP7_75t_SL g8349 ( 
.A(n_8064),
.Y(n_8349)
);

OAI22xp33_ASAP7_75t_L g8350 ( 
.A1(n_7823),
.A2(n_4509),
.B1(n_4511),
.B2(n_4507),
.Y(n_8350)
);

O2A1O1Ixp33_ASAP7_75t_L g8351 ( 
.A1(n_8017),
.A2(n_4730),
.B(n_4735),
.C(n_4717),
.Y(n_8351)
);

AOI22xp5_ASAP7_75t_L g8352 ( 
.A1(n_7739),
.A2(n_4515),
.B1(n_4516),
.B2(n_4513),
.Y(n_8352)
);

NAND2xp5_ASAP7_75t_SL g8353 ( 
.A(n_7837),
.B(n_4518),
.Y(n_8353)
);

NOR3xp33_ASAP7_75t_L g8354 ( 
.A(n_7746),
.B(n_4743),
.C(n_4740),
.Y(n_8354)
);

NAND2xp33_ASAP7_75t_L g8355 ( 
.A(n_7982),
.B(n_4519),
.Y(n_8355)
);

INVx2_ASAP7_75t_SL g8356 ( 
.A(n_8064),
.Y(n_8356)
);

INVx2_ASAP7_75t_SL g8357 ( 
.A(n_8112),
.Y(n_8357)
);

NAND2xp5_ASAP7_75t_L g8358 ( 
.A(n_8040),
.B(n_4744),
.Y(n_8358)
);

AND2x2_ASAP7_75t_L g8359 ( 
.A(n_7915),
.B(n_4520),
.Y(n_8359)
);

NOR2xp33_ASAP7_75t_L g8360 ( 
.A(n_7769),
.B(n_4521),
.Y(n_8360)
);

INVx3_ASAP7_75t_L g8361 ( 
.A(n_8112),
.Y(n_8361)
);

NAND2xp5_ASAP7_75t_L g8362 ( 
.A(n_8062),
.B(n_4746),
.Y(n_8362)
);

BUFx6f_ASAP7_75t_SL g8363 ( 
.A(n_7726),
.Y(n_8363)
);

NAND2xp5_ASAP7_75t_L g8364 ( 
.A(n_7861),
.B(n_4747),
.Y(n_8364)
);

INVx1_ASAP7_75t_L g8365 ( 
.A(n_7743),
.Y(n_8365)
);

INVxp67_ASAP7_75t_SL g8366 ( 
.A(n_7922),
.Y(n_8366)
);

BUFx3_ASAP7_75t_L g8367 ( 
.A(n_7776),
.Y(n_8367)
);

NAND2xp5_ASAP7_75t_L g8368 ( 
.A(n_7873),
.B(n_4748),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_7744),
.Y(n_8369)
);

AOI22xp5_ASAP7_75t_L g8370 ( 
.A1(n_7795),
.A2(n_4523),
.B1(n_4525),
.B2(n_4522),
.Y(n_8370)
);

NAND2xp5_ASAP7_75t_SL g8371 ( 
.A(n_7710),
.B(n_4527),
.Y(n_8371)
);

OAI22xp5_ASAP7_75t_L g8372 ( 
.A1(n_7748),
.A2(n_4530),
.B1(n_4532),
.B2(n_4529),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7750),
.Y(n_8373)
);

NOR2xp33_ASAP7_75t_L g8374 ( 
.A(n_8047),
.B(n_4534),
.Y(n_8374)
);

INVx2_ASAP7_75t_L g8375 ( 
.A(n_7753),
.Y(n_8375)
);

NOR2xp67_ASAP7_75t_L g8376 ( 
.A(n_7859),
.B(n_3413),
.Y(n_8376)
);

A2O1A1Ixp33_ASAP7_75t_L g8377 ( 
.A1(n_8144),
.A2(n_4752),
.B(n_4753),
.C(n_4750),
.Y(n_8377)
);

NAND2xp5_ASAP7_75t_L g8378 ( 
.A(n_7754),
.B(n_7756),
.Y(n_8378)
);

NAND2xp5_ASAP7_75t_L g8379 ( 
.A(n_7757),
.B(n_4754),
.Y(n_8379)
);

NAND2xp5_ASAP7_75t_L g8380 ( 
.A(n_7758),
.B(n_4759),
.Y(n_8380)
);

BUFx6f_ASAP7_75t_L g8381 ( 
.A(n_7838),
.Y(n_8381)
);

BUFx3_ASAP7_75t_L g8382 ( 
.A(n_7778),
.Y(n_8382)
);

NAND2xp5_ASAP7_75t_L g8383 ( 
.A(n_7760),
.B(n_4760),
.Y(n_8383)
);

BUFx6f_ASAP7_75t_L g8384 ( 
.A(n_7974),
.Y(n_8384)
);

AOI221xp5_ASAP7_75t_L g8385 ( 
.A1(n_8106),
.A2(n_4770),
.B1(n_4771),
.B2(n_4767),
.C(n_4765),
.Y(n_8385)
);

AND2x2_ASAP7_75t_L g8386 ( 
.A(n_7917),
.B(n_4537),
.Y(n_8386)
);

AND2x4_ASAP7_75t_SL g8387 ( 
.A(n_7779),
.B(n_4774),
.Y(n_8387)
);

AND2x2_ASAP7_75t_L g8388 ( 
.A(n_8050),
.B(n_4538),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7761),
.Y(n_8389)
);

INVx8_ASAP7_75t_L g8390 ( 
.A(n_8005),
.Y(n_8390)
);

NAND2xp5_ASAP7_75t_L g8391 ( 
.A(n_7762),
.B(n_4777),
.Y(n_8391)
);

AOI22xp33_ASAP7_75t_L g8392 ( 
.A1(n_8188),
.A2(n_4786),
.B1(n_4791),
.B2(n_4779),
.Y(n_8392)
);

INVx1_ASAP7_75t_L g8393 ( 
.A(n_7813),
.Y(n_8393)
);

NOR2xp67_ASAP7_75t_L g8394 ( 
.A(n_7874),
.B(n_3414),
.Y(n_8394)
);

NAND2xp5_ASAP7_75t_SL g8395 ( 
.A(n_7832),
.B(n_4540),
.Y(n_8395)
);

BUFx3_ASAP7_75t_L g8396 ( 
.A(n_7877),
.Y(n_8396)
);

NAND2xp5_ASAP7_75t_SL g8397 ( 
.A(n_8163),
.B(n_4542),
.Y(n_8397)
);

NAND2xp5_ASAP7_75t_L g8398 ( 
.A(n_7763),
.B(n_4792),
.Y(n_8398)
);

INVx2_ASAP7_75t_L g8399 ( 
.A(n_7972),
.Y(n_8399)
);

OAI22xp5_ASAP7_75t_L g8400 ( 
.A1(n_7814),
.A2(n_4549),
.B1(n_4550),
.B2(n_4547),
.Y(n_8400)
);

INVx2_ASAP7_75t_L g8401 ( 
.A(n_7973),
.Y(n_8401)
);

NAND2xp5_ASAP7_75t_L g8402 ( 
.A(n_7764),
.B(n_4794),
.Y(n_8402)
);

INVx3_ASAP7_75t_L g8403 ( 
.A(n_8177),
.Y(n_8403)
);

INVx1_ASAP7_75t_L g8404 ( 
.A(n_7815),
.Y(n_8404)
);

NAND2xp5_ASAP7_75t_L g8405 ( 
.A(n_7766),
.B(n_4798),
.Y(n_8405)
);

OR2x6_ASAP7_75t_L g8406 ( 
.A(n_7720),
.B(n_4810),
.Y(n_8406)
);

INVx3_ASAP7_75t_L g8407 ( 
.A(n_8072),
.Y(n_8407)
);

INVx1_ASAP7_75t_L g8408 ( 
.A(n_7818),
.Y(n_8408)
);

AO22x1_ASAP7_75t_L g8409 ( 
.A1(n_7845),
.A2(n_4553),
.B1(n_4554),
.B2(n_4551),
.Y(n_8409)
);

NAND2xp5_ASAP7_75t_L g8410 ( 
.A(n_7773),
.B(n_4815),
.Y(n_8410)
);

NAND2xp5_ASAP7_75t_SL g8411 ( 
.A(n_8164),
.B(n_4555),
.Y(n_8411)
);

NAND2xp5_ASAP7_75t_SL g8412 ( 
.A(n_8165),
.B(n_4559),
.Y(n_8412)
);

NOR2xp33_ASAP7_75t_L g8413 ( 
.A(n_8108),
.B(n_4564),
.Y(n_8413)
);

AND2x2_ASAP7_75t_L g8414 ( 
.A(n_7901),
.B(n_4566),
.Y(n_8414)
);

INVx2_ASAP7_75t_L g8415 ( 
.A(n_7980),
.Y(n_8415)
);

INVxp67_ASAP7_75t_L g8416 ( 
.A(n_7857),
.Y(n_8416)
);

NAND2xp5_ASAP7_75t_L g8417 ( 
.A(n_7777),
.B(n_4820),
.Y(n_8417)
);

INVx2_ASAP7_75t_L g8418 ( 
.A(n_7981),
.Y(n_8418)
);

BUFx6f_ASAP7_75t_L g8419 ( 
.A(n_8023),
.Y(n_8419)
);

NAND2xp5_ASAP7_75t_L g8420 ( 
.A(n_7780),
.B(n_4829),
.Y(n_8420)
);

NAND2xp5_ASAP7_75t_L g8421 ( 
.A(n_7782),
.B(n_4844),
.Y(n_8421)
);

NAND2xp5_ASAP7_75t_SL g8422 ( 
.A(n_8075),
.B(n_4567),
.Y(n_8422)
);

AOI22xp33_ASAP7_75t_SL g8423 ( 
.A1(n_8018),
.A2(n_8125),
.B1(n_8120),
.B2(n_8121),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_7819),
.Y(n_8424)
);

AOI22xp5_ASAP7_75t_L g8425 ( 
.A1(n_8078),
.A2(n_4572),
.B1(n_4575),
.B2(n_4568),
.Y(n_8425)
);

NAND2xp5_ASAP7_75t_L g8426 ( 
.A(n_7785),
.B(n_7789),
.Y(n_8426)
);

NAND2xp5_ASAP7_75t_L g8427 ( 
.A(n_7790),
.B(n_4846),
.Y(n_8427)
);

NAND2xp5_ASAP7_75t_L g8428 ( 
.A(n_7793),
.B(n_4849),
.Y(n_8428)
);

INVx1_ASAP7_75t_L g8429 ( 
.A(n_7820),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_7821),
.Y(n_8430)
);

NAND2xp5_ASAP7_75t_L g8431 ( 
.A(n_7796),
.B(n_7798),
.Y(n_8431)
);

INVx2_ASAP7_75t_SL g8432 ( 
.A(n_8140),
.Y(n_8432)
);

INVx2_ASAP7_75t_L g8433 ( 
.A(n_7983),
.Y(n_8433)
);

AOI22xp5_ASAP7_75t_L g8434 ( 
.A1(n_8011),
.A2(n_4577),
.B1(n_4579),
.B2(n_4576),
.Y(n_8434)
);

INVx1_ASAP7_75t_L g8435 ( 
.A(n_7824),
.Y(n_8435)
);

O2A1O1Ixp33_ASAP7_75t_L g8436 ( 
.A1(n_8171),
.A2(n_4861),
.B(n_4863),
.C(n_4855),
.Y(n_8436)
);

NOR2xp67_ASAP7_75t_L g8437 ( 
.A(n_7902),
.B(n_7923),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7825),
.Y(n_8438)
);

OR2x2_ASAP7_75t_L g8439 ( 
.A(n_7876),
.B(n_4581),
.Y(n_8439)
);

INVx1_ASAP7_75t_L g8440 ( 
.A(n_7826),
.Y(n_8440)
);

A2O1A1Ixp33_ASAP7_75t_L g8441 ( 
.A1(n_8124),
.A2(n_4878),
.B(n_4879),
.C(n_4866),
.Y(n_8441)
);

NOR2xp33_ASAP7_75t_L g8442 ( 
.A(n_8088),
.B(n_7791),
.Y(n_8442)
);

INVx2_ASAP7_75t_L g8443 ( 
.A(n_7984),
.Y(n_8443)
);

NOR2xp33_ASAP7_75t_L g8444 ( 
.A(n_7872),
.B(n_4582),
.Y(n_8444)
);

NOR2xp33_ASAP7_75t_L g8445 ( 
.A(n_7834),
.B(n_8161),
.Y(n_8445)
);

NAND2xp5_ASAP7_75t_L g8446 ( 
.A(n_7800),
.B(n_7801),
.Y(n_8446)
);

NAND2xp5_ASAP7_75t_L g8447 ( 
.A(n_7803),
.B(n_7805),
.Y(n_8447)
);

OAI21xp5_ASAP7_75t_L g8448 ( 
.A1(n_8160),
.A2(n_4894),
.B(n_4893),
.Y(n_8448)
);

NAND2xp5_ASAP7_75t_L g8449 ( 
.A(n_7808),
.B(n_4902),
.Y(n_8449)
);

OR2x6_ASAP7_75t_L g8450 ( 
.A(n_7690),
.B(n_7706),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7828),
.Y(n_8451)
);

NAND2xp5_ASAP7_75t_L g8452 ( 
.A(n_7810),
.B(n_4916),
.Y(n_8452)
);

NAND2xp5_ASAP7_75t_SL g8453 ( 
.A(n_8030),
.B(n_4583),
.Y(n_8453)
);

NAND2xp5_ASAP7_75t_L g8454 ( 
.A(n_7811),
.B(n_4917),
.Y(n_8454)
);

INVxp67_ASAP7_75t_SL g8455 ( 
.A(n_7831),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_7812),
.B(n_4918),
.Y(n_8456)
);

AND2x6_ASAP7_75t_SL g8457 ( 
.A(n_7716),
.B(n_4921),
.Y(n_8457)
);

HB1xp67_ASAP7_75t_L g8458 ( 
.A(n_8035),
.Y(n_8458)
);

CKINVDCx20_ASAP7_75t_R g8459 ( 
.A(n_7699),
.Y(n_8459)
);

AOI22xp33_ASAP7_75t_L g8460 ( 
.A1(n_8044),
.A2(n_4926),
.B1(n_4936),
.B2(n_4924),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_7835),
.Y(n_8461)
);

HB1xp67_ASAP7_75t_L g8462 ( 
.A(n_8043),
.Y(n_8462)
);

OR2x6_ASAP7_75t_L g8463 ( 
.A(n_7767),
.B(n_8136),
.Y(n_8463)
);

INVx2_ASAP7_75t_L g8464 ( 
.A(n_7985),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_L g8465 ( 
.A(n_7836),
.B(n_4937),
.Y(n_8465)
);

INVx2_ASAP7_75t_L g8466 ( 
.A(n_7839),
.Y(n_8466)
);

AND2x2_ASAP7_75t_L g8467 ( 
.A(n_7993),
.B(n_4590),
.Y(n_8467)
);

NAND2xp5_ASAP7_75t_L g8468 ( 
.A(n_7840),
.B(n_4941),
.Y(n_8468)
);

BUFx5_ASAP7_75t_L g8469 ( 
.A(n_8130),
.Y(n_8469)
);

BUFx6f_ASAP7_75t_SL g8470 ( 
.A(n_7880),
.Y(n_8470)
);

NOR2xp33_ASAP7_75t_L g8471 ( 
.A(n_7988),
.B(n_4595),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_7844),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_7846),
.B(n_7848),
.Y(n_8473)
);

INVx2_ASAP7_75t_L g8474 ( 
.A(n_7856),
.Y(n_8474)
);

NOR2xp33_ASAP7_75t_L g8475 ( 
.A(n_7708),
.B(n_4599),
.Y(n_8475)
);

NAND2xp5_ASAP7_75t_SL g8476 ( 
.A(n_8175),
.B(n_4604),
.Y(n_8476)
);

AOI22xp33_ASAP7_75t_L g8477 ( 
.A1(n_8046),
.A2(n_4955),
.B1(n_4956),
.B2(n_4944),
.Y(n_8477)
);

NAND2xp5_ASAP7_75t_L g8478 ( 
.A(n_7860),
.B(n_4606),
.Y(n_8478)
);

INVx2_ASAP7_75t_L g8479 ( 
.A(n_7862),
.Y(n_8479)
);

NOR2xp33_ASAP7_75t_L g8480 ( 
.A(n_7963),
.B(n_4613),
.Y(n_8480)
);

INVx2_ASAP7_75t_L g8481 ( 
.A(n_7863),
.Y(n_8481)
);

NAND2xp5_ASAP7_75t_L g8482 ( 
.A(n_7765),
.B(n_7774),
.Y(n_8482)
);

INVx1_ASAP7_75t_L g8483 ( 
.A(n_7827),
.Y(n_8483)
);

AOI22xp33_ASAP7_75t_L g8484 ( 
.A1(n_8104),
.A2(n_4615),
.B1(n_4618),
.B2(n_4614),
.Y(n_8484)
);

NOR3xp33_ASAP7_75t_L g8485 ( 
.A(n_8107),
.B(n_4625),
.C(n_4624),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_7698),
.Y(n_8486)
);

NOR2xp33_ASAP7_75t_L g8487 ( 
.A(n_7916),
.B(n_4628),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_7747),
.Y(n_8488)
);

INVx1_ASAP7_75t_L g8489 ( 
.A(n_7865),
.Y(n_8489)
);

AOI21xp5_ASAP7_75t_L g8490 ( 
.A1(n_8071),
.A2(n_3416),
.B(n_3415),
.Y(n_8490)
);

BUFx6f_ASAP7_75t_SL g8491 ( 
.A(n_8055),
.Y(n_8491)
);

NAND2xp5_ASAP7_75t_L g8492 ( 
.A(n_7783),
.B(n_4630),
.Y(n_8492)
);

INVx2_ASAP7_75t_L g8493 ( 
.A(n_8054),
.Y(n_8493)
);

NAND2xp5_ASAP7_75t_SL g8494 ( 
.A(n_8028),
.B(n_4632),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_7868),
.Y(n_8495)
);

AOI22xp5_ASAP7_75t_L g8496 ( 
.A1(n_8147),
.A2(n_4634),
.B1(n_4638),
.B2(n_4633),
.Y(n_8496)
);

NOR3xp33_ASAP7_75t_L g8497 ( 
.A(n_7998),
.B(n_4640),
.C(n_4639),
.Y(n_8497)
);

NAND2xp5_ASAP7_75t_L g8498 ( 
.A(n_7784),
.B(n_4643),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_7786),
.B(n_4644),
.Y(n_8499)
);

NAND2xp5_ASAP7_75t_L g8500 ( 
.A(n_7788),
.B(n_7792),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7887),
.Y(n_8501)
);

NAND2xp5_ASAP7_75t_L g8502 ( 
.A(n_7807),
.B(n_4645),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_L g8503 ( 
.A(n_7888),
.B(n_7893),
.Y(n_8503)
);

NAND2xp5_ASAP7_75t_L g8504 ( 
.A(n_7896),
.B(n_4646),
.Y(n_8504)
);

NAND2xp5_ASAP7_75t_SL g8505 ( 
.A(n_8082),
.B(n_4649),
.Y(n_8505)
);

AOI22xp33_ASAP7_75t_L g8506 ( 
.A1(n_8109),
.A2(n_4651),
.B1(n_4655),
.B2(n_4650),
.Y(n_8506)
);

INVx2_ASAP7_75t_L g8507 ( 
.A(n_7830),
.Y(n_8507)
);

NAND2xp5_ASAP7_75t_SL g8508 ( 
.A(n_7920),
.B(n_4656),
.Y(n_8508)
);

NOR2xp33_ASAP7_75t_SL g8509 ( 
.A(n_8029),
.B(n_4658),
.Y(n_8509)
);

NOR2xp33_ASAP7_75t_L g8510 ( 
.A(n_8096),
.B(n_8115),
.Y(n_8510)
);

NAND2xp5_ASAP7_75t_L g8511 ( 
.A(n_7897),
.B(n_4664),
.Y(n_8511)
);

AOI22xp5_ASAP7_75t_L g8512 ( 
.A1(n_8123),
.A2(n_4666),
.B1(n_4668),
.B2(n_4665),
.Y(n_8512)
);

INVx2_ASAP7_75t_L g8513 ( 
.A(n_7968),
.Y(n_8513)
);

INVx2_ASAP7_75t_L g8514 ( 
.A(n_7969),
.Y(n_8514)
);

NAND2xp5_ASAP7_75t_L g8515 ( 
.A(n_7990),
.B(n_4672),
.Y(n_8515)
);

NAND2xp5_ASAP7_75t_L g8516 ( 
.A(n_8122),
.B(n_4674),
.Y(n_8516)
);

INVx2_ASAP7_75t_L g8517 ( 
.A(n_7841),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_7992),
.Y(n_8518)
);

INVx2_ASAP7_75t_SL g8519 ( 
.A(n_8158),
.Y(n_8519)
);

NAND2xp5_ASAP7_75t_L g8520 ( 
.A(n_8168),
.B(n_4675),
.Y(n_8520)
);

NAND2xp5_ASAP7_75t_SL g8521 ( 
.A(n_8113),
.B(n_8129),
.Y(n_8521)
);

BUFx5_ASAP7_75t_L g8522 ( 
.A(n_8132),
.Y(n_8522)
);

HB1xp67_ASAP7_75t_L g8523 ( 
.A(n_8169),
.Y(n_8523)
);

CKINVDCx5p33_ASAP7_75t_R g8524 ( 
.A(n_7732),
.Y(n_8524)
);

NAND2xp5_ASAP7_75t_L g8525 ( 
.A(n_8191),
.B(n_7905),
.Y(n_8525)
);

NOR3xp33_ASAP7_75t_L g8526 ( 
.A(n_8086),
.B(n_4681),
.C(n_4679),
.Y(n_8526)
);

CKINVDCx5p33_ASAP7_75t_R g8527 ( 
.A(n_8016),
.Y(n_8527)
);

INVx2_ASAP7_75t_L g8528 ( 
.A(n_7842),
.Y(n_8528)
);

INVx2_ASAP7_75t_L g8529 ( 
.A(n_7843),
.Y(n_8529)
);

OAI22xp5_ASAP7_75t_SL g8530 ( 
.A1(n_7940),
.A2(n_4686),
.B1(n_4689),
.B2(n_4684),
.Y(n_8530)
);

INVx2_ASAP7_75t_L g8531 ( 
.A(n_7852),
.Y(n_8531)
);

BUFx12f_ASAP7_75t_SL g8532 ( 
.A(n_8084),
.Y(n_8532)
);

AOI22xp33_ASAP7_75t_L g8533 ( 
.A1(n_8152),
.A2(n_4691),
.B1(n_4692),
.B2(n_4690),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_L g8534 ( 
.A(n_7906),
.B(n_4693),
.Y(n_8534)
);

NOR2xp33_ASAP7_75t_SL g8535 ( 
.A(n_7879),
.B(n_4695),
.Y(n_8535)
);

INVx2_ASAP7_75t_L g8536 ( 
.A(n_7854),
.Y(n_8536)
);

AOI22xp33_ASAP7_75t_L g8537 ( 
.A1(n_7947),
.A2(n_4697),
.B1(n_4698),
.B2(n_4696),
.Y(n_8537)
);

OAI22xp33_ASAP7_75t_L g8538 ( 
.A1(n_7904),
.A2(n_4701),
.B1(n_4703),
.B2(n_4700),
.Y(n_8538)
);

A2O1A1Ixp33_ASAP7_75t_L g8539 ( 
.A1(n_7759),
.A2(n_4707),
.B(n_4708),
.C(n_4705),
.Y(n_8539)
);

OAI22xp5_ASAP7_75t_L g8540 ( 
.A1(n_7907),
.A2(n_4713),
.B1(n_4714),
.B2(n_4712),
.Y(n_8540)
);

BUFx6f_ASAP7_75t_L g8541 ( 
.A(n_8117),
.Y(n_8541)
);

NAND3xp33_ASAP7_75t_L g8542 ( 
.A(n_8137),
.B(n_4720),
.C(n_4719),
.Y(n_8542)
);

NAND2xp5_ASAP7_75t_L g8543 ( 
.A(n_7908),
.B(n_4721),
.Y(n_8543)
);

NAND2xp5_ASAP7_75t_SL g8544 ( 
.A(n_8141),
.B(n_4722),
.Y(n_8544)
);

NAND2xp5_ASAP7_75t_L g8545 ( 
.A(n_7909),
.B(n_4725),
.Y(n_8545)
);

AOI22xp33_ASAP7_75t_L g8546 ( 
.A1(n_8090),
.A2(n_4728),
.B1(n_4729),
.B2(n_4726),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_7912),
.B(n_4731),
.Y(n_8547)
);

OAI221xp5_ASAP7_75t_L g8548 ( 
.A1(n_8012),
.A2(n_4736),
.B1(n_4737),
.B2(n_4733),
.C(n_4732),
.Y(n_8548)
);

NAND2xp5_ASAP7_75t_L g8549 ( 
.A(n_7914),
.B(n_7921),
.Y(n_8549)
);

INVx1_ASAP7_75t_L g8550 ( 
.A(n_7924),
.Y(n_8550)
);

INVx2_ASAP7_75t_SL g8551 ( 
.A(n_8167),
.Y(n_8551)
);

NAND2xp5_ASAP7_75t_L g8552 ( 
.A(n_7925),
.B(n_7927),
.Y(n_8552)
);

NAND2xp5_ASAP7_75t_L g8553 ( 
.A(n_7928),
.B(n_4739),
.Y(n_8553)
);

NAND2xp5_ASAP7_75t_L g8554 ( 
.A(n_7929),
.B(n_4741),
.Y(n_8554)
);

NOR2xp33_ASAP7_75t_L g8555 ( 
.A(n_8111),
.B(n_4742),
.Y(n_8555)
);

INVx2_ASAP7_75t_L g8556 ( 
.A(n_7878),
.Y(n_8556)
);

INVx2_ASAP7_75t_L g8557 ( 
.A(n_7900),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_7933),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_7934),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_7911),
.Y(n_8560)
);

NOR2xp33_ASAP7_75t_L g8561 ( 
.A(n_8126),
.B(n_4745),
.Y(n_8561)
);

AOI22xp5_ASAP7_75t_L g8562 ( 
.A1(n_8131),
.A2(n_4755),
.B1(n_4761),
.B2(n_4749),
.Y(n_8562)
);

NAND2xp5_ASAP7_75t_L g8563 ( 
.A(n_7936),
.B(n_4762),
.Y(n_8563)
);

OAI21xp5_ASAP7_75t_L g8564 ( 
.A1(n_8048),
.A2(n_4769),
.B(n_4768),
.Y(n_8564)
);

AND2x2_ASAP7_75t_L g8565 ( 
.A(n_7926),
.B(n_4772),
.Y(n_8565)
);

NOR2xp33_ASAP7_75t_SL g8566 ( 
.A(n_7937),
.B(n_4773),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7938),
.Y(n_8567)
);

NOR2xp33_ASAP7_75t_L g8568 ( 
.A(n_8143),
.B(n_4775),
.Y(n_8568)
);

INVx2_ASAP7_75t_L g8569 ( 
.A(n_7913),
.Y(n_8569)
);

AND2x2_ASAP7_75t_L g8570 ( 
.A(n_8068),
.B(n_4778),
.Y(n_8570)
);

INVx1_ASAP7_75t_L g8571 ( 
.A(n_7942),
.Y(n_8571)
);

OAI22xp5_ASAP7_75t_L g8572 ( 
.A1(n_7943),
.A2(n_4787),
.B1(n_4788),
.B2(n_4782),
.Y(n_8572)
);

NAND2xp5_ASAP7_75t_L g8573 ( 
.A(n_7945),
.B(n_4789),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_7946),
.Y(n_8574)
);

NAND2xp5_ASAP7_75t_L g8575 ( 
.A(n_7948),
.B(n_4790),
.Y(n_8575)
);

INVx3_ASAP7_75t_L g8576 ( 
.A(n_8178),
.Y(n_8576)
);

O2A1O1Ixp33_ASAP7_75t_L g8577 ( 
.A1(n_8156),
.A2(n_4795),
.B(n_4796),
.C(n_4793),
.Y(n_8577)
);

NAND2xp5_ASAP7_75t_L g8578 ( 
.A(n_7951),
.B(n_4797),
.Y(n_8578)
);

NAND2xp5_ASAP7_75t_SL g8579 ( 
.A(n_8151),
.B(n_8099),
.Y(n_8579)
);

NAND2xp5_ASAP7_75t_L g8580 ( 
.A(n_7954),
.B(n_4799),
.Y(n_8580)
);

BUFx6f_ASAP7_75t_L g8581 ( 
.A(n_8138),
.Y(n_8581)
);

INVx2_ASAP7_75t_SL g8582 ( 
.A(n_8166),
.Y(n_8582)
);

NOR2xp33_ASAP7_75t_SL g8583 ( 
.A(n_7886),
.B(n_4805),
.Y(n_8583)
);

INVx2_ASAP7_75t_L g8584 ( 
.A(n_7952),
.Y(n_8584)
);

INVx1_ASAP7_75t_L g8585 ( 
.A(n_7955),
.Y(n_8585)
);

INVxp67_ASAP7_75t_L g8586 ( 
.A(n_8186),
.Y(n_8586)
);

INVx2_ASAP7_75t_L g8587 ( 
.A(n_7953),
.Y(n_8587)
);

HB1xp67_ASAP7_75t_L g8588 ( 
.A(n_8045),
.Y(n_8588)
);

BUFx3_ASAP7_75t_L g8589 ( 
.A(n_8148),
.Y(n_8589)
);

NOR2xp67_ASAP7_75t_L g8590 ( 
.A(n_8093),
.B(n_3417),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_7959),
.Y(n_8591)
);

NAND2xp5_ASAP7_75t_L g8592 ( 
.A(n_7960),
.B(n_4807),
.Y(n_8592)
);

NOR2xp33_ASAP7_75t_L g8593 ( 
.A(n_8094),
.B(n_4808),
.Y(n_8593)
);

NOR2xp33_ASAP7_75t_L g8594 ( 
.A(n_8097),
.B(n_4809),
.Y(n_8594)
);

NAND2xp5_ASAP7_75t_L g8595 ( 
.A(n_7962),
.B(n_4811),
.Y(n_8595)
);

INVxp67_ASAP7_75t_L g8596 ( 
.A(n_8081),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_7964),
.B(n_7965),
.Y(n_8597)
);

NOR2xp33_ASAP7_75t_L g8598 ( 
.A(n_8100),
.B(n_4812),
.Y(n_8598)
);

INVx2_ASAP7_75t_L g8599 ( 
.A(n_7979),
.Y(n_8599)
);

NAND2xp5_ASAP7_75t_SL g8600 ( 
.A(n_8001),
.B(n_4813),
.Y(n_8600)
);

CKINVDCx20_ASAP7_75t_R g8601 ( 
.A(n_7977),
.Y(n_8601)
);

NAND2xp5_ASAP7_75t_SL g8602 ( 
.A(n_8128),
.B(n_4814),
.Y(n_8602)
);

NAND2xp5_ASAP7_75t_L g8603 ( 
.A(n_7966),
.B(n_4816),
.Y(n_8603)
);

AND2x2_ASAP7_75t_L g8604 ( 
.A(n_7898),
.B(n_4818),
.Y(n_8604)
);

INVx2_ASAP7_75t_L g8605 ( 
.A(n_7989),
.Y(n_8605)
);

INVx5_ASAP7_75t_L g8606 ( 
.A(n_7982),
.Y(n_8606)
);

NAND2xp5_ASAP7_75t_L g8607 ( 
.A(n_7971),
.B(n_4821),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_7999),
.Y(n_8608)
);

AOI21xp5_ASAP7_75t_L g8609 ( 
.A1(n_8103),
.A2(n_3419),
.B(n_3418),
.Y(n_8609)
);

NAND2xp5_ASAP7_75t_L g8610 ( 
.A(n_8000),
.B(n_4822),
.Y(n_8610)
);

AND2x2_ASAP7_75t_L g8611 ( 
.A(n_7987),
.B(n_4824),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_8007),
.Y(n_8612)
);

OAI22xp33_ASAP7_75t_L g8613 ( 
.A1(n_7930),
.A2(n_4827),
.B1(n_4828),
.B2(n_4825),
.Y(n_8613)
);

INVx3_ASAP7_75t_L g8614 ( 
.A(n_8114),
.Y(n_8614)
);

NAND2xp5_ASAP7_75t_L g8615 ( 
.A(n_8004),
.B(n_4830),
.Y(n_8615)
);

NAND2xp5_ASAP7_75t_L g8616 ( 
.A(n_8008),
.B(n_4831),
.Y(n_8616)
);

NOR2xp67_ASAP7_75t_L g8617 ( 
.A(n_8154),
.B(n_3420),
.Y(n_8617)
);

NAND2xp5_ASAP7_75t_L g8618 ( 
.A(n_8013),
.B(n_4832),
.Y(n_8618)
);

AOI221xp5_ASAP7_75t_L g8619 ( 
.A1(n_7931),
.A2(n_4838),
.B1(n_4841),
.B2(n_4837),
.C(n_4834),
.Y(n_8619)
);

NAND2xp5_ASAP7_75t_L g8620 ( 
.A(n_8014),
.B(n_8015),
.Y(n_8620)
);

NAND2xp5_ASAP7_75t_SL g8621 ( 
.A(n_8155),
.B(n_4842),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_8070),
.Y(n_8622)
);

NOR2xp33_ASAP7_75t_L g8623 ( 
.A(n_8073),
.B(n_4845),
.Y(n_8623)
);

OAI21xp5_ASAP7_75t_L g8624 ( 
.A1(n_8034),
.A2(n_4853),
.B(n_4850),
.Y(n_8624)
);

NAND2xp5_ASAP7_75t_L g8625 ( 
.A(n_7982),
.B(n_4856),
.Y(n_8625)
);

INVx2_ASAP7_75t_L g8626 ( 
.A(n_8074),
.Y(n_8626)
);

NAND2xp5_ASAP7_75t_L g8627 ( 
.A(n_8076),
.B(n_4857),
.Y(n_8627)
);

A2O1A1Ixp33_ASAP7_75t_L g8628 ( 
.A1(n_8133),
.A2(n_4862),
.B(n_4864),
.C(n_4858),
.Y(n_8628)
);

AOI221xp5_ASAP7_75t_L g8629 ( 
.A1(n_8105),
.A2(n_4870),
.B1(n_4873),
.B2(n_4867),
.C(n_4865),
.Y(n_8629)
);

BUFx3_ASAP7_75t_L g8630 ( 
.A(n_8173),
.Y(n_8630)
);

INVx2_ASAP7_75t_L g8631 ( 
.A(n_8077),
.Y(n_8631)
);

NAND2xp5_ASAP7_75t_L g8632 ( 
.A(n_8079),
.B(n_4874),
.Y(n_8632)
);

INVx2_ASAP7_75t_L g8633 ( 
.A(n_8080),
.Y(n_8633)
);

NAND2xp33_ASAP7_75t_SL g8634 ( 
.A(n_7961),
.B(n_4876),
.Y(n_8634)
);

NAND2xp5_ASAP7_75t_L g8635 ( 
.A(n_8085),
.B(n_4882),
.Y(n_8635)
);

NAND2xp5_ASAP7_75t_SL g8636 ( 
.A(n_8157),
.B(n_4883),
.Y(n_8636)
);

AND2x6_ASAP7_75t_SL g8637 ( 
.A(n_8170),
.B(n_4884),
.Y(n_8637)
);

OAI221xp5_ASAP7_75t_L g8638 ( 
.A1(n_8049),
.A2(n_4889),
.B1(n_4897),
.B2(n_4886),
.C(n_4885),
.Y(n_8638)
);

NAND2xp5_ASAP7_75t_L g8639 ( 
.A(n_8184),
.B(n_4900),
.Y(n_8639)
);

INVx2_ASAP7_75t_L g8640 ( 
.A(n_7781),
.Y(n_8640)
);

NAND2xp5_ASAP7_75t_L g8641 ( 
.A(n_8095),
.B(n_4901),
.Y(n_8641)
);

NAND2xp5_ASAP7_75t_L g8642 ( 
.A(n_8139),
.B(n_4905),
.Y(n_8642)
);

OAI22xp5_ASAP7_75t_L g8643 ( 
.A1(n_8149),
.A2(n_4911),
.B1(n_4912),
.B2(n_4906),
.Y(n_8643)
);

NOR2xp33_ASAP7_75t_L g8644 ( 
.A(n_7787),
.B(n_4913),
.Y(n_8644)
);

OR2x6_ASAP7_75t_L g8645 ( 
.A(n_7749),
.B(n_3421),
.Y(n_8645)
);

INVx3_ASAP7_75t_L g8646 ( 
.A(n_8176),
.Y(n_8646)
);

AOI22x1_ASAP7_75t_L g8647 ( 
.A1(n_8150),
.A2(n_4923),
.B1(n_4925),
.B2(n_4922),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8067),
.Y(n_8648)
);

AOI22xp33_ASAP7_75t_L g8649 ( 
.A1(n_7994),
.A2(n_4928),
.B1(n_4931),
.B2(n_4927),
.Y(n_8649)
);

NAND2xp5_ASAP7_75t_L g8650 ( 
.A(n_7775),
.B(n_4933),
.Y(n_8650)
);

HB1xp67_ASAP7_75t_L g8651 ( 
.A(n_8179),
.Y(n_8651)
);

NOR2xp33_ASAP7_75t_L g8652 ( 
.A(n_8180),
.B(n_4935),
.Y(n_8652)
);

NAND2xp5_ASAP7_75t_L g8653 ( 
.A(n_8182),
.B(n_4938),
.Y(n_8653)
);

INVx1_ASAP7_75t_L g8654 ( 
.A(n_8183),
.Y(n_8654)
);

AOI22xp33_ASAP7_75t_L g8655 ( 
.A1(n_8185),
.A2(n_4940),
.B1(n_4943),
.B2(n_4939),
.Y(n_8655)
);

INVx2_ASAP7_75t_L g8656 ( 
.A(n_8021),
.Y(n_8656)
);

INVx1_ASAP7_75t_L g8657 ( 
.A(n_8187),
.Y(n_8657)
);

NAND3xp33_ASAP7_75t_L g8658 ( 
.A(n_7949),
.B(n_4947),
.C(n_4946),
.Y(n_8658)
);

NOR2xp33_ASAP7_75t_SL g8659 ( 
.A(n_7883),
.B(n_4948),
.Y(n_8659)
);

NOR2xp33_ASAP7_75t_L g8660 ( 
.A(n_8189),
.B(n_4950),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_8032),
.Y(n_8661)
);

INVx2_ASAP7_75t_L g8662 ( 
.A(n_8146),
.Y(n_8662)
);

INVx2_ASAP7_75t_SL g8663 ( 
.A(n_8193),
.Y(n_8663)
);

NAND2xp5_ASAP7_75t_SL g8664 ( 
.A(n_7996),
.B(n_4951),
.Y(n_8664)
);

INVx2_ASAP7_75t_SL g8665 ( 
.A(n_8116),
.Y(n_8665)
);

NAND2xp5_ASAP7_75t_L g8666 ( 
.A(n_8091),
.B(n_4952),
.Y(n_8666)
);

NAND2xp5_ASAP7_75t_L g8667 ( 
.A(n_7970),
.B(n_7847),
.Y(n_8667)
);

A2O1A1Ixp33_ASAP7_75t_L g8668 ( 
.A1(n_8009),
.A2(n_4958),
.B(n_4959),
.C(n_4957),
.Y(n_8668)
);

NOR2xp33_ASAP7_75t_L g8669 ( 
.A(n_7870),
.B(n_4960),
.Y(n_8669)
);

NAND2xp5_ASAP7_75t_SL g8670 ( 
.A(n_8116),
.B(n_4963),
.Y(n_8670)
);

NAND2xp5_ASAP7_75t_L g8671 ( 
.A(n_8172),
.B(n_4965),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_7975),
.Y(n_8672)
);

AND2x2_ASAP7_75t_L g8673 ( 
.A(n_8159),
.B(n_4966),
.Y(n_8673)
);

NAND2xp5_ASAP7_75t_L g8674 ( 
.A(n_7755),
.B(n_4967),
.Y(n_8674)
);

OAI22xp33_ASAP7_75t_L g8675 ( 
.A1(n_7723),
.A2(n_4969),
.B1(n_4972),
.B2(n_4968),
.Y(n_8675)
);

OR2x6_ASAP7_75t_L g8676 ( 
.A(n_7714),
.B(n_3422),
.Y(n_8676)
);

NAND2xp5_ASAP7_75t_L g8677 ( 
.A(n_7755),
.B(n_4973),
.Y(n_8677)
);

NOR2xp33_ASAP7_75t_L g8678 ( 
.A(n_7723),
.B(n_4974),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_7755),
.B(n_4975),
.Y(n_8679)
);

NAND2xp5_ASAP7_75t_L g8680 ( 
.A(n_7755),
.B(n_4976),
.Y(n_8680)
);

AND2x2_ASAP7_75t_L g8681 ( 
.A(n_7715),
.B(n_8),
.Y(n_8681)
);

A2O1A1Ixp33_ASAP7_75t_L g8682 ( 
.A1(n_7755),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_8682)
);

NAND2xp5_ASAP7_75t_L g8683 ( 
.A(n_7755),
.B(n_9),
.Y(n_8683)
);

NAND2xp5_ASAP7_75t_L g8684 ( 
.A(n_7755),
.B(n_10),
.Y(n_8684)
);

NAND2xp5_ASAP7_75t_L g8685 ( 
.A(n_7755),
.B(n_11),
.Y(n_8685)
);

BUFx3_ASAP7_75t_L g8686 ( 
.A(n_8102),
.Y(n_8686)
);

NOR2xp33_ASAP7_75t_L g8687 ( 
.A(n_7723),
.B(n_11),
.Y(n_8687)
);

INVx1_ASAP7_75t_L g8688 ( 
.A(n_7684),
.Y(n_8688)
);

INVx3_ASAP7_75t_L g8689 ( 
.A(n_7884),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_7684),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_L g8691 ( 
.A(n_7755),
.B(n_12),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_7684),
.Y(n_8692)
);

INVxp67_ASAP7_75t_L g8693 ( 
.A(n_7691),
.Y(n_8693)
);

AOI22xp33_ASAP7_75t_L g8694 ( 
.A1(n_7755),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_8694)
);

NOR2xp33_ASAP7_75t_L g8695 ( 
.A(n_7723),
.B(n_13),
.Y(n_8695)
);

NAND2xp5_ASAP7_75t_L g8696 ( 
.A(n_7755),
.B(n_15),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_7684),
.Y(n_8697)
);

INVx1_ASAP7_75t_L g8698 ( 
.A(n_7684),
.Y(n_8698)
);

INVx2_ASAP7_75t_L g8699 ( 
.A(n_7684),
.Y(n_8699)
);

BUFx3_ASAP7_75t_L g8700 ( 
.A(n_8102),
.Y(n_8700)
);

NAND2xp5_ASAP7_75t_L g8701 ( 
.A(n_7755),
.B(n_16),
.Y(n_8701)
);

AOI21xp5_ASAP7_75t_L g8702 ( 
.A1(n_7804),
.A2(n_3424),
.B(n_3423),
.Y(n_8702)
);

A2O1A1Ixp33_ASAP7_75t_L g8703 ( 
.A1(n_7755),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_8703)
);

NAND2xp5_ASAP7_75t_SL g8704 ( 
.A(n_7723),
.B(n_17),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_7684),
.Y(n_8705)
);

INVx1_ASAP7_75t_L g8706 ( 
.A(n_7684),
.Y(n_8706)
);

INVx2_ASAP7_75t_L g8707 ( 
.A(n_7684),
.Y(n_8707)
);

AND2x4_ASAP7_75t_L g8708 ( 
.A(n_8223),
.B(n_3426),
.Y(n_8708)
);

INVx2_ASAP7_75t_L g8709 ( 
.A(n_8201),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_8378),
.Y(n_8710)
);

INVx2_ASAP7_75t_L g8711 ( 
.A(n_8207),
.Y(n_8711)
);

O2A1O1Ixp33_ASAP7_75t_L g8712 ( 
.A1(n_8259),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_8712)
);

NAND2xp5_ASAP7_75t_L g8713 ( 
.A(n_8237),
.B(n_8240),
.Y(n_8713)
);

INVx2_ASAP7_75t_L g8714 ( 
.A(n_8219),
.Y(n_8714)
);

CKINVDCx5p33_ASAP7_75t_R g8715 ( 
.A(n_8459),
.Y(n_8715)
);

BUFx3_ASAP7_75t_L g8716 ( 
.A(n_8205),
.Y(n_8716)
);

AND2x4_ASAP7_75t_L g8717 ( 
.A(n_8225),
.B(n_3428),
.Y(n_8717)
);

INVx1_ASAP7_75t_L g8718 ( 
.A(n_8473),
.Y(n_8718)
);

A2O1A1Ixp33_ASAP7_75t_L g8719 ( 
.A1(n_8300),
.A2(n_8413),
.B(n_8442),
.C(n_8487),
.Y(n_8719)
);

INVxp67_ASAP7_75t_SL g8720 ( 
.A(n_8291),
.Y(n_8720)
);

INVx2_ASAP7_75t_SL g8721 ( 
.A(n_8390),
.Y(n_8721)
);

BUFx6f_ASAP7_75t_L g8722 ( 
.A(n_8205),
.Y(n_8722)
);

OR2x2_ASAP7_75t_L g8723 ( 
.A(n_8264),
.B(n_19),
.Y(n_8723)
);

INVx2_ASAP7_75t_L g8724 ( 
.A(n_8222),
.Y(n_8724)
);

AOI22xp5_ASAP7_75t_L g8725 ( 
.A1(n_8423),
.A2(n_8286),
.B1(n_8302),
.B2(n_8260),
.Y(n_8725)
);

NAND2xp5_ASAP7_75t_L g8726 ( 
.A(n_8209),
.B(n_20),
.Y(n_8726)
);

INVx2_ASAP7_75t_L g8727 ( 
.A(n_8233),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_8503),
.Y(n_8728)
);

BUFx3_ASAP7_75t_L g8729 ( 
.A(n_8236),
.Y(n_8729)
);

NAND2xp5_ASAP7_75t_L g8730 ( 
.A(n_8195),
.B(n_21),
.Y(n_8730)
);

AOI22xp33_ASAP7_75t_L g8731 ( 
.A1(n_8214),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_8731)
);

HB1xp67_ASAP7_75t_L g8732 ( 
.A(n_8216),
.Y(n_8732)
);

BUFx3_ASAP7_75t_L g8733 ( 
.A(n_8236),
.Y(n_8733)
);

NAND2xp5_ASAP7_75t_SL g8734 ( 
.A(n_8204),
.B(n_23),
.Y(n_8734)
);

BUFx6f_ASAP7_75t_L g8735 ( 
.A(n_8347),
.Y(n_8735)
);

BUFx3_ASAP7_75t_L g8736 ( 
.A(n_8689),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_8239),
.Y(n_8737)
);

NOR2xp33_ASAP7_75t_L g8738 ( 
.A(n_8310),
.B(n_3429),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_SL g8739 ( 
.A(n_8249),
.B(n_24),
.Y(n_8739)
);

INVx2_ASAP7_75t_L g8740 ( 
.A(n_8246),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_L g8741 ( 
.A(n_8678),
.B(n_8674),
.Y(n_8741)
);

NAND2xp5_ASAP7_75t_SL g8742 ( 
.A(n_8197),
.B(n_25),
.Y(n_8742)
);

AOI22xp33_ASAP7_75t_L g8743 ( 
.A1(n_8687),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_8743)
);

INVx1_ASAP7_75t_L g8744 ( 
.A(n_8247),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_L g8745 ( 
.A(n_8677),
.B(n_28),
.Y(n_8745)
);

AOI22xp33_ASAP7_75t_SL g8746 ( 
.A1(n_8695),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_8746)
);

NOR2xp33_ASAP7_75t_L g8747 ( 
.A(n_8316),
.B(n_8639),
.Y(n_8747)
);

NAND2xp5_ASAP7_75t_L g8748 ( 
.A(n_8679),
.B(n_29),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_8294),
.Y(n_8749)
);

INVx2_ASAP7_75t_SL g8750 ( 
.A(n_8390),
.Y(n_8750)
);

NAND2xp5_ASAP7_75t_L g8751 ( 
.A(n_8680),
.B(n_30),
.Y(n_8751)
);

AND2x2_ASAP7_75t_L g8752 ( 
.A(n_8336),
.B(n_31),
.Y(n_8752)
);

INVx2_ASAP7_75t_L g8753 ( 
.A(n_8307),
.Y(n_8753)
);

HB1xp67_ASAP7_75t_L g8754 ( 
.A(n_8458),
.Y(n_8754)
);

INVx3_ASAP7_75t_L g8755 ( 
.A(n_8384),
.Y(n_8755)
);

NAND2xp5_ASAP7_75t_L g8756 ( 
.A(n_8279),
.B(n_32),
.Y(n_8756)
);

INVx2_ASAP7_75t_L g8757 ( 
.A(n_8311),
.Y(n_8757)
);

INVxp67_ASAP7_75t_L g8758 ( 
.A(n_8462),
.Y(n_8758)
);

NAND2xp5_ASAP7_75t_L g8759 ( 
.A(n_8270),
.B(n_32),
.Y(n_8759)
);

INVx3_ASAP7_75t_L g8760 ( 
.A(n_8384),
.Y(n_8760)
);

INVx1_ASAP7_75t_L g8761 ( 
.A(n_8313),
.Y(n_8761)
);

AND2x2_ASAP7_75t_SL g8762 ( 
.A(n_8694),
.B(n_33),
.Y(n_8762)
);

OR2x6_ASAP7_75t_L g8763 ( 
.A(n_8348),
.B(n_3431),
.Y(n_8763)
);

AND2x4_ASAP7_75t_L g8764 ( 
.A(n_8403),
.B(n_3432),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_SL g8765 ( 
.A(n_8230),
.B(n_33),
.Y(n_8765)
);

NAND2xp5_ASAP7_75t_L g8766 ( 
.A(n_8213),
.B(n_35),
.Y(n_8766)
);

NAND2xp5_ASAP7_75t_L g8767 ( 
.A(n_8215),
.B(n_8273),
.Y(n_8767)
);

NAND2xp5_ASAP7_75t_SL g8768 ( 
.A(n_8445),
.B(n_35),
.Y(n_8768)
);

BUFx3_ASAP7_75t_L g8769 ( 
.A(n_8348),
.Y(n_8769)
);

OR2x6_ASAP7_75t_L g8770 ( 
.A(n_8227),
.B(n_3433),
.Y(n_8770)
);

AND2x6_ASAP7_75t_SL g8771 ( 
.A(n_8644),
.B(n_36),
.Y(n_8771)
);

INVx2_ASAP7_75t_L g8772 ( 
.A(n_8328),
.Y(n_8772)
);

OAI21xp33_ASAP7_75t_L g8773 ( 
.A1(n_8292),
.A2(n_36),
.B(n_37),
.Y(n_8773)
);

INVx4_ASAP7_75t_L g8774 ( 
.A(n_8419),
.Y(n_8774)
);

INVx3_ASAP7_75t_L g8775 ( 
.A(n_8419),
.Y(n_8775)
);

AND2x2_ASAP7_75t_L g8776 ( 
.A(n_8681),
.B(n_37),
.Y(n_8776)
);

AOI22xp5_ASAP7_75t_L g8777 ( 
.A1(n_8475),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_8777)
);

AND2x2_ASAP7_75t_L g8778 ( 
.A(n_8194),
.B(n_38),
.Y(n_8778)
);

INVx2_ASAP7_75t_L g8779 ( 
.A(n_8329),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_SL g8780 ( 
.A(n_8211),
.B(n_41),
.Y(n_8780)
);

INVx2_ASAP7_75t_SL g8781 ( 
.A(n_8361),
.Y(n_8781)
);

INVx2_ASAP7_75t_L g8782 ( 
.A(n_8331),
.Y(n_8782)
);

BUFx3_ASAP7_75t_L g8783 ( 
.A(n_8589),
.Y(n_8783)
);

AND2x2_ASAP7_75t_L g8784 ( 
.A(n_8565),
.B(n_42),
.Y(n_8784)
);

INVx1_ASAP7_75t_L g8785 ( 
.A(n_8375),
.Y(n_8785)
);

NAND2xp5_ASAP7_75t_L g8786 ( 
.A(n_8200),
.B(n_44),
.Y(n_8786)
);

BUFx6f_ASAP7_75t_L g8787 ( 
.A(n_8541),
.Y(n_8787)
);

OAI22xp33_ASAP7_75t_L g8788 ( 
.A1(n_8548),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_8788)
);

NAND2xp5_ASAP7_75t_L g8789 ( 
.A(n_8596),
.B(n_45),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_8683),
.B(n_46),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_8399),
.Y(n_8791)
);

INVx1_ASAP7_75t_SL g8792 ( 
.A(n_8301),
.Y(n_8792)
);

INVx1_ASAP7_75t_L g8793 ( 
.A(n_8401),
.Y(n_8793)
);

NAND2xp5_ASAP7_75t_L g8794 ( 
.A(n_8684),
.B(n_47),
.Y(n_8794)
);

NOR3xp33_ASAP7_75t_SL g8795 ( 
.A(n_8226),
.B(n_48),
.C(n_49),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_SL g8796 ( 
.A(n_8196),
.B(n_48),
.Y(n_8796)
);

CKINVDCx5p33_ASAP7_75t_R g8797 ( 
.A(n_8524),
.Y(n_8797)
);

NAND2xp5_ASAP7_75t_L g8798 ( 
.A(n_8685),
.B(n_49),
.Y(n_8798)
);

HB1xp67_ASAP7_75t_L g8799 ( 
.A(n_8212),
.Y(n_8799)
);

NAND2xp5_ASAP7_75t_L g8800 ( 
.A(n_8691),
.B(n_50),
.Y(n_8800)
);

INVx1_ASAP7_75t_L g8801 ( 
.A(n_8415),
.Y(n_8801)
);

INVx2_ASAP7_75t_L g8802 ( 
.A(n_8418),
.Y(n_8802)
);

INVx2_ASAP7_75t_L g8803 ( 
.A(n_8433),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_8443),
.Y(n_8804)
);

INVx2_ASAP7_75t_SL g8805 ( 
.A(n_8202),
.Y(n_8805)
);

AND2x4_ASAP7_75t_L g8806 ( 
.A(n_8337),
.B(n_3435),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_L g8807 ( 
.A(n_8696),
.B(n_50),
.Y(n_8807)
);

NAND3xp33_ASAP7_75t_L g8808 ( 
.A(n_8297),
.B(n_51),
.C(n_52),
.Y(n_8808)
);

INVx2_ASAP7_75t_L g8809 ( 
.A(n_8464),
.Y(n_8809)
);

NAND2xp5_ASAP7_75t_L g8810 ( 
.A(n_8701),
.B(n_52),
.Y(n_8810)
);

INVx3_ASAP7_75t_L g8811 ( 
.A(n_8314),
.Y(n_8811)
);

NAND2xp5_ASAP7_75t_L g8812 ( 
.A(n_8304),
.B(n_8305),
.Y(n_8812)
);

NOR2xp33_ASAP7_75t_L g8813 ( 
.A(n_8641),
.B(n_3437),
.Y(n_8813)
);

AO22x1_ASAP7_75t_L g8814 ( 
.A1(n_8606),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8466),
.Y(n_8815)
);

NAND2xp5_ASAP7_75t_SL g8816 ( 
.A(n_8248),
.B(n_53),
.Y(n_8816)
);

INVx4_ASAP7_75t_L g8817 ( 
.A(n_8224),
.Y(n_8817)
);

NAND2xp5_ASAP7_75t_L g8818 ( 
.A(n_8360),
.B(n_54),
.Y(n_8818)
);

OR2x2_ASAP7_75t_L g8819 ( 
.A(n_8272),
.B(n_56),
.Y(n_8819)
);

INVx1_ASAP7_75t_L g8820 ( 
.A(n_8472),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_L g8821 ( 
.A(n_8414),
.B(n_56),
.Y(n_8821)
);

NAND2xp5_ASAP7_75t_SL g8822 ( 
.A(n_8525),
.B(n_58),
.Y(n_8822)
);

INVx1_ASAP7_75t_L g8823 ( 
.A(n_8474),
.Y(n_8823)
);

OR2x4_ASAP7_75t_L g8824 ( 
.A(n_8243),
.B(n_59),
.Y(n_8824)
);

INVx1_ASAP7_75t_L g8825 ( 
.A(n_8479),
.Y(n_8825)
);

HB1xp67_ASAP7_75t_L g8826 ( 
.A(n_8693),
.Y(n_8826)
);

NAND2xp5_ASAP7_75t_SL g8827 ( 
.A(n_8218),
.B(n_60),
.Y(n_8827)
);

NAND2xp5_ASAP7_75t_L g8828 ( 
.A(n_8467),
.B(n_60),
.Y(n_8828)
);

AND2x2_ASAP7_75t_L g8829 ( 
.A(n_8388),
.B(n_8570),
.Y(n_8829)
);

NAND2xp5_ASAP7_75t_L g8830 ( 
.A(n_8480),
.B(n_61),
.Y(n_8830)
);

INVx2_ASAP7_75t_L g8831 ( 
.A(n_8481),
.Y(n_8831)
);

NAND2xp5_ASAP7_75t_L g8832 ( 
.A(n_8250),
.B(n_8251),
.Y(n_8832)
);

NAND2xp5_ASAP7_75t_L g8833 ( 
.A(n_8275),
.B(n_61),
.Y(n_8833)
);

NAND2xp5_ASAP7_75t_SL g8834 ( 
.A(n_8267),
.B(n_62),
.Y(n_8834)
);

OR2x2_ASAP7_75t_SL g8835 ( 
.A(n_8381),
.B(n_63),
.Y(n_8835)
);

NAND2xp5_ASAP7_75t_SL g8836 ( 
.A(n_8203),
.B(n_63),
.Y(n_8836)
);

NOR2xp33_ASAP7_75t_L g8837 ( 
.A(n_8671),
.B(n_8277),
.Y(n_8837)
);

INVx2_ASAP7_75t_L g8838 ( 
.A(n_8692),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_8699),
.Y(n_8839)
);

BUFx12f_ASAP7_75t_L g8840 ( 
.A(n_8381),
.Y(n_8840)
);

AOI22xp33_ASAP7_75t_L g8841 ( 
.A1(n_8263),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_8841)
);

NAND2xp5_ASAP7_75t_SL g8842 ( 
.A(n_8232),
.B(n_64),
.Y(n_8842)
);

NAND2xp5_ASAP7_75t_L g8843 ( 
.A(n_8280),
.B(n_65),
.Y(n_8843)
);

NAND2xp5_ASAP7_75t_L g8844 ( 
.A(n_8282),
.B(n_68),
.Y(n_8844)
);

A2O1A1Ixp33_ASAP7_75t_L g8845 ( 
.A1(n_8542),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_8845)
);

NAND2xp5_ASAP7_75t_SL g8846 ( 
.A(n_8206),
.B(n_71),
.Y(n_8846)
);

OR2x2_ASAP7_75t_L g8847 ( 
.A(n_8320),
.B(n_71),
.Y(n_8847)
);

INVx2_ASAP7_75t_L g8848 ( 
.A(n_8705),
.Y(n_8848)
);

NOR2xp33_ASAP7_75t_R g8849 ( 
.A(n_8315),
.B(n_3439),
.Y(n_8849)
);

NAND2xp5_ASAP7_75t_L g8850 ( 
.A(n_8284),
.B(n_72),
.Y(n_8850)
);

INVx2_ASAP7_75t_L g8851 ( 
.A(n_8707),
.Y(n_8851)
);

INVx2_ASAP7_75t_L g8852 ( 
.A(n_8513),
.Y(n_8852)
);

CKINVDCx5p33_ASAP7_75t_R g8853 ( 
.A(n_8527),
.Y(n_8853)
);

AND2x4_ASAP7_75t_L g8854 ( 
.A(n_8463),
.B(n_3440),
.Y(n_8854)
);

INVx1_ASAP7_75t_L g8855 ( 
.A(n_8199),
.Y(n_8855)
);

BUFx2_ASAP7_75t_L g8856 ( 
.A(n_8245),
.Y(n_8856)
);

AOI22xp5_ASAP7_75t_L g8857 ( 
.A1(n_8392),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_8857)
);

NAND2xp5_ASAP7_75t_L g8858 ( 
.A(n_8288),
.B(n_8235),
.Y(n_8858)
);

INVx1_ASAP7_75t_L g8859 ( 
.A(n_8208),
.Y(n_8859)
);

BUFx8_ASAP7_75t_L g8860 ( 
.A(n_8491),
.Y(n_8860)
);

INVx1_ASAP7_75t_L g8861 ( 
.A(n_8238),
.Y(n_8861)
);

NAND2xp5_ASAP7_75t_SL g8862 ( 
.A(n_8538),
.B(n_73),
.Y(n_8862)
);

INVx1_ASAP7_75t_L g8863 ( 
.A(n_8242),
.Y(n_8863)
);

AND2x4_ASAP7_75t_L g8864 ( 
.A(n_8463),
.B(n_8614),
.Y(n_8864)
);

OR2x6_ASAP7_75t_L g8865 ( 
.A(n_8676),
.B(n_3446),
.Y(n_8865)
);

AOI22xp5_ASAP7_75t_L g8866 ( 
.A1(n_8471),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_8866)
);

NOR2xp67_ASAP7_75t_L g8867 ( 
.A(n_8576),
.B(n_3447),
.Y(n_8867)
);

INVx2_ASAP7_75t_L g8868 ( 
.A(n_8514),
.Y(n_8868)
);

INVx1_ASAP7_75t_L g8869 ( 
.A(n_8244),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_8256),
.Y(n_8870)
);

OR2x6_ASAP7_75t_L g8871 ( 
.A(n_8676),
.B(n_3448),
.Y(n_8871)
);

AND2x6_ASAP7_75t_L g8872 ( 
.A(n_8258),
.B(n_3452),
.Y(n_8872)
);

NOR2xp33_ASAP7_75t_L g8873 ( 
.A(n_8658),
.B(n_3453),
.Y(n_8873)
);

BUFx6f_ASAP7_75t_L g8874 ( 
.A(n_8541),
.Y(n_8874)
);

INVx2_ASAP7_75t_L g8875 ( 
.A(n_8626),
.Y(n_8875)
);

AOI22xp5_ASAP7_75t_L g8876 ( 
.A1(n_8634),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_8876)
);

BUFx6f_ASAP7_75t_L g8877 ( 
.A(n_8581),
.Y(n_8877)
);

OAI22xp5_ASAP7_75t_L g8878 ( 
.A1(n_8455),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_8878)
);

NAND2xp5_ASAP7_75t_L g8879 ( 
.A(n_8341),
.B(n_79),
.Y(n_8879)
);

INVx5_ASAP7_75t_L g8880 ( 
.A(n_8338),
.Y(n_8880)
);

INVx1_ASAP7_75t_L g8881 ( 
.A(n_8274),
.Y(n_8881)
);

INVx2_ASAP7_75t_L g8882 ( 
.A(n_8631),
.Y(n_8882)
);

BUFx3_ASAP7_75t_L g8883 ( 
.A(n_8228),
.Y(n_8883)
);

AOI22xp5_ASAP7_75t_L g8884 ( 
.A1(n_8526),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_8884)
);

INVx2_ASAP7_75t_L g8885 ( 
.A(n_8633),
.Y(n_8885)
);

AND2x2_ASAP7_75t_L g8886 ( 
.A(n_8299),
.B(n_81),
.Y(n_8886)
);

INVx3_ASAP7_75t_L g8887 ( 
.A(n_8367),
.Y(n_8887)
);

INVx2_ASAP7_75t_L g8888 ( 
.A(n_8507),
.Y(n_8888)
);

INVx3_ASAP7_75t_L g8889 ( 
.A(n_8382),
.Y(n_8889)
);

BUFx2_ASAP7_75t_L g8890 ( 
.A(n_8366),
.Y(n_8890)
);

NAND2xp5_ASAP7_75t_L g8891 ( 
.A(n_8358),
.B(n_82),
.Y(n_8891)
);

AND2x4_ASAP7_75t_L g8892 ( 
.A(n_8665),
.B(n_8345),
.Y(n_8892)
);

NAND2xp5_ASAP7_75t_SL g8893 ( 
.A(n_8229),
.B(n_83),
.Y(n_8893)
);

AOI22xp33_ASAP7_75t_L g8894 ( 
.A1(n_8448),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_8894)
);

INVx3_ASAP7_75t_SL g8895 ( 
.A(n_8601),
.Y(n_8895)
);

AND2x4_ASAP7_75t_L g8896 ( 
.A(n_8265),
.B(n_3454),
.Y(n_8896)
);

AND2x4_ASAP7_75t_L g8897 ( 
.A(n_8281),
.B(n_3459),
.Y(n_8897)
);

NAND2xp5_ASAP7_75t_SL g8898 ( 
.A(n_8613),
.B(n_84),
.Y(n_8898)
);

INVx2_ASAP7_75t_L g8899 ( 
.A(n_8517),
.Y(n_8899)
);

INVx4_ASAP7_75t_L g8900 ( 
.A(n_8224),
.Y(n_8900)
);

BUFx4f_ASAP7_75t_L g8901 ( 
.A(n_8581),
.Y(n_8901)
);

INVx1_ASAP7_75t_L g8902 ( 
.A(n_8287),
.Y(n_8902)
);

INVx2_ASAP7_75t_L g8903 ( 
.A(n_8528),
.Y(n_8903)
);

INVx1_ASAP7_75t_L g8904 ( 
.A(n_8289),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8362),
.B(n_86),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_8364),
.B(n_87),
.Y(n_8906)
);

INVx1_ASAP7_75t_SL g8907 ( 
.A(n_8510),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8529),
.Y(n_8908)
);

AND2x4_ASAP7_75t_L g8909 ( 
.A(n_8293),
.B(n_3461),
.Y(n_8909)
);

INVx1_ASAP7_75t_L g8910 ( 
.A(n_8296),
.Y(n_8910)
);

AOI22xp5_ASAP7_75t_L g8911 ( 
.A1(n_8669),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_8911)
);

NOR2xp33_ASAP7_75t_L g8912 ( 
.A(n_8672),
.B(n_3463),
.Y(n_8912)
);

INVx2_ASAP7_75t_SL g8913 ( 
.A(n_8349),
.Y(n_8913)
);

NAND2xp5_ASAP7_75t_L g8914 ( 
.A(n_8368),
.B(n_91),
.Y(n_8914)
);

BUFx10_ASAP7_75t_L g8915 ( 
.A(n_8470),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_SL g8916 ( 
.A(n_8675),
.B(n_92),
.Y(n_8916)
);

INVx2_ASAP7_75t_L g8917 ( 
.A(n_8531),
.Y(n_8917)
);

INVx1_ASAP7_75t_L g8918 ( 
.A(n_8303),
.Y(n_8918)
);

NOR2xp33_ASAP7_75t_L g8919 ( 
.A(n_8673),
.B(n_3464),
.Y(n_8919)
);

INVx2_ASAP7_75t_L g8920 ( 
.A(n_8536),
.Y(n_8920)
);

NAND2x1_ASAP7_75t_L g8921 ( 
.A(n_8656),
.B(n_3465),
.Y(n_8921)
);

NAND2xp5_ASAP7_75t_L g8922 ( 
.A(n_8269),
.B(n_94),
.Y(n_8922)
);

INVx3_ASAP7_75t_L g8923 ( 
.A(n_8407),
.Y(n_8923)
);

INVx4_ASAP7_75t_L g8924 ( 
.A(n_8262),
.Y(n_8924)
);

INVx3_ASAP7_75t_L g8925 ( 
.A(n_8396),
.Y(n_8925)
);

AOI22xp33_ASAP7_75t_L g8926 ( 
.A1(n_8564),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_8926)
);

AOI22xp33_ASAP7_75t_L g8927 ( 
.A1(n_8704),
.A2(n_8624),
.B1(n_8395),
.B2(n_8332),
.Y(n_8927)
);

AND2x4_ASAP7_75t_L g8928 ( 
.A(n_8356),
.B(n_3466),
.Y(n_8928)
);

NOR2xp33_ASAP7_75t_L g8929 ( 
.A(n_8530),
.B(n_3468),
.Y(n_8929)
);

OR2x6_ASAP7_75t_L g8930 ( 
.A(n_8198),
.B(n_3469),
.Y(n_8930)
);

A2O1A1Ixp33_ASAP7_75t_L g8931 ( 
.A1(n_8351),
.A2(n_8340),
.B(n_8241),
.C(n_8577),
.Y(n_8931)
);

INVx1_ASAP7_75t_L g8932 ( 
.A(n_8317),
.Y(n_8932)
);

NAND2xp5_ASAP7_75t_L g8933 ( 
.A(n_8271),
.B(n_95),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8318),
.Y(n_8934)
);

BUFx2_ASAP7_75t_L g8935 ( 
.A(n_8532),
.Y(n_8935)
);

INVx2_ASAP7_75t_SL g8936 ( 
.A(n_8357),
.Y(n_8936)
);

AND2x2_ASAP7_75t_L g8937 ( 
.A(n_8309),
.B(n_98),
.Y(n_8937)
);

INVx1_ASAP7_75t_L g8938 ( 
.A(n_8325),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8327),
.Y(n_8939)
);

INVx1_ASAP7_75t_L g8940 ( 
.A(n_8335),
.Y(n_8940)
);

BUFx3_ASAP7_75t_L g8941 ( 
.A(n_8686),
.Y(n_8941)
);

INVx2_ASAP7_75t_L g8942 ( 
.A(n_8556),
.Y(n_8942)
);

CKINVDCx5p33_ASAP7_75t_R g8943 ( 
.A(n_8268),
.Y(n_8943)
);

AND2x6_ASAP7_75t_SL g8944 ( 
.A(n_8450),
.B(n_98),
.Y(n_8944)
);

NOR2xp33_ASAP7_75t_L g8945 ( 
.A(n_8583),
.B(n_3470),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8343),
.Y(n_8946)
);

AO21x1_ASAP7_75t_L g8947 ( 
.A1(n_8210),
.A2(n_99),
.B(n_100),
.Y(n_8947)
);

NAND2xp5_ASAP7_75t_L g8948 ( 
.A(n_8323),
.B(n_99),
.Y(n_8948)
);

AND2x4_ASAP7_75t_L g8949 ( 
.A(n_8346),
.B(n_3471),
.Y(n_8949)
);

INVx2_ASAP7_75t_L g8950 ( 
.A(n_8557),
.Y(n_8950)
);

AOI22xp33_ASAP7_75t_SL g8951 ( 
.A1(n_8220),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_8951)
);

INVx2_ASAP7_75t_SL g8952 ( 
.A(n_8432),
.Y(n_8952)
);

BUFx2_ASAP7_75t_L g8953 ( 
.A(n_8523),
.Y(n_8953)
);

NAND2x1p5_ASAP7_75t_L g8954 ( 
.A(n_8606),
.B(n_3473),
.Y(n_8954)
);

AOI22xp33_ASAP7_75t_L g8955 ( 
.A1(n_8354),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_8955)
);

NAND2xp5_ASAP7_75t_L g8956 ( 
.A(n_8339),
.B(n_104),
.Y(n_8956)
);

NAND2xp5_ASAP7_75t_SL g8957 ( 
.A(n_8254),
.B(n_104),
.Y(n_8957)
);

AND2x2_ASAP7_75t_L g8958 ( 
.A(n_8359),
.B(n_105),
.Y(n_8958)
);

INVxp67_ASAP7_75t_L g8959 ( 
.A(n_8276),
.Y(n_8959)
);

NAND2xp5_ASAP7_75t_SL g8960 ( 
.A(n_8234),
.B(n_105),
.Y(n_8960)
);

NOR2xp33_ASAP7_75t_L g8961 ( 
.A(n_8333),
.B(n_3474),
.Y(n_8961)
);

INVx1_ASAP7_75t_L g8962 ( 
.A(n_8365),
.Y(n_8962)
);

NAND2xp5_ASAP7_75t_SL g8963 ( 
.A(n_8606),
.B(n_106),
.Y(n_8963)
);

INVx1_ASAP7_75t_SL g8964 ( 
.A(n_8255),
.Y(n_8964)
);

OAI21xp33_ASAP7_75t_L g8965 ( 
.A1(n_8321),
.A2(n_8533),
.B(n_8537),
.Y(n_8965)
);

CKINVDCx8_ASAP7_75t_R g8966 ( 
.A(n_8637),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_8386),
.B(n_106),
.Y(n_8967)
);

OR2x6_ASAP7_75t_L g8968 ( 
.A(n_8450),
.B(n_8700),
.Y(n_8968)
);

INVx2_ASAP7_75t_L g8969 ( 
.A(n_8560),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_8369),
.Y(n_8970)
);

AOI22xp33_ASAP7_75t_L g8971 ( 
.A1(n_8546),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_8971)
);

HB1xp67_ASAP7_75t_L g8972 ( 
.A(n_8588),
.Y(n_8972)
);

CKINVDCx20_ASAP7_75t_R g8973 ( 
.A(n_8387),
.Y(n_8973)
);

NAND2xp5_ASAP7_75t_L g8974 ( 
.A(n_8285),
.B(n_8324),
.Y(n_8974)
);

AND2x2_ASAP7_75t_L g8975 ( 
.A(n_8604),
.B(n_108),
.Y(n_8975)
);

INVx1_ASAP7_75t_SL g8976 ( 
.A(n_8231),
.Y(n_8976)
);

NAND2xp5_ASAP7_75t_L g8977 ( 
.A(n_8444),
.B(n_110),
.Y(n_8977)
);

INVx1_ASAP7_75t_SL g8978 ( 
.A(n_8630),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_8373),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_8389),
.Y(n_8980)
);

INVx2_ASAP7_75t_L g8981 ( 
.A(n_8569),
.Y(n_8981)
);

NAND2xp5_ASAP7_75t_SL g8982 ( 
.A(n_8416),
.B(n_110),
.Y(n_8982)
);

BUFx6f_ASAP7_75t_L g8983 ( 
.A(n_8338),
.Y(n_8983)
);

INVx5_ASAP7_75t_L g8984 ( 
.A(n_8645),
.Y(n_8984)
);

INVx1_ASAP7_75t_L g8985 ( 
.A(n_8393),
.Y(n_8985)
);

NAND2xp5_ASAP7_75t_L g8986 ( 
.A(n_8520),
.B(n_111),
.Y(n_8986)
);

INVx1_ASAP7_75t_L g8987 ( 
.A(n_8404),
.Y(n_8987)
);

INVx2_ASAP7_75t_L g8988 ( 
.A(n_8584),
.Y(n_8988)
);

NOR2xp33_ASAP7_75t_L g8989 ( 
.A(n_8667),
.B(n_3475),
.Y(n_8989)
);

INVx2_ASAP7_75t_L g8990 ( 
.A(n_8587),
.Y(n_8990)
);

OR2x6_ASAP7_75t_L g8991 ( 
.A(n_8645),
.B(n_3477),
.Y(n_8991)
);

NAND2xp5_ASAP7_75t_SL g8992 ( 
.A(n_8509),
.B(n_111),
.Y(n_8992)
);

NAND2xp5_ASAP7_75t_L g8993 ( 
.A(n_8623),
.B(n_112),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8599),
.Y(n_8994)
);

NAND2xp5_ASAP7_75t_L g8995 ( 
.A(n_8611),
.B(n_112),
.Y(n_8995)
);

OAI21xp5_ASAP7_75t_L g8996 ( 
.A1(n_8344),
.A2(n_113),
.B(n_114),
.Y(n_8996)
);

AOI22xp33_ASAP7_75t_L g8997 ( 
.A1(n_8295),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_8408),
.Y(n_8998)
);

NAND2xp5_ASAP7_75t_SL g8999 ( 
.A(n_8659),
.B(n_115),
.Y(n_8999)
);

INVx2_ASAP7_75t_L g9000 ( 
.A(n_8605),
.Y(n_9000)
);

NAND2xp33_ASAP7_75t_SL g9001 ( 
.A(n_8363),
.B(n_116),
.Y(n_9001)
);

NAND2xp5_ASAP7_75t_L g9002 ( 
.A(n_8319),
.B(n_117),
.Y(n_9002)
);

NAND2xp5_ASAP7_75t_L g9003 ( 
.A(n_8593),
.B(n_117),
.Y(n_9003)
);

CKINVDCx5p33_ASAP7_75t_R g9004 ( 
.A(n_8457),
.Y(n_9004)
);

BUFx3_ASAP7_75t_L g9005 ( 
.A(n_8519),
.Y(n_9005)
);

AOI22xp5_ASAP7_75t_L g9006 ( 
.A1(n_8485),
.A2(n_8253),
.B1(n_8330),
.B2(n_8497),
.Y(n_9006)
);

NOR2xp33_ASAP7_75t_L g9007 ( 
.A(n_8261),
.B(n_3478),
.Y(n_9007)
);

NAND2xp5_ASAP7_75t_L g9008 ( 
.A(n_8594),
.B(n_119),
.Y(n_9008)
);

BUFx6f_ASAP7_75t_L g9009 ( 
.A(n_8551),
.Y(n_9009)
);

INVx1_ASAP7_75t_SL g9010 ( 
.A(n_8651),
.Y(n_9010)
);

INVx1_ASAP7_75t_L g9011 ( 
.A(n_8424),
.Y(n_9011)
);

NOR2xp33_ASAP7_75t_L g9012 ( 
.A(n_8638),
.B(n_3481),
.Y(n_9012)
);

NAND2xp5_ASAP7_75t_L g9013 ( 
.A(n_8598),
.B(n_120),
.Y(n_9013)
);

BUFx8_ASAP7_75t_L g9014 ( 
.A(n_8654),
.Y(n_9014)
);

AOI21xp33_ASAP7_75t_L g9015 ( 
.A1(n_8278),
.A2(n_120),
.B(n_121),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_8429),
.Y(n_9016)
);

NAND3xp33_ASAP7_75t_SL g9017 ( 
.A(n_8649),
.B(n_121),
.C(n_122),
.Y(n_9017)
);

OAI22xp5_ASAP7_75t_L g9018 ( 
.A1(n_8586),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_9018)
);

NAND2xp5_ASAP7_75t_SL g9019 ( 
.A(n_8535),
.B(n_8426),
.Y(n_9019)
);

AOI22xp5_ASAP7_75t_L g9020 ( 
.A1(n_8453),
.A2(n_8494),
.B1(n_8355),
.B2(n_8476),
.Y(n_9020)
);

INVx1_ASAP7_75t_L g9021 ( 
.A(n_8430),
.Y(n_9021)
);

INVx1_ASAP7_75t_L g9022 ( 
.A(n_8435),
.Y(n_9022)
);

NOR2xp33_ASAP7_75t_L g9023 ( 
.A(n_8508),
.B(n_3482),
.Y(n_9023)
);

NAND2xp5_ASAP7_75t_L g9024 ( 
.A(n_8431),
.B(n_123),
.Y(n_9024)
);

NAND2xp5_ASAP7_75t_SL g9025 ( 
.A(n_8446),
.B(n_124),
.Y(n_9025)
);

INVx1_ASAP7_75t_L g9026 ( 
.A(n_8438),
.Y(n_9026)
);

AND2x2_ASAP7_75t_L g9027 ( 
.A(n_8483),
.B(n_125),
.Y(n_9027)
);

BUFx2_ASAP7_75t_L g9028 ( 
.A(n_8646),
.Y(n_9028)
);

AOI22xp5_ASAP7_75t_L g9029 ( 
.A1(n_8374),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_9029)
);

BUFx6f_ASAP7_75t_L g9030 ( 
.A(n_8582),
.Y(n_9030)
);

OR2x4_ASAP7_75t_L g9031 ( 
.A(n_8555),
.B(n_8561),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8440),
.Y(n_9032)
);

NOR3xp33_ASAP7_75t_SL g9033 ( 
.A(n_8283),
.B(n_128),
.C(n_129),
.Y(n_9033)
);

OR2x2_ASAP7_75t_L g9034 ( 
.A(n_8447),
.B(n_128),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_L g9035 ( 
.A(n_8308),
.B(n_130),
.Y(n_9035)
);

INVxp67_ASAP7_75t_L g9036 ( 
.A(n_8568),
.Y(n_9036)
);

OAI22xp5_ASAP7_75t_L g9037 ( 
.A1(n_8217),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_9037)
);

AND2x6_ASAP7_75t_SL g9038 ( 
.A(n_8406),
.B(n_131),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8451),
.Y(n_9039)
);

BUFx12f_ASAP7_75t_L g9040 ( 
.A(n_8298),
.Y(n_9040)
);

NAND2xp5_ASAP7_75t_L g9041 ( 
.A(n_8482),
.B(n_134),
.Y(n_9041)
);

INVx1_ASAP7_75t_L g9042 ( 
.A(n_8461),
.Y(n_9042)
);

INVxp67_ASAP7_75t_SL g9043 ( 
.A(n_8549),
.Y(n_9043)
);

AOI22xp33_ASAP7_75t_L g9044 ( 
.A1(n_8629),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_8688),
.Y(n_9045)
);

CKINVDCx5p33_ASAP7_75t_R g9046 ( 
.A(n_8406),
.Y(n_9046)
);

NAND2xp5_ASAP7_75t_SL g9047 ( 
.A(n_8552),
.B(n_135),
.Y(n_9047)
);

O2A1O1Ixp33_ASAP7_75t_L g9048 ( 
.A1(n_8682),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_9048)
);

NAND2xp5_ASAP7_75t_L g9049 ( 
.A(n_8500),
.B(n_137),
.Y(n_9049)
);

OAI22xp5_ASAP7_75t_SL g9050 ( 
.A1(n_8334),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_9050)
);

NAND2xp5_ASAP7_75t_L g9051 ( 
.A(n_8516),
.B(n_139),
.Y(n_9051)
);

NAND2xp5_ASAP7_75t_L g9052 ( 
.A(n_8690),
.B(n_140),
.Y(n_9052)
);

INVx2_ASAP7_75t_L g9053 ( 
.A(n_8697),
.Y(n_9053)
);

BUFx2_ASAP7_75t_L g9054 ( 
.A(n_8663),
.Y(n_9054)
);

BUFx6f_ASAP7_75t_L g9055 ( 
.A(n_8257),
.Y(n_9055)
);

OR2x6_ASAP7_75t_L g9056 ( 
.A(n_8437),
.B(n_8376),
.Y(n_9056)
);

NAND2xp5_ASAP7_75t_L g9057 ( 
.A(n_8698),
.B(n_141),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_8706),
.Y(n_9058)
);

HB1xp67_ASAP7_75t_L g9059 ( 
.A(n_8489),
.Y(n_9059)
);

INVx2_ASAP7_75t_L g9060 ( 
.A(n_8486),
.Y(n_9060)
);

BUFx3_ASAP7_75t_L g9061 ( 
.A(n_8657),
.Y(n_9061)
);

OR2x2_ASAP7_75t_L g9062 ( 
.A(n_8597),
.B(n_8620),
.Y(n_9062)
);

AND2x4_ASAP7_75t_L g9063 ( 
.A(n_8488),
.B(n_3483),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_8493),
.Y(n_9064)
);

NOR2x1p5_ASAP7_75t_L g9065 ( 
.A(n_8625),
.B(n_3485),
.Y(n_9065)
);

NAND2xp5_ASAP7_75t_SL g9066 ( 
.A(n_8290),
.B(n_142),
.Y(n_9066)
);

NOR2x1p5_ASAP7_75t_L g9067 ( 
.A(n_8650),
.B(n_3486),
.Y(n_9067)
);

NAND2xp5_ASAP7_75t_L g9068 ( 
.A(n_8370),
.B(n_142),
.Y(n_9068)
);

NAND2xp5_ASAP7_75t_L g9069 ( 
.A(n_8312),
.B(n_8439),
.Y(n_9069)
);

INVxp67_ASAP7_75t_L g9070 ( 
.A(n_8371),
.Y(n_9070)
);

CKINVDCx5p33_ASAP7_75t_R g9071 ( 
.A(n_8353),
.Y(n_9071)
);

CKINVDCx5p33_ASAP7_75t_R g9072 ( 
.A(n_8670),
.Y(n_9072)
);

CKINVDCx20_ASAP7_75t_R g9073 ( 
.A(n_8505),
.Y(n_9073)
);

BUFx4f_ASAP7_75t_L g9074 ( 
.A(n_8622),
.Y(n_9074)
);

INVx3_ASAP7_75t_L g9075 ( 
.A(n_8495),
.Y(n_9075)
);

INVx2_ASAP7_75t_SL g9076 ( 
.A(n_8221),
.Y(n_9076)
);

OAI22xp5_ASAP7_75t_SL g9077 ( 
.A1(n_8266),
.A2(n_8306),
.B1(n_8512),
.B2(n_8352),
.Y(n_9077)
);

NAND2xp5_ASAP7_75t_L g9078 ( 
.A(n_8478),
.B(n_143),
.Y(n_9078)
);

INVx3_ASAP7_75t_L g9079 ( 
.A(n_8501),
.Y(n_9079)
);

BUFx5_ASAP7_75t_L g9080 ( 
.A(n_8648),
.Y(n_9080)
);

NAND2xp5_ASAP7_75t_SL g9081 ( 
.A(n_8566),
.B(n_143),
.Y(n_9081)
);

NAND2xp5_ASAP7_75t_L g9082 ( 
.A(n_8518),
.B(n_145),
.Y(n_9082)
);

AND2x2_ASAP7_75t_L g9083 ( 
.A(n_8652),
.B(n_145),
.Y(n_9083)
);

NOR2xp33_ASAP7_75t_L g9084 ( 
.A(n_8425),
.B(n_3487),
.Y(n_9084)
);

NAND2xp5_ASAP7_75t_L g9085 ( 
.A(n_8379),
.B(n_146),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_8550),
.Y(n_9086)
);

NAND2xp5_ASAP7_75t_L g9087 ( 
.A(n_8380),
.B(n_146),
.Y(n_9087)
);

AOI22xp5_ASAP7_75t_L g9088 ( 
.A1(n_8664),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_9088)
);

BUFx6f_ASAP7_75t_L g9089 ( 
.A(n_8579),
.Y(n_9089)
);

INVxp67_ASAP7_75t_L g9090 ( 
.A(n_8660),
.Y(n_9090)
);

INVx5_ASAP7_75t_L g9091 ( 
.A(n_8661),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_L g9092 ( 
.A(n_8383),
.B(n_148),
.Y(n_9092)
);

AOI22xp33_ASAP7_75t_L g9093 ( 
.A1(n_8647),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_9093)
);

AOI21xp5_ASAP7_75t_L g9094 ( 
.A1(n_8609),
.A2(n_3489),
.B(n_3488),
.Y(n_9094)
);

NAND2xp5_ASAP7_75t_L g9095 ( 
.A(n_8391),
.B(n_8465),
.Y(n_9095)
);

INVx1_ASAP7_75t_L g9096 ( 
.A(n_8558),
.Y(n_9096)
);

INVx2_ASAP7_75t_L g9097 ( 
.A(n_8559),
.Y(n_9097)
);

INVx2_ASAP7_75t_L g9098 ( 
.A(n_8567),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_8571),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8574),
.Y(n_9100)
);

AOI22xp33_ASAP7_75t_L g9101 ( 
.A1(n_8385),
.A2(n_153),
.B1(n_150),
.B2(n_152),
.Y(n_9101)
);

INVx2_ASAP7_75t_L g9102 ( 
.A(n_8585),
.Y(n_9102)
);

INVxp33_ASAP7_75t_L g9103 ( 
.A(n_8653),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_8591),
.Y(n_9104)
);

NAND2x1p5_ASAP7_75t_L g9105 ( 
.A(n_8521),
.B(n_3490),
.Y(n_9105)
);

BUFx3_ASAP7_75t_L g9106 ( 
.A(n_8608),
.Y(n_9106)
);

HB1xp67_ASAP7_75t_L g9107 ( 
.A(n_8612),
.Y(n_9107)
);

NAND2xp5_ASAP7_75t_L g9108 ( 
.A(n_8468),
.B(n_152),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_8398),
.Y(n_9109)
);

INVx1_ASAP7_75t_L g9110 ( 
.A(n_8402),
.Y(n_9110)
);

CKINVDCx5p33_ASAP7_75t_R g9111 ( 
.A(n_8434),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8405),
.Y(n_9112)
);

AND2x2_ASAP7_75t_L g9113 ( 
.A(n_8460),
.B(n_153),
.Y(n_9113)
);

AOI22xp33_ASAP7_75t_L g9114 ( 
.A1(n_8350),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_9114)
);

NAND2xp5_ASAP7_75t_L g9115 ( 
.A(n_8410),
.B(n_155),
.Y(n_9115)
);

AND2x4_ASAP7_75t_L g9116 ( 
.A(n_8544),
.B(n_3491),
.Y(n_9116)
);

A2O1A1Ixp33_ASAP7_75t_L g9117 ( 
.A1(n_8252),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8417),
.Y(n_9118)
);

OR2x6_ASAP7_75t_L g9119 ( 
.A(n_8394),
.B(n_3492),
.Y(n_9119)
);

INVx2_ASAP7_75t_L g9120 ( 
.A(n_8469),
.Y(n_9120)
);

BUFx2_ASAP7_75t_L g9121 ( 
.A(n_8469),
.Y(n_9121)
);

INVx2_ASAP7_75t_L g9122 ( 
.A(n_8469),
.Y(n_9122)
);

NAND2xp5_ASAP7_75t_L g9123 ( 
.A(n_8420),
.B(n_157),
.Y(n_9123)
);

A2O1A1Ixp33_ASAP7_75t_L g9124 ( 
.A1(n_8441),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_9124)
);

INVx5_ASAP7_75t_L g9125 ( 
.A(n_8662),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_8421),
.Y(n_9126)
);

AND2x4_ASAP7_75t_L g9127 ( 
.A(n_8621),
.B(n_3493),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_8427),
.B(n_160),
.Y(n_9128)
);

AND2x4_ASAP7_75t_L g9129 ( 
.A(n_8636),
.B(n_3494),
.Y(n_9129)
);

BUFx3_ASAP7_75t_L g9130 ( 
.A(n_8469),
.Y(n_9130)
);

NOR3xp33_ASAP7_75t_SL g9131 ( 
.A(n_8668),
.B(n_161),
.C(n_162),
.Y(n_9131)
);

INVx3_ASAP7_75t_L g9132 ( 
.A(n_8522),
.Y(n_9132)
);

NAND2xp5_ASAP7_75t_SL g9133 ( 
.A(n_8666),
.B(n_161),
.Y(n_9133)
);

INVx2_ASAP7_75t_L g9134 ( 
.A(n_8522),
.Y(n_9134)
);

INVx1_ASAP7_75t_L g9135 ( 
.A(n_8428),
.Y(n_9135)
);

NAND2xp5_ASAP7_75t_L g9136 ( 
.A(n_8449),
.B(n_163),
.Y(n_9136)
);

AND2x2_ASAP7_75t_L g9137 ( 
.A(n_8477),
.B(n_163),
.Y(n_9137)
);

INVxp67_ASAP7_75t_L g9138 ( 
.A(n_8492),
.Y(n_9138)
);

CKINVDCx5p33_ASAP7_75t_R g9139 ( 
.A(n_8562),
.Y(n_9139)
);

INVx2_ASAP7_75t_L g9140 ( 
.A(n_8522),
.Y(n_9140)
);

NAND2xp5_ASAP7_75t_L g9141 ( 
.A(n_8452),
.B(n_164),
.Y(n_9141)
);

INVx1_ASAP7_75t_L g9142 ( 
.A(n_8454),
.Y(n_9142)
);

NAND2xp5_ASAP7_75t_SL g9143 ( 
.A(n_8590),
.B(n_164),
.Y(n_9143)
);

INVx1_ASAP7_75t_L g9144 ( 
.A(n_8456),
.Y(n_9144)
);

INVx1_ASAP7_75t_L g9145 ( 
.A(n_8640),
.Y(n_9145)
);

NOR2xp33_ASAP7_75t_R g9146 ( 
.A(n_8522),
.B(n_3495),
.Y(n_9146)
);

AND2x2_ASAP7_75t_SL g9147 ( 
.A(n_8642),
.B(n_165),
.Y(n_9147)
);

INVx1_ASAP7_75t_L g9148 ( 
.A(n_8322),
.Y(n_9148)
);

INVx3_ASAP7_75t_L g9149 ( 
.A(n_8498),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_8615),
.Y(n_9150)
);

NAND2xp5_ASAP7_75t_L g9151 ( 
.A(n_8504),
.B(n_166),
.Y(n_9151)
);

INVx4_ASAP7_75t_L g9152 ( 
.A(n_8617),
.Y(n_9152)
);

INVx1_ASAP7_75t_L g9153 ( 
.A(n_8534),
.Y(n_9153)
);

INVx2_ASAP7_75t_L g9154 ( 
.A(n_8499),
.Y(n_9154)
);

INVxp67_ASAP7_75t_SL g9155 ( 
.A(n_8502),
.Y(n_9155)
);

OAI22xp5_ASAP7_75t_SL g9156 ( 
.A1(n_8496),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.Y(n_9156)
);

BUFx6f_ASAP7_75t_L g9157 ( 
.A(n_8422),
.Y(n_9157)
);

BUFx6f_ASAP7_75t_L g9158 ( 
.A(n_8397),
.Y(n_9158)
);

NOR3xp33_ASAP7_75t_SL g9159 ( 
.A(n_8703),
.B(n_8539),
.C(n_8326),
.Y(n_9159)
);

NOR2xp33_ASAP7_75t_L g9160 ( 
.A(n_8411),
.B(n_3496),
.Y(n_9160)
);

INVx1_ASAP7_75t_L g9161 ( 
.A(n_8543),
.Y(n_9161)
);

NOR2x2_ASAP7_75t_L g9162 ( 
.A(n_8409),
.B(n_168),
.Y(n_9162)
);

INVx1_ASAP7_75t_L g9163 ( 
.A(n_8545),
.Y(n_9163)
);

AOI21xp5_ASAP7_75t_L g9164 ( 
.A1(n_8490),
.A2(n_3498),
.B(n_3497),
.Y(n_9164)
);

AOI22xp33_ASAP7_75t_L g9165 ( 
.A1(n_8602),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_9165)
);

NAND2xp5_ASAP7_75t_L g9166 ( 
.A(n_8511),
.B(n_170),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_L g9167 ( 
.A(n_8515),
.B(n_8547),
.Y(n_9167)
);

BUFx2_ASAP7_75t_L g9168 ( 
.A(n_8553),
.Y(n_9168)
);

NAND2xp33_ASAP7_75t_SL g9169 ( 
.A(n_8412),
.B(n_173),
.Y(n_9169)
);

OAI22xp5_ASAP7_75t_L g9170 ( 
.A1(n_8627),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_9170)
);

INVx2_ASAP7_75t_L g9171 ( 
.A(n_8554),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_8563),
.Y(n_9172)
);

NOR2xp33_ASAP7_75t_L g9173 ( 
.A(n_8600),
.B(n_3499),
.Y(n_9173)
);

AND2x2_ASAP7_75t_SL g9174 ( 
.A(n_8632),
.B(n_175),
.Y(n_9174)
);

AND2x4_ASAP7_75t_L g9175 ( 
.A(n_8628),
.B(n_3500),
.Y(n_9175)
);

NAND2xp5_ASAP7_75t_L g9176 ( 
.A(n_8573),
.B(n_177),
.Y(n_9176)
);

INVx1_ASAP7_75t_SL g9177 ( 
.A(n_8575),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_8578),
.Y(n_9178)
);

INVx1_ASAP7_75t_L g9179 ( 
.A(n_8580),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_8592),
.Y(n_9180)
);

INVxp67_ASAP7_75t_L g9181 ( 
.A(n_8635),
.Y(n_9181)
);

INVx1_ASAP7_75t_SL g9182 ( 
.A(n_8595),
.Y(n_9182)
);

AOI22xp5_ASAP7_75t_L g9183 ( 
.A1(n_8342),
.A2(n_180),
.B1(n_177),
.B2(n_179),
.Y(n_9183)
);

AOI21xp5_ASAP7_75t_L g9184 ( 
.A1(n_8702),
.A2(n_3503),
.B(n_3502),
.Y(n_9184)
);

BUFx8_ASAP7_75t_SL g9185 ( 
.A(n_8603),
.Y(n_9185)
);

BUFx8_ASAP7_75t_L g9186 ( 
.A(n_8377),
.Y(n_9186)
);

INVx1_ASAP7_75t_L g9187 ( 
.A(n_8607),
.Y(n_9187)
);

NAND2xp5_ASAP7_75t_SL g9188 ( 
.A(n_8610),
.B(n_179),
.Y(n_9188)
);

BUFx6f_ASAP7_75t_L g9189 ( 
.A(n_8616),
.Y(n_9189)
);

NAND2xp5_ASAP7_75t_L g9190 ( 
.A(n_8618),
.B(n_180),
.Y(n_9190)
);

INVx3_ASAP7_75t_L g9191 ( 
.A(n_8655),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_8436),
.Y(n_9192)
);

BUFx4f_ASAP7_75t_L g9193 ( 
.A(n_8484),
.Y(n_9193)
);

INVx2_ASAP7_75t_SL g9194 ( 
.A(n_8540),
.Y(n_9194)
);

HB1xp67_ASAP7_75t_L g9195 ( 
.A(n_8643),
.Y(n_9195)
);

INVx2_ASAP7_75t_L g9196 ( 
.A(n_8572),
.Y(n_9196)
);

CKINVDCx5p33_ASAP7_75t_R g9197 ( 
.A(n_8372),
.Y(n_9197)
);

BUFx6f_ASAP7_75t_L g9198 ( 
.A(n_8506),
.Y(n_9198)
);

NAND2x1p5_ASAP7_75t_L g9199 ( 
.A(n_8400),
.B(n_3505),
.Y(n_9199)
);

NOR2xp33_ASAP7_75t_L g9200 ( 
.A(n_8619),
.B(n_3508),
.Y(n_9200)
);

INVx2_ASAP7_75t_SL g9201 ( 
.A(n_8390),
.Y(n_9201)
);

INVx2_ASAP7_75t_L g9202 ( 
.A(n_8201),
.Y(n_9202)
);

INVx2_ASAP7_75t_SL g9203 ( 
.A(n_8390),
.Y(n_9203)
);

O2A1O1Ixp5_ASAP7_75t_L g9204 ( 
.A1(n_8259),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_9204)
);

INVx1_ASAP7_75t_L g9205 ( 
.A(n_8378),
.Y(n_9205)
);

NOR3x1_ASAP7_75t_L g9206 ( 
.A(n_8206),
.B(n_184),
.C(n_185),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_8378),
.Y(n_9207)
);

NAND2x1p5_ASAP7_75t_L g9208 ( 
.A(n_8347),
.B(n_3509),
.Y(n_9208)
);

AND2x4_ASAP7_75t_L g9209 ( 
.A(n_8223),
.B(n_3510),
.Y(n_9209)
);

NOR2xp33_ASAP7_75t_L g9210 ( 
.A(n_8442),
.B(n_3511),
.Y(n_9210)
);

BUFx2_ASAP7_75t_L g9211 ( 
.A(n_8315),
.Y(n_9211)
);

INVx1_ASAP7_75t_L g9212 ( 
.A(n_8378),
.Y(n_9212)
);

NOR2xp33_ASAP7_75t_R g9213 ( 
.A(n_8459),
.B(n_3514),
.Y(n_9213)
);

INVx1_ASAP7_75t_L g9214 ( 
.A(n_8378),
.Y(n_9214)
);

INVx2_ASAP7_75t_L g9215 ( 
.A(n_8201),
.Y(n_9215)
);

AND2x4_ASAP7_75t_L g9216 ( 
.A(n_8223),
.B(n_3516),
.Y(n_9216)
);

INVx2_ASAP7_75t_L g9217 ( 
.A(n_8201),
.Y(n_9217)
);

BUFx6f_ASAP7_75t_L g9218 ( 
.A(n_8205),
.Y(n_9218)
);

NAND2xp5_ASAP7_75t_SL g9219 ( 
.A(n_8300),
.B(n_186),
.Y(n_9219)
);

AND2x6_ASAP7_75t_L g9220 ( 
.A(n_8204),
.B(n_3517),
.Y(n_9220)
);

NAND2xp5_ASAP7_75t_SL g9221 ( 
.A(n_8300),
.B(n_186),
.Y(n_9221)
);

INVx4_ASAP7_75t_L g9222 ( 
.A(n_8347),
.Y(n_9222)
);

AND2x4_ASAP7_75t_L g9223 ( 
.A(n_8223),
.B(n_3518),
.Y(n_9223)
);

NAND2xp5_ASAP7_75t_SL g9224 ( 
.A(n_8300),
.B(n_187),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_SL g9225 ( 
.A(n_8300),
.B(n_187),
.Y(n_9225)
);

AND2x4_ASAP7_75t_L g9226 ( 
.A(n_8223),
.B(n_3519),
.Y(n_9226)
);

BUFx6f_ASAP7_75t_L g9227 ( 
.A(n_8205),
.Y(n_9227)
);

BUFx3_ASAP7_75t_L g9228 ( 
.A(n_8223),
.Y(n_9228)
);

BUFx12f_ASAP7_75t_L g9229 ( 
.A(n_8381),
.Y(n_9229)
);

NOR2xp33_ASAP7_75t_L g9230 ( 
.A(n_8442),
.B(n_3521),
.Y(n_9230)
);

NAND2xp5_ASAP7_75t_L g9231 ( 
.A(n_8237),
.B(n_188),
.Y(n_9231)
);

NAND2xp5_ASAP7_75t_L g9232 ( 
.A(n_8237),
.B(n_189),
.Y(n_9232)
);

AND2x2_ASAP7_75t_L g9233 ( 
.A(n_8336),
.B(n_189),
.Y(n_9233)
);

NAND2xp5_ASAP7_75t_L g9234 ( 
.A(n_8237),
.B(n_190),
.Y(n_9234)
);

NAND2xp5_ASAP7_75t_SL g9235 ( 
.A(n_8300),
.B(n_191),
.Y(n_9235)
);

INVx2_ASAP7_75t_SL g9236 ( 
.A(n_8390),
.Y(n_9236)
);

NAND2xp5_ASAP7_75t_L g9237 ( 
.A(n_8237),
.B(n_191),
.Y(n_9237)
);

INVx2_ASAP7_75t_L g9238 ( 
.A(n_8201),
.Y(n_9238)
);

OR2x2_ASAP7_75t_L g9239 ( 
.A(n_8264),
.B(n_192),
.Y(n_9239)
);

INVx1_ASAP7_75t_L g9240 ( 
.A(n_8378),
.Y(n_9240)
);

NAND2xp5_ASAP7_75t_SL g9241 ( 
.A(n_8300),
.B(n_193),
.Y(n_9241)
);

CKINVDCx5p33_ASAP7_75t_R g9242 ( 
.A(n_8459),
.Y(n_9242)
);

INVx2_ASAP7_75t_L g9243 ( 
.A(n_8201),
.Y(n_9243)
);

INVx2_ASAP7_75t_L g9244 ( 
.A(n_8201),
.Y(n_9244)
);

INVx5_ASAP7_75t_L g9245 ( 
.A(n_8347),
.Y(n_9245)
);

AND2x2_ASAP7_75t_L g9246 ( 
.A(n_8336),
.B(n_193),
.Y(n_9246)
);

AND2x2_ASAP7_75t_L g9247 ( 
.A(n_8336),
.B(n_194),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_8378),
.Y(n_9248)
);

INVx2_ASAP7_75t_L g9249 ( 
.A(n_8201),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_8378),
.Y(n_9250)
);

NOR2xp67_ASAP7_75t_L g9251 ( 
.A(n_8314),
.B(n_3522),
.Y(n_9251)
);

AOI22xp33_ASAP7_75t_L g9252 ( 
.A1(n_8300),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.Y(n_9252)
);

INVx2_ASAP7_75t_L g9253 ( 
.A(n_8201),
.Y(n_9253)
);

NOR2xp33_ASAP7_75t_R g9254 ( 
.A(n_8459),
.B(n_3524),
.Y(n_9254)
);

INVx1_ASAP7_75t_L g9255 ( 
.A(n_8378),
.Y(n_9255)
);

INVx1_ASAP7_75t_L g9256 ( 
.A(n_8378),
.Y(n_9256)
);

AOI22xp33_ASAP7_75t_L g9257 ( 
.A1(n_8300),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_9257)
);

NAND2xp5_ASAP7_75t_L g9258 ( 
.A(n_8237),
.B(n_199),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_8378),
.Y(n_9259)
);

NOR2xp33_ASAP7_75t_L g9260 ( 
.A(n_8442),
.B(n_3528),
.Y(n_9260)
);

INVx1_ASAP7_75t_L g9261 ( 
.A(n_8378),
.Y(n_9261)
);

INVx1_ASAP7_75t_L g9262 ( 
.A(n_8378),
.Y(n_9262)
);

INVx2_ASAP7_75t_L g9263 ( 
.A(n_8201),
.Y(n_9263)
);

INVx2_ASAP7_75t_L g9264 ( 
.A(n_8201),
.Y(n_9264)
);

AOI22xp33_ASAP7_75t_L g9265 ( 
.A1(n_8300),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_9265)
);

INVx2_ASAP7_75t_L g9266 ( 
.A(n_8201),
.Y(n_9266)
);

NAND2xp5_ASAP7_75t_L g9267 ( 
.A(n_8237),
.B(n_202),
.Y(n_9267)
);

INVx1_ASAP7_75t_L g9268 ( 
.A(n_8378),
.Y(n_9268)
);

NAND2xp5_ASAP7_75t_L g9269 ( 
.A(n_8237),
.B(n_202),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_8237),
.B(n_203),
.Y(n_9270)
);

NAND2xp5_ASAP7_75t_SL g9271 ( 
.A(n_8300),
.B(n_204),
.Y(n_9271)
);

AOI22x1_ASAP7_75t_L g9272 ( 
.A1(n_8448),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_9272)
);

NOR2x1_ASAP7_75t_L g9273 ( 
.A(n_8437),
.B(n_3529),
.Y(n_9273)
);

AOI22xp33_ASAP7_75t_L g9274 ( 
.A1(n_8300),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_9274)
);

NAND2xp5_ASAP7_75t_SL g9275 ( 
.A(n_8300),
.B(n_208),
.Y(n_9275)
);

AOI22xp5_ASAP7_75t_L g9276 ( 
.A1(n_8300),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_9276)
);

XNOR2xp5_ASAP7_75t_L g9277 ( 
.A(n_8459),
.B(n_3530),
.Y(n_9277)
);

AND2x4_ASAP7_75t_L g9278 ( 
.A(n_8223),
.B(n_3531),
.Y(n_9278)
);

INVx1_ASAP7_75t_L g9279 ( 
.A(n_8378),
.Y(n_9279)
);

INVx2_ASAP7_75t_L g9280 ( 
.A(n_8201),
.Y(n_9280)
);

BUFx3_ASAP7_75t_L g9281 ( 
.A(n_8223),
.Y(n_9281)
);

AND2x6_ASAP7_75t_SL g9282 ( 
.A(n_8644),
.B(n_210),
.Y(n_9282)
);

HB1xp67_ASAP7_75t_L g9283 ( 
.A(n_8216),
.Y(n_9283)
);

INVx2_ASAP7_75t_L g9284 ( 
.A(n_8201),
.Y(n_9284)
);

INVx2_ASAP7_75t_L g9285 ( 
.A(n_8201),
.Y(n_9285)
);

AND2x6_ASAP7_75t_L g9286 ( 
.A(n_8204),
.B(n_3532),
.Y(n_9286)
);

INVx2_ASAP7_75t_L g9287 ( 
.A(n_8201),
.Y(n_9287)
);

NOR2xp33_ASAP7_75t_L g9288 ( 
.A(n_8442),
.B(n_3535),
.Y(n_9288)
);

INVx1_ASAP7_75t_L g9289 ( 
.A(n_8378),
.Y(n_9289)
);

AND2x2_ASAP7_75t_L g9290 ( 
.A(n_8336),
.B(n_211),
.Y(n_9290)
);

AOI22xp5_ASAP7_75t_L g9291 ( 
.A1(n_8300),
.A2(n_215),
.B1(n_212),
.B2(n_213),
.Y(n_9291)
);

INVx2_ASAP7_75t_SL g9292 ( 
.A(n_8390),
.Y(n_9292)
);

INVx3_ASAP7_75t_L g9293 ( 
.A(n_8347),
.Y(n_9293)
);

NOR2xp33_ASAP7_75t_R g9294 ( 
.A(n_8459),
.B(n_3536),
.Y(n_9294)
);

BUFx3_ASAP7_75t_L g9295 ( 
.A(n_8223),
.Y(n_9295)
);

INVx1_ASAP7_75t_SL g9296 ( 
.A(n_8216),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8378),
.Y(n_9297)
);

INVx2_ASAP7_75t_L g9298 ( 
.A(n_8201),
.Y(n_9298)
);

INVx1_ASAP7_75t_L g9299 ( 
.A(n_8378),
.Y(n_9299)
);

INVx2_ASAP7_75t_SL g9300 ( 
.A(n_8390),
.Y(n_9300)
);

INVx1_ASAP7_75t_L g9301 ( 
.A(n_9059),
.Y(n_9301)
);

HB1xp67_ASAP7_75t_L g9302 ( 
.A(n_8856),
.Y(n_9302)
);

CKINVDCx5p33_ASAP7_75t_R g9303 ( 
.A(n_8853),
.Y(n_9303)
);

NAND2xp5_ASAP7_75t_L g9304 ( 
.A(n_8713),
.B(n_213),
.Y(n_9304)
);

HB1xp67_ASAP7_75t_L g9305 ( 
.A(n_8890),
.Y(n_9305)
);

NOR2xp33_ASAP7_75t_R g9306 ( 
.A(n_8715),
.B(n_3539),
.Y(n_9306)
);

BUFx6f_ASAP7_75t_L g9307 ( 
.A(n_8722),
.Y(n_9307)
);

BUFx12f_ASAP7_75t_L g9308 ( 
.A(n_8840),
.Y(n_9308)
);

BUFx4f_ASAP7_75t_L g9309 ( 
.A(n_9229),
.Y(n_9309)
);

INVx1_ASAP7_75t_SL g9310 ( 
.A(n_8907),
.Y(n_9310)
);

INVx5_ASAP7_75t_L g9311 ( 
.A(n_8722),
.Y(n_9311)
);

A2O1A1Ixp33_ASAP7_75t_L g9312 ( 
.A1(n_8719),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_9312)
);

NAND2xp5_ASAP7_75t_L g9313 ( 
.A(n_8767),
.B(n_216),
.Y(n_9313)
);

BUFx2_ASAP7_75t_L g9314 ( 
.A(n_8754),
.Y(n_9314)
);

AOI22xp33_ASAP7_75t_L g9315 ( 
.A1(n_9193),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_9315)
);

BUFx6f_ASAP7_75t_L g9316 ( 
.A(n_9218),
.Y(n_9316)
);

AND2x4_ASAP7_75t_L g9317 ( 
.A(n_8864),
.B(n_3542),
.Y(n_9317)
);

NAND2xp5_ASAP7_75t_L g9318 ( 
.A(n_9043),
.B(n_218),
.Y(n_9318)
);

INVxp67_ASAP7_75t_L g9319 ( 
.A(n_8732),
.Y(n_9319)
);

INVx1_ASAP7_75t_L g9320 ( 
.A(n_9107),
.Y(n_9320)
);

NAND2xp5_ASAP7_75t_L g9321 ( 
.A(n_8832),
.B(n_219),
.Y(n_9321)
);

HB1xp67_ASAP7_75t_L g9322 ( 
.A(n_8953),
.Y(n_9322)
);

INVx1_ASAP7_75t_L g9323 ( 
.A(n_8855),
.Y(n_9323)
);

CKINVDCx5p33_ASAP7_75t_R g9324 ( 
.A(n_8797),
.Y(n_9324)
);

HB1xp67_ASAP7_75t_L g9325 ( 
.A(n_8972),
.Y(n_9325)
);

NAND2xp5_ASAP7_75t_L g9326 ( 
.A(n_8812),
.B(n_220),
.Y(n_9326)
);

NAND2xp5_ASAP7_75t_L g9327 ( 
.A(n_9155),
.B(n_221),
.Y(n_9327)
);

INVx3_ASAP7_75t_SL g9328 ( 
.A(n_9242),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_8859),
.Y(n_9329)
);

AND2x4_ASAP7_75t_L g9330 ( 
.A(n_8783),
.B(n_3543),
.Y(n_9330)
);

AND2x2_ASAP7_75t_L g9331 ( 
.A(n_8778),
.B(n_3544),
.Y(n_9331)
);

NAND2xp5_ASAP7_75t_L g9332 ( 
.A(n_8741),
.B(n_222),
.Y(n_9332)
);

INVx4_ASAP7_75t_L g9333 ( 
.A(n_9245),
.Y(n_9333)
);

BUFx2_ASAP7_75t_L g9334 ( 
.A(n_9283),
.Y(n_9334)
);

AND2x2_ASAP7_75t_L g9335 ( 
.A(n_8752),
.B(n_3545),
.Y(n_9335)
);

INVx6_ASAP7_75t_L g9336 ( 
.A(n_8860),
.Y(n_9336)
);

NOR2xp33_ASAP7_75t_L g9337 ( 
.A(n_8837),
.B(n_3546),
.Y(n_9337)
);

AND2x2_ASAP7_75t_L g9338 ( 
.A(n_9290),
.B(n_3547),
.Y(n_9338)
);

INVxp67_ASAP7_75t_L g9339 ( 
.A(n_8799),
.Y(n_9339)
);

INVx1_ASAP7_75t_SL g9340 ( 
.A(n_9296),
.Y(n_9340)
);

AND2x4_ASAP7_75t_L g9341 ( 
.A(n_8968),
.B(n_3548),
.Y(n_9341)
);

BUFx2_ASAP7_75t_L g9342 ( 
.A(n_9074),
.Y(n_9342)
);

INVx1_ASAP7_75t_L g9343 ( 
.A(n_8861),
.Y(n_9343)
);

INVx2_ASAP7_75t_L g9344 ( 
.A(n_8709),
.Y(n_9344)
);

INVx3_ASAP7_75t_L g9345 ( 
.A(n_8736),
.Y(n_9345)
);

INVx1_ASAP7_75t_L g9346 ( 
.A(n_8863),
.Y(n_9346)
);

INVx2_ASAP7_75t_L g9347 ( 
.A(n_8711),
.Y(n_9347)
);

AND2x2_ASAP7_75t_L g9348 ( 
.A(n_9233),
.B(n_3555),
.Y(n_9348)
);

NOR2xp33_ASAP7_75t_L g9349 ( 
.A(n_8959),
.B(n_3559),
.Y(n_9349)
);

NAND2xp5_ASAP7_75t_L g9350 ( 
.A(n_8710),
.B(n_223),
.Y(n_9350)
);

INVx4_ASAP7_75t_L g9351 ( 
.A(n_9245),
.Y(n_9351)
);

INVx3_ASAP7_75t_L g9352 ( 
.A(n_8774),
.Y(n_9352)
);

INVx3_ASAP7_75t_L g9353 ( 
.A(n_9228),
.Y(n_9353)
);

NAND2xp5_ASAP7_75t_L g9354 ( 
.A(n_8718),
.B(n_223),
.Y(n_9354)
);

INVx1_ASAP7_75t_L g9355 ( 
.A(n_8869),
.Y(n_9355)
);

BUFx2_ASAP7_75t_L g9356 ( 
.A(n_9028),
.Y(n_9356)
);

BUFx12f_ASAP7_75t_L g9357 ( 
.A(n_8943),
.Y(n_9357)
);

INVx1_ASAP7_75t_L g9358 ( 
.A(n_8870),
.Y(n_9358)
);

NAND2xp5_ASAP7_75t_L g9359 ( 
.A(n_8728),
.B(n_224),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_9205),
.B(n_224),
.Y(n_9360)
);

NOR3xp33_ASAP7_75t_SL g9361 ( 
.A(n_9197),
.B(n_225),
.C(n_226),
.Y(n_9361)
);

BUFx2_ASAP7_75t_L g9362 ( 
.A(n_8968),
.Y(n_9362)
);

HB1xp67_ASAP7_75t_L g9363 ( 
.A(n_9010),
.Y(n_9363)
);

INVx2_ASAP7_75t_SL g9364 ( 
.A(n_9218),
.Y(n_9364)
);

AOI22xp5_ASAP7_75t_L g9365 ( 
.A1(n_9077),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_8881),
.Y(n_9366)
);

INVx2_ASAP7_75t_L g9367 ( 
.A(n_8714),
.Y(n_9367)
);

NOR3xp33_ASAP7_75t_SL g9368 ( 
.A(n_9219),
.B(n_9224),
.C(n_9221),
.Y(n_9368)
);

INVx2_ASAP7_75t_L g9369 ( 
.A(n_8724),
.Y(n_9369)
);

NAND2xp5_ASAP7_75t_L g9370 ( 
.A(n_9207),
.B(n_227),
.Y(n_9370)
);

NOR2xp33_ASAP7_75t_R g9371 ( 
.A(n_8973),
.B(n_3560),
.Y(n_9371)
);

INVx2_ASAP7_75t_L g9372 ( 
.A(n_8727),
.Y(n_9372)
);

BUFx6f_ASAP7_75t_L g9373 ( 
.A(n_9227),
.Y(n_9373)
);

BUFx2_ASAP7_75t_L g9374 ( 
.A(n_8758),
.Y(n_9374)
);

NAND2xp5_ASAP7_75t_L g9375 ( 
.A(n_9212),
.B(n_228),
.Y(n_9375)
);

BUFx4f_ASAP7_75t_SL g9376 ( 
.A(n_9040),
.Y(n_9376)
);

INVx2_ASAP7_75t_L g9377 ( 
.A(n_8740),
.Y(n_9377)
);

NAND2xp5_ASAP7_75t_L g9378 ( 
.A(n_9214),
.B(n_229),
.Y(n_9378)
);

CKINVDCx5p33_ASAP7_75t_R g9379 ( 
.A(n_8895),
.Y(n_9379)
);

NAND2xp5_ASAP7_75t_L g9380 ( 
.A(n_9240),
.B(n_230),
.Y(n_9380)
);

NAND2xp5_ASAP7_75t_L g9381 ( 
.A(n_9248),
.B(n_230),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8902),
.Y(n_9382)
);

AND3x1_ASAP7_75t_L g9383 ( 
.A(n_8929),
.B(n_231),
.C(n_232),
.Y(n_9383)
);

AND2x4_ASAP7_75t_L g9384 ( 
.A(n_8769),
.B(n_3562),
.Y(n_9384)
);

INVx1_ASAP7_75t_L g9385 ( 
.A(n_8904),
.Y(n_9385)
);

AND2x4_ASAP7_75t_L g9386 ( 
.A(n_8923),
.B(n_3563),
.Y(n_9386)
);

AND3x1_ASAP7_75t_SL g9387 ( 
.A(n_9065),
.B(n_231),
.C(n_233),
.Y(n_9387)
);

CKINVDCx5p33_ASAP7_75t_R g9388 ( 
.A(n_8901),
.Y(n_9388)
);

NAND2xp5_ASAP7_75t_L g9389 ( 
.A(n_9250),
.B(n_233),
.Y(n_9389)
);

NAND2xp5_ASAP7_75t_L g9390 ( 
.A(n_9255),
.B(n_234),
.Y(n_9390)
);

NOR3xp33_ASAP7_75t_SL g9391 ( 
.A(n_9225),
.B(n_9241),
.C(n_9235),
.Y(n_9391)
);

INVx2_ASAP7_75t_L g9392 ( 
.A(n_8749),
.Y(n_9392)
);

INVx2_ASAP7_75t_L g9393 ( 
.A(n_8753),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_8910),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_8918),
.Y(n_9395)
);

BUFx8_ASAP7_75t_L g9396 ( 
.A(n_9211),
.Y(n_9396)
);

INVx2_ASAP7_75t_L g9397 ( 
.A(n_8757),
.Y(n_9397)
);

INVx1_ASAP7_75t_L g9398 ( 
.A(n_8932),
.Y(n_9398)
);

NOR3xp33_ASAP7_75t_SL g9399 ( 
.A(n_9271),
.B(n_234),
.C(n_235),
.Y(n_9399)
);

INVx1_ASAP7_75t_L g9400 ( 
.A(n_8934),
.Y(n_9400)
);

NOR2xp33_ASAP7_75t_L g9401 ( 
.A(n_9090),
.B(n_3564),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_8772),
.Y(n_9402)
);

AND2x6_ASAP7_75t_L g9403 ( 
.A(n_9206),
.B(n_3565),
.Y(n_9403)
);

OR2x6_ASAP7_75t_L g9404 ( 
.A(n_8865),
.B(n_3566),
.Y(n_9404)
);

OR2x6_ASAP7_75t_L g9405 ( 
.A(n_8865),
.B(n_3567),
.Y(n_9405)
);

INVx1_ASAP7_75t_L g9406 ( 
.A(n_8938),
.Y(n_9406)
);

A2O1A1Ixp33_ASAP7_75t_L g9407 ( 
.A1(n_8725),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_9407)
);

BUFx6f_ASAP7_75t_L g9408 ( 
.A(n_9227),
.Y(n_9408)
);

INVx3_ASAP7_75t_L g9409 ( 
.A(n_9281),
.Y(n_9409)
);

NAND2xp5_ASAP7_75t_L g9410 ( 
.A(n_9256),
.B(n_236),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_8939),
.Y(n_9411)
);

AND2x4_ASAP7_75t_L g9412 ( 
.A(n_8887),
.B(n_3568),
.Y(n_9412)
);

AND2x2_ASAP7_75t_L g9413 ( 
.A(n_9246),
.B(n_3569),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_8940),
.Y(n_9414)
);

INVx2_ASAP7_75t_L g9415 ( 
.A(n_8779),
.Y(n_9415)
);

BUFx2_ASAP7_75t_L g9416 ( 
.A(n_8925),
.Y(n_9416)
);

BUFx6f_ASAP7_75t_L g9417 ( 
.A(n_8716),
.Y(n_9417)
);

NAND2xp5_ASAP7_75t_L g9418 ( 
.A(n_9259),
.B(n_237),
.Y(n_9418)
);

INVx5_ASAP7_75t_L g9419 ( 
.A(n_8735),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_8946),
.Y(n_9420)
);

INVx2_ASAP7_75t_L g9421 ( 
.A(n_8782),
.Y(n_9421)
);

BUFx6f_ASAP7_75t_L g9422 ( 
.A(n_8729),
.Y(n_9422)
);

NOR2xp33_ASAP7_75t_R g9423 ( 
.A(n_9072),
.B(n_3570),
.Y(n_9423)
);

INVx3_ASAP7_75t_L g9424 ( 
.A(n_9295),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_8962),
.Y(n_9425)
);

AND2x4_ASAP7_75t_L g9426 ( 
.A(n_8889),
.B(n_3572),
.Y(n_9426)
);

AND2x2_ASAP7_75t_L g9427 ( 
.A(n_9247),
.B(n_3574),
.Y(n_9427)
);

INVx2_ASAP7_75t_L g9428 ( 
.A(n_8802),
.Y(n_9428)
);

NAND2xp5_ASAP7_75t_L g9429 ( 
.A(n_9261),
.B(n_238),
.Y(n_9429)
);

INVx2_ASAP7_75t_L g9430 ( 
.A(n_8803),
.Y(n_9430)
);

AND2x4_ASAP7_75t_L g9431 ( 
.A(n_8978),
.B(n_3575),
.Y(n_9431)
);

AND2x4_ASAP7_75t_L g9432 ( 
.A(n_8721),
.B(n_3576),
.Y(n_9432)
);

AOI22xp33_ASAP7_75t_L g9433 ( 
.A1(n_8965),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_9433)
);

NOR3xp33_ASAP7_75t_SL g9434 ( 
.A(n_9275),
.B(n_239),
.C(n_240),
.Y(n_9434)
);

NAND2xp5_ASAP7_75t_L g9435 ( 
.A(n_9262),
.B(n_241),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_8970),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_8979),
.Y(n_9437)
);

O2A1O1Ixp33_ASAP7_75t_L g9438 ( 
.A1(n_8893),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_9438)
);

NOR2xp33_ASAP7_75t_L g9439 ( 
.A(n_9036),
.B(n_3577),
.Y(n_9439)
);

INVx1_ASAP7_75t_L g9440 ( 
.A(n_8980),
.Y(n_9440)
);

NAND2xp33_ASAP7_75t_SL g9441 ( 
.A(n_9146),
.B(n_244),
.Y(n_9441)
);

INVx1_ASAP7_75t_L g9442 ( 
.A(n_8985),
.Y(n_9442)
);

INVx2_ASAP7_75t_L g9443 ( 
.A(n_8809),
.Y(n_9443)
);

BUFx4f_ASAP7_75t_L g9444 ( 
.A(n_8735),
.Y(n_9444)
);

NAND2xp33_ASAP7_75t_SL g9445 ( 
.A(n_8849),
.B(n_245),
.Y(n_9445)
);

NOR2xp33_ASAP7_75t_R g9446 ( 
.A(n_9071),
.B(n_3578),
.Y(n_9446)
);

INVx2_ASAP7_75t_L g9447 ( 
.A(n_8831),
.Y(n_9447)
);

HB1xp67_ASAP7_75t_L g9448 ( 
.A(n_9106),
.Y(n_9448)
);

BUFx6f_ASAP7_75t_L g9449 ( 
.A(n_8733),
.Y(n_9449)
);

INVx1_ASAP7_75t_SL g9450 ( 
.A(n_8964),
.Y(n_9450)
);

INVxp67_ASAP7_75t_L g9451 ( 
.A(n_8826),
.Y(n_9451)
);

BUFx6f_ASAP7_75t_L g9452 ( 
.A(n_8787),
.Y(n_9452)
);

INVx2_ASAP7_75t_L g9453 ( 
.A(n_8838),
.Y(n_9453)
);

AOI22xp5_ASAP7_75t_L g9454 ( 
.A1(n_8961),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_9454)
);

INVx1_ASAP7_75t_L g9455 ( 
.A(n_8987),
.Y(n_9455)
);

BUFx2_ASAP7_75t_L g9456 ( 
.A(n_9054),
.Y(n_9456)
);

OR2x4_ASAP7_75t_L g9457 ( 
.A(n_9210),
.B(n_246),
.Y(n_9457)
);

AND2x4_ASAP7_75t_L g9458 ( 
.A(n_8750),
.B(n_3579),
.Y(n_9458)
);

BUFx2_ASAP7_75t_L g9459 ( 
.A(n_9061),
.Y(n_9459)
);

INVx4_ASAP7_75t_L g9460 ( 
.A(n_8787),
.Y(n_9460)
);

BUFx2_ASAP7_75t_L g9461 ( 
.A(n_8792),
.Y(n_9461)
);

AND2x4_ASAP7_75t_L g9462 ( 
.A(n_9201),
.B(n_3584),
.Y(n_9462)
);

NOR2xp33_ASAP7_75t_L g9463 ( 
.A(n_9103),
.B(n_3585),
.Y(n_9463)
);

BUFx2_ASAP7_75t_L g9464 ( 
.A(n_8720),
.Y(n_9464)
);

INVx1_ASAP7_75t_L g9465 ( 
.A(n_8998),
.Y(n_9465)
);

BUFx3_ASAP7_75t_L g9466 ( 
.A(n_8755),
.Y(n_9466)
);

OR2x2_ASAP7_75t_L g9467 ( 
.A(n_8730),
.B(n_247),
.Y(n_9467)
);

BUFx4f_ASAP7_75t_L g9468 ( 
.A(n_8874),
.Y(n_9468)
);

NOR2xp33_ASAP7_75t_L g9469 ( 
.A(n_8747),
.B(n_3586),
.Y(n_9469)
);

AND2x2_ASAP7_75t_L g9470 ( 
.A(n_8776),
.B(n_3587),
.Y(n_9470)
);

AOI22xp5_ASAP7_75t_L g9471 ( 
.A1(n_9084),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_9471)
);

BUFx2_ASAP7_75t_L g9472 ( 
.A(n_9030),
.Y(n_9472)
);

BUFx6f_ASAP7_75t_L g9473 ( 
.A(n_8874),
.Y(n_9473)
);

HB1xp67_ASAP7_75t_L g9474 ( 
.A(n_9075),
.Y(n_9474)
);

NAND2xp5_ASAP7_75t_L g9475 ( 
.A(n_9268),
.B(n_9279),
.Y(n_9475)
);

INVx2_ASAP7_75t_SL g9476 ( 
.A(n_8915),
.Y(n_9476)
);

NAND2xp5_ASAP7_75t_L g9477 ( 
.A(n_9289),
.B(n_248),
.Y(n_9477)
);

BUFx6f_ASAP7_75t_L g9478 ( 
.A(n_8877),
.Y(n_9478)
);

INVx2_ASAP7_75t_L g9479 ( 
.A(n_8839),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_9011),
.Y(n_9480)
);

INVx2_ASAP7_75t_L g9481 ( 
.A(n_8848),
.Y(n_9481)
);

INVx1_ASAP7_75t_L g9482 ( 
.A(n_9016),
.Y(n_9482)
);

NAND2xp5_ASAP7_75t_SL g9483 ( 
.A(n_8858),
.B(n_3588),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_9021),
.Y(n_9484)
);

INVx1_ASAP7_75t_L g9485 ( 
.A(n_9022),
.Y(n_9485)
);

INVx2_ASAP7_75t_L g9486 ( 
.A(n_8851),
.Y(n_9486)
);

AND2x4_ASAP7_75t_L g9487 ( 
.A(n_9203),
.B(n_3589),
.Y(n_9487)
);

INVx1_ASAP7_75t_L g9488 ( 
.A(n_9026),
.Y(n_9488)
);

NOR2xp33_ASAP7_75t_L g9489 ( 
.A(n_9139),
.B(n_3591),
.Y(n_9489)
);

INVx1_ASAP7_75t_L g9490 ( 
.A(n_9032),
.Y(n_9490)
);

NAND2xp5_ASAP7_75t_SL g9491 ( 
.A(n_9189),
.B(n_3593),
.Y(n_9491)
);

INVx1_ASAP7_75t_L g9492 ( 
.A(n_9039),
.Y(n_9492)
);

BUFx5_ASAP7_75t_L g9493 ( 
.A(n_8872),
.Y(n_9493)
);

BUFx2_ASAP7_75t_L g9494 ( 
.A(n_9030),
.Y(n_9494)
);

NAND2xp5_ASAP7_75t_SL g9495 ( 
.A(n_9189),
.B(n_3594),
.Y(n_9495)
);

NOR2xp33_ASAP7_75t_R g9496 ( 
.A(n_9073),
.B(n_3595),
.Y(n_9496)
);

BUFx3_ASAP7_75t_L g9497 ( 
.A(n_8760),
.Y(n_9497)
);

OAI22xp5_ASAP7_75t_L g9498 ( 
.A1(n_8927),
.A2(n_8976),
.B1(n_9191),
.B2(n_8984),
.Y(n_9498)
);

NAND2xp5_ASAP7_75t_L g9499 ( 
.A(n_9297),
.B(n_250),
.Y(n_9499)
);

AND2x4_ASAP7_75t_L g9500 ( 
.A(n_9236),
.B(n_3597),
.Y(n_9500)
);

NAND2xp5_ASAP7_75t_SL g9501 ( 
.A(n_9177),
.B(n_3598),
.Y(n_9501)
);

BUFx3_ASAP7_75t_L g9502 ( 
.A(n_8775),
.Y(n_9502)
);

AOI21xp5_ASAP7_75t_L g9503 ( 
.A1(n_8931),
.A2(n_3601),
.B(n_3600),
.Y(n_9503)
);

INVx4_ASAP7_75t_L g9504 ( 
.A(n_8877),
.Y(n_9504)
);

INVx1_ASAP7_75t_L g9505 ( 
.A(n_9042),
.Y(n_9505)
);

NAND3xp33_ASAP7_75t_SL g9506 ( 
.A(n_8830),
.B(n_252),
.C(n_253),
.Y(n_9506)
);

INVx1_ASAP7_75t_L g9507 ( 
.A(n_9045),
.Y(n_9507)
);

HB1xp67_ASAP7_75t_L g9508 ( 
.A(n_9079),
.Y(n_9508)
);

BUFx3_ASAP7_75t_L g9509 ( 
.A(n_8883),
.Y(n_9509)
);

NOR2xp33_ASAP7_75t_L g9510 ( 
.A(n_9111),
.B(n_3602),
.Y(n_9510)
);

INVx3_ASAP7_75t_L g9511 ( 
.A(n_9222),
.Y(n_9511)
);

NAND2xp5_ASAP7_75t_SL g9512 ( 
.A(n_9182),
.B(n_3603),
.Y(n_9512)
);

INVx2_ASAP7_75t_L g9513 ( 
.A(n_8852),
.Y(n_9513)
);

INVx1_ASAP7_75t_L g9514 ( 
.A(n_9058),
.Y(n_9514)
);

AOI22xp5_ASAP7_75t_L g9515 ( 
.A1(n_9012),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_9515)
);

HB1xp67_ASAP7_75t_L g9516 ( 
.A(n_9091),
.Y(n_9516)
);

BUFx6f_ASAP7_75t_L g9517 ( 
.A(n_9009),
.Y(n_9517)
);

NAND2xp5_ASAP7_75t_L g9518 ( 
.A(n_9299),
.B(n_255),
.Y(n_9518)
);

BUFx6f_ASAP7_75t_L g9519 ( 
.A(n_9009),
.Y(n_9519)
);

INVx1_ASAP7_75t_L g9520 ( 
.A(n_9086),
.Y(n_9520)
);

INVx2_ASAP7_75t_L g9521 ( 
.A(n_8868),
.Y(n_9521)
);

INVx3_ASAP7_75t_L g9522 ( 
.A(n_9005),
.Y(n_9522)
);

INVx3_ASAP7_75t_L g9523 ( 
.A(n_8811),
.Y(n_9523)
);

OR2x6_ASAP7_75t_L g9524 ( 
.A(n_8871),
.B(n_3604),
.Y(n_9524)
);

INVx1_ASAP7_75t_L g9525 ( 
.A(n_9096),
.Y(n_9525)
);

OAI22xp33_ASAP7_75t_L g9526 ( 
.A1(n_8777),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_9526)
);

INVx2_ASAP7_75t_SL g9527 ( 
.A(n_8892),
.Y(n_9527)
);

AOI22xp33_ASAP7_75t_L g9528 ( 
.A1(n_8762),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_9528)
);

O2A1O1Ixp33_ASAP7_75t_L g9529 ( 
.A1(n_8759),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_9529)
);

BUFx2_ASAP7_75t_L g9530 ( 
.A(n_9091),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_9099),
.Y(n_9531)
);

HB1xp67_ASAP7_75t_L g9532 ( 
.A(n_9053),
.Y(n_9532)
);

AOI22xp33_ASAP7_75t_SL g9533 ( 
.A1(n_9220),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_9533)
);

INVx1_ASAP7_75t_L g9534 ( 
.A(n_9100),
.Y(n_9534)
);

NAND2xp33_ASAP7_75t_L g9535 ( 
.A(n_9220),
.B(n_263),
.Y(n_9535)
);

HB1xp67_ASAP7_75t_L g9536 ( 
.A(n_9097),
.Y(n_9536)
);

NAND2xp5_ASAP7_75t_L g9537 ( 
.A(n_9109),
.B(n_9110),
.Y(n_9537)
);

INVx2_ASAP7_75t_L g9538 ( 
.A(n_8875),
.Y(n_9538)
);

INVx2_ASAP7_75t_SL g9539 ( 
.A(n_8781),
.Y(n_9539)
);

INVx1_ASAP7_75t_L g9540 ( 
.A(n_9104),
.Y(n_9540)
);

AND2x4_ASAP7_75t_L g9541 ( 
.A(n_9292),
.B(n_3605),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_9098),
.Y(n_9542)
);

NAND2xp5_ASAP7_75t_L g9543 ( 
.A(n_9112),
.B(n_9118),
.Y(n_9543)
);

NOR3xp33_ASAP7_75t_SL g9544 ( 
.A(n_9017),
.B(n_263),
.C(n_264),
.Y(n_9544)
);

INVx1_ASAP7_75t_L g9545 ( 
.A(n_9102),
.Y(n_9545)
);

BUFx2_ASAP7_75t_L g9546 ( 
.A(n_9014),
.Y(n_9546)
);

NAND2xp5_ASAP7_75t_L g9547 ( 
.A(n_9126),
.B(n_9135),
.Y(n_9547)
);

AND3x1_ASAP7_75t_SL g9548 ( 
.A(n_9067),
.B(n_264),
.C(n_265),
.Y(n_9548)
);

AND2x2_ASAP7_75t_L g9549 ( 
.A(n_9168),
.B(n_3606),
.Y(n_9549)
);

INVx2_ASAP7_75t_L g9550 ( 
.A(n_8882),
.Y(n_9550)
);

AOI22xp33_ASAP7_75t_L g9551 ( 
.A1(n_9200),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9145),
.Y(n_9552)
);

INVx4_ASAP7_75t_L g9553 ( 
.A(n_8880),
.Y(n_9553)
);

INVx2_ASAP7_75t_L g9554 ( 
.A(n_8885),
.Y(n_9554)
);

INVx5_ASAP7_75t_L g9555 ( 
.A(n_8991),
.Y(n_9555)
);

OR2x6_ASAP7_75t_L g9556 ( 
.A(n_8871),
.B(n_3607),
.Y(n_9556)
);

BUFx12f_ASAP7_75t_L g9557 ( 
.A(n_8924),
.Y(n_9557)
);

NAND2xp5_ASAP7_75t_L g9558 ( 
.A(n_9142),
.B(n_266),
.Y(n_9558)
);

OAI22xp33_ASAP7_75t_L g9559 ( 
.A1(n_8866),
.A2(n_9291),
.B1(n_9276),
.B2(n_8911),
.Y(n_9559)
);

BUFx4f_ASAP7_75t_L g9560 ( 
.A(n_8991),
.Y(n_9560)
);

A2O1A1Ixp33_ASAP7_75t_L g9561 ( 
.A1(n_8712),
.A2(n_270),
.B(n_267),
.C(n_269),
.Y(n_9561)
);

BUFx8_ASAP7_75t_L g9562 ( 
.A(n_8935),
.Y(n_9562)
);

INVx3_ASAP7_75t_L g9563 ( 
.A(n_9293),
.Y(n_9563)
);

INVx3_ASAP7_75t_L g9564 ( 
.A(n_8817),
.Y(n_9564)
);

AND3x1_ASAP7_75t_SL g9565 ( 
.A(n_9153),
.B(n_269),
.C(n_270),
.Y(n_9565)
);

BUFx12f_ASAP7_75t_L g9566 ( 
.A(n_8983),
.Y(n_9566)
);

NAND2xp5_ASAP7_75t_L g9567 ( 
.A(n_9144),
.B(n_271),
.Y(n_9567)
);

INVx2_ASAP7_75t_L g9568 ( 
.A(n_9202),
.Y(n_9568)
);

BUFx4_ASAP7_75t_SL g9569 ( 
.A(n_8944),
.Y(n_9569)
);

AND2x2_ASAP7_75t_L g9570 ( 
.A(n_9027),
.B(n_3608),
.Y(n_9570)
);

NOR3xp33_ASAP7_75t_SL g9571 ( 
.A(n_9004),
.B(n_271),
.C(n_272),
.Y(n_9571)
);

INVx1_ASAP7_75t_L g9572 ( 
.A(n_8737),
.Y(n_9572)
);

INVx1_ASAP7_75t_L g9573 ( 
.A(n_8744),
.Y(n_9573)
);

INVx3_ASAP7_75t_L g9574 ( 
.A(n_8900),
.Y(n_9574)
);

INVx3_ASAP7_75t_L g9575 ( 
.A(n_8941),
.Y(n_9575)
);

INVx3_ASAP7_75t_L g9576 ( 
.A(n_8708),
.Y(n_9576)
);

NAND2xp33_ASAP7_75t_SL g9577 ( 
.A(n_9213),
.B(n_9254),
.Y(n_9577)
);

INVx2_ASAP7_75t_SL g9578 ( 
.A(n_8805),
.Y(n_9578)
);

INVx1_ASAP7_75t_SL g9579 ( 
.A(n_8829),
.Y(n_9579)
);

NOR3xp33_ASAP7_75t_SL g9580 ( 
.A(n_9156),
.B(n_272),
.C(n_273),
.Y(n_9580)
);

CKINVDCx5p33_ASAP7_75t_R g9581 ( 
.A(n_9185),
.Y(n_9581)
);

NAND2xp5_ASAP7_75t_SL g9582 ( 
.A(n_8984),
.B(n_3610),
.Y(n_9582)
);

BUFx2_ASAP7_75t_L g9583 ( 
.A(n_9076),
.Y(n_9583)
);

INVx1_ASAP7_75t_L g9584 ( 
.A(n_8761),
.Y(n_9584)
);

INVx1_ASAP7_75t_L g9585 ( 
.A(n_8785),
.Y(n_9585)
);

NOR2xp33_ASAP7_75t_L g9586 ( 
.A(n_9031),
.B(n_3611),
.Y(n_9586)
);

INVx5_ASAP7_75t_L g9587 ( 
.A(n_9056),
.Y(n_9587)
);

NAND2xp5_ASAP7_75t_L g9588 ( 
.A(n_9062),
.B(n_274),
.Y(n_9588)
);

OR2x2_ASAP7_75t_L g9589 ( 
.A(n_8786),
.B(n_275),
.Y(n_9589)
);

NAND2xp5_ASAP7_75t_L g9590 ( 
.A(n_9161),
.B(n_275),
.Y(n_9590)
);

INVx3_ASAP7_75t_L g9591 ( 
.A(n_9209),
.Y(n_9591)
);

INVx1_ASAP7_75t_L g9592 ( 
.A(n_8791),
.Y(n_9592)
);

AND2x2_ASAP7_75t_L g9593 ( 
.A(n_9171),
.B(n_3612),
.Y(n_9593)
);

BUFx6f_ASAP7_75t_L g9594 ( 
.A(n_8983),
.Y(n_9594)
);

NOR2xp33_ASAP7_75t_L g9595 ( 
.A(n_9181),
.B(n_3614),
.Y(n_9595)
);

NAND2xp5_ASAP7_75t_SL g9596 ( 
.A(n_9149),
.B(n_3616),
.Y(n_9596)
);

NOR2xp33_ASAP7_75t_L g9597 ( 
.A(n_8989),
.B(n_9230),
.Y(n_9597)
);

NAND2xp5_ASAP7_75t_L g9598 ( 
.A(n_9163),
.B(n_276),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_9215),
.Y(n_9599)
);

BUFx6f_ASAP7_75t_L g9600 ( 
.A(n_9300),
.Y(n_9600)
);

AOI22xp5_ASAP7_75t_L g9601 ( 
.A1(n_8796),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_9601)
);

BUFx3_ASAP7_75t_L g9602 ( 
.A(n_8913),
.Y(n_9602)
);

CKINVDCx5p33_ASAP7_75t_R g9603 ( 
.A(n_8966),
.Y(n_9603)
);

INVx2_ASAP7_75t_SL g9604 ( 
.A(n_8936),
.Y(n_9604)
);

HB1xp67_ASAP7_75t_L g9605 ( 
.A(n_8793),
.Y(n_9605)
);

CKINVDCx20_ASAP7_75t_R g9606 ( 
.A(n_9294),
.Y(n_9606)
);

INVx1_ASAP7_75t_L g9607 ( 
.A(n_8801),
.Y(n_9607)
);

NAND3xp33_ASAP7_75t_SL g9608 ( 
.A(n_8818),
.B(n_277),
.C(n_278),
.Y(n_9608)
);

INVx1_ASAP7_75t_L g9609 ( 
.A(n_8804),
.Y(n_9609)
);

INVx1_ASAP7_75t_L g9610 ( 
.A(n_8815),
.Y(n_9610)
);

BUFx2_ASAP7_75t_L g9611 ( 
.A(n_9157),
.Y(n_9611)
);

NAND2xp5_ASAP7_75t_L g9612 ( 
.A(n_9172),
.B(n_279),
.Y(n_9612)
);

INVx3_ASAP7_75t_L g9613 ( 
.A(n_9216),
.Y(n_9613)
);

BUFx3_ASAP7_75t_L g9614 ( 
.A(n_8952),
.Y(n_9614)
);

OR2x2_ASAP7_75t_SL g9615 ( 
.A(n_8808),
.B(n_279),
.Y(n_9615)
);

OR2x6_ASAP7_75t_L g9616 ( 
.A(n_8770),
.B(n_3617),
.Y(n_9616)
);

AOI22xp33_ASAP7_75t_L g9617 ( 
.A1(n_9050),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_9617)
);

NOR2xp33_ASAP7_75t_R g9618 ( 
.A(n_9046),
.B(n_3618),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_8820),
.Y(n_9619)
);

INVx2_ASAP7_75t_L g9620 ( 
.A(n_9217),
.Y(n_9620)
);

INVx1_ASAP7_75t_L g9621 ( 
.A(n_8823),
.Y(n_9621)
);

AND2x6_ASAP7_75t_SL g9622 ( 
.A(n_8919),
.B(n_280),
.Y(n_9622)
);

BUFx6f_ASAP7_75t_L g9623 ( 
.A(n_9223),
.Y(n_9623)
);

INVx2_ASAP7_75t_L g9624 ( 
.A(n_9238),
.Y(n_9624)
);

BUFx6f_ASAP7_75t_L g9625 ( 
.A(n_9226),
.Y(n_9625)
);

INVx2_ASAP7_75t_L g9626 ( 
.A(n_9243),
.Y(n_9626)
);

AND2x2_ASAP7_75t_L g9627 ( 
.A(n_9180),
.B(n_9154),
.Y(n_9627)
);

AOI211xp5_ASAP7_75t_L g9628 ( 
.A1(n_8788),
.A2(n_8993),
.B(n_9008),
.C(n_9003),
.Y(n_9628)
);

INVx3_ASAP7_75t_SL g9629 ( 
.A(n_8880),
.Y(n_9629)
);

NAND2xp5_ASAP7_75t_L g9630 ( 
.A(n_9178),
.B(n_281),
.Y(n_9630)
);

HB1xp67_ASAP7_75t_L g9631 ( 
.A(n_8825),
.Y(n_9631)
);

INVx2_ASAP7_75t_SL g9632 ( 
.A(n_9278),
.Y(n_9632)
);

INVx2_ASAP7_75t_L g9633 ( 
.A(n_9244),
.Y(n_9633)
);

OAI21x1_ASAP7_75t_L g9634 ( 
.A1(n_9164),
.A2(n_9184),
.B(n_9094),
.Y(n_9634)
);

BUFx6f_ASAP7_75t_L g9635 ( 
.A(n_9157),
.Y(n_9635)
);

INVxp67_ASAP7_75t_SL g9636 ( 
.A(n_9249),
.Y(n_9636)
);

AND2x4_ASAP7_75t_L g9637 ( 
.A(n_8854),
.B(n_3619),
.Y(n_9637)
);

NOR3xp33_ASAP7_75t_SL g9638 ( 
.A(n_8827),
.B(n_282),
.C(n_283),
.Y(n_9638)
);

INVx3_ASAP7_75t_SL g9639 ( 
.A(n_9158),
.Y(n_9639)
);

INVx4_ASAP7_75t_L g9640 ( 
.A(n_8806),
.Y(n_9640)
);

NAND2xp5_ASAP7_75t_SL g9641 ( 
.A(n_9260),
.B(n_9288),
.Y(n_9641)
);

INVxp67_ASAP7_75t_SL g9642 ( 
.A(n_9253),
.Y(n_9642)
);

NAND2xp5_ASAP7_75t_L g9643 ( 
.A(n_9179),
.B(n_9187),
.Y(n_9643)
);

NAND2xp5_ASAP7_75t_L g9644 ( 
.A(n_9150),
.B(n_283),
.Y(n_9644)
);

OR2x6_ASAP7_75t_L g9645 ( 
.A(n_8770),
.B(n_3620),
.Y(n_9645)
);

BUFx3_ASAP7_75t_L g9646 ( 
.A(n_9158),
.Y(n_9646)
);

AND2x2_ASAP7_75t_L g9647 ( 
.A(n_8784),
.B(n_3621),
.Y(n_9647)
);

BUFx6f_ASAP7_75t_L g9648 ( 
.A(n_8717),
.Y(n_9648)
);

AND2x4_ASAP7_75t_L g9649 ( 
.A(n_8764),
.B(n_3623),
.Y(n_9649)
);

INVx2_ASAP7_75t_L g9650 ( 
.A(n_9263),
.Y(n_9650)
);

AND2x4_ASAP7_75t_L g9651 ( 
.A(n_9056),
.B(n_3624),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_9060),
.Y(n_9652)
);

NOR3xp33_ASAP7_75t_SL g9653 ( 
.A(n_8960),
.B(n_8765),
.C(n_8816),
.Y(n_9653)
);

INVx1_ASAP7_75t_L g9654 ( 
.A(n_9264),
.Y(n_9654)
);

BUFx3_ASAP7_75t_L g9655 ( 
.A(n_8949),
.Y(n_9655)
);

INVx1_ASAP7_75t_L g9656 ( 
.A(n_9266),
.Y(n_9656)
);

NAND3xp33_ASAP7_75t_SL g9657 ( 
.A(n_8884),
.B(n_285),
.C(n_286),
.Y(n_9657)
);

INVx2_ASAP7_75t_L g9658 ( 
.A(n_9280),
.Y(n_9658)
);

AOI21xp5_ASAP7_75t_L g9659 ( 
.A1(n_8996),
.A2(n_3626),
.B(n_3625),
.Y(n_9659)
);

NAND2xp5_ASAP7_75t_L g9660 ( 
.A(n_9095),
.B(n_285),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_9298),
.Y(n_9661)
);

INVx2_ASAP7_75t_L g9662 ( 
.A(n_9284),
.Y(n_9662)
);

BUFx3_ASAP7_75t_L g9663 ( 
.A(n_8896),
.Y(n_9663)
);

INVx2_ASAP7_75t_SL g9664 ( 
.A(n_8897),
.Y(n_9664)
);

INVx1_ASAP7_75t_L g9665 ( 
.A(n_9287),
.Y(n_9665)
);

OR2x6_ASAP7_75t_L g9666 ( 
.A(n_8763),
.B(n_8954),
.Y(n_9666)
);

NAND2xp5_ASAP7_75t_SL g9667 ( 
.A(n_9006),
.B(n_3627),
.Y(n_9667)
);

NAND2xp5_ASAP7_75t_SL g9668 ( 
.A(n_9020),
.B(n_3630),
.Y(n_9668)
);

NOR2xp33_ASAP7_75t_L g9669 ( 
.A(n_8974),
.B(n_3631),
.Y(n_9669)
);

CKINVDCx20_ASAP7_75t_R g9670 ( 
.A(n_9277),
.Y(n_9670)
);

NOR3xp33_ASAP7_75t_SL g9671 ( 
.A(n_9001),
.B(n_287),
.C(n_288),
.Y(n_9671)
);

OAI21xp33_ASAP7_75t_L g9672 ( 
.A1(n_9033),
.A2(n_288),
.B(n_289),
.Y(n_9672)
);

INVx2_ASAP7_75t_L g9673 ( 
.A(n_9285),
.Y(n_9673)
);

OAI22xp33_ASAP7_75t_L g9674 ( 
.A1(n_9029),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_9674)
);

INVx1_ASAP7_75t_L g9675 ( 
.A(n_9080),
.Y(n_9675)
);

AND2x4_ASAP7_75t_L g9676 ( 
.A(n_9063),
.B(n_9055),
.Y(n_9676)
);

INVx1_ASAP7_75t_L g9677 ( 
.A(n_9080),
.Y(n_9677)
);

OR2x6_ASAP7_75t_L g9678 ( 
.A(n_8763),
.B(n_291),
.Y(n_9678)
);

NAND2xp5_ASAP7_75t_L g9679 ( 
.A(n_9167),
.B(n_292),
.Y(n_9679)
);

INVx2_ASAP7_75t_SL g9680 ( 
.A(n_8909),
.Y(n_9680)
);

AOI22xp33_ASAP7_75t_L g9681 ( 
.A1(n_8916),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_9681)
);

INVx1_ASAP7_75t_L g9682 ( 
.A(n_9080),
.Y(n_9682)
);

INVx2_ASAP7_75t_L g9683 ( 
.A(n_8888),
.Y(n_9683)
);

BUFx6f_ASAP7_75t_L g9684 ( 
.A(n_9089),
.Y(n_9684)
);

BUFx2_ASAP7_75t_L g9685 ( 
.A(n_9130),
.Y(n_9685)
);

INVx1_ASAP7_75t_L g9686 ( 
.A(n_8899),
.Y(n_9686)
);

INVx1_ASAP7_75t_L g9687 ( 
.A(n_8903),
.Y(n_9687)
);

NAND2xp5_ASAP7_75t_L g9688 ( 
.A(n_8742),
.B(n_293),
.Y(n_9688)
);

INVx2_ASAP7_75t_L g9689 ( 
.A(n_8908),
.Y(n_9689)
);

NAND2xp5_ASAP7_75t_L g9690 ( 
.A(n_9138),
.B(n_9231),
.Y(n_9690)
);

INVx3_ASAP7_75t_L g9691 ( 
.A(n_9089),
.Y(n_9691)
);

NAND2xp5_ASAP7_75t_SL g9692 ( 
.A(n_9198),
.B(n_295),
.Y(n_9692)
);

INVx3_ASAP7_75t_L g9693 ( 
.A(n_8928),
.Y(n_9693)
);

NOR2xp33_ASAP7_75t_R g9694 ( 
.A(n_9169),
.B(n_297),
.Y(n_9694)
);

CKINVDCx5p33_ASAP7_75t_R g9695 ( 
.A(n_9038),
.Y(n_9695)
);

AOI22xp33_ASAP7_75t_SL g9696 ( 
.A1(n_9286),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_9696)
);

NOR3xp33_ASAP7_75t_SL g9697 ( 
.A(n_9170),
.B(n_298),
.C(n_299),
.Y(n_9697)
);

INVx1_ASAP7_75t_L g9698 ( 
.A(n_8917),
.Y(n_9698)
);

INVx1_ASAP7_75t_L g9699 ( 
.A(n_8920),
.Y(n_9699)
);

OAI22xp5_ASAP7_75t_L g9700 ( 
.A1(n_9198),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_9700)
);

NAND2xp5_ASAP7_75t_SL g9701 ( 
.A(n_9019),
.B(n_9194),
.Y(n_9701)
);

NAND2xp5_ASAP7_75t_L g9702 ( 
.A(n_9232),
.B(n_9234),
.Y(n_9702)
);

BUFx3_ASAP7_75t_L g9703 ( 
.A(n_8824),
.Y(n_9703)
);

NOR2xp67_ASAP7_75t_L g9704 ( 
.A(n_9070),
.B(n_300),
.Y(n_9704)
);

INVx4_ASAP7_75t_L g9705 ( 
.A(n_9055),
.Y(n_9705)
);

INVx1_ASAP7_75t_L g9706 ( 
.A(n_8942),
.Y(n_9706)
);

BUFx12f_ASAP7_75t_L g9707 ( 
.A(n_8930),
.Y(n_9707)
);

CKINVDCx16_ASAP7_75t_R g9708 ( 
.A(n_8975),
.Y(n_9708)
);

INVx4_ASAP7_75t_L g9709 ( 
.A(n_8930),
.Y(n_9709)
);

NOR2xp33_ASAP7_75t_R g9710 ( 
.A(n_9186),
.B(n_301),
.Y(n_9710)
);

NOR2xp33_ASAP7_75t_L g9711 ( 
.A(n_9069),
.B(n_303),
.Y(n_9711)
);

AND2x2_ASAP7_75t_L g9712 ( 
.A(n_8886),
.B(n_303),
.Y(n_9712)
);

NAND2x1p5_ASAP7_75t_L g9713 ( 
.A(n_9152),
.B(n_304),
.Y(n_9713)
);

INVxp67_ASAP7_75t_L g9714 ( 
.A(n_8789),
.Y(n_9714)
);

NAND2xp5_ASAP7_75t_L g9715 ( 
.A(n_9237),
.B(n_9258),
.Y(n_9715)
);

CKINVDCx5p33_ASAP7_75t_R g9716 ( 
.A(n_8771),
.Y(n_9716)
);

INVx2_ASAP7_75t_SL g9717 ( 
.A(n_8950),
.Y(n_9717)
);

OR2x2_ASAP7_75t_L g9718 ( 
.A(n_8723),
.B(n_304),
.Y(n_9718)
);

AO22x1_ASAP7_75t_L g9719 ( 
.A1(n_9220),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_9719)
);

NAND2xp5_ASAP7_75t_SL g9720 ( 
.A(n_9175),
.B(n_305),
.Y(n_9720)
);

AND2x2_ASAP7_75t_L g9721 ( 
.A(n_8937),
.B(n_306),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_8969),
.Y(n_9722)
);

BUFx8_ASAP7_75t_SL g9723 ( 
.A(n_8948),
.Y(n_9723)
);

BUFx6f_ASAP7_75t_L g9724 ( 
.A(n_8981),
.Y(n_9724)
);

INVx1_ASAP7_75t_SL g9725 ( 
.A(n_8958),
.Y(n_9725)
);

INVx1_ASAP7_75t_SL g9726 ( 
.A(n_8995),
.Y(n_9726)
);

BUFx3_ASAP7_75t_L g9727 ( 
.A(n_9121),
.Y(n_9727)
);

BUFx6f_ASAP7_75t_L g9728 ( 
.A(n_8988),
.Y(n_9728)
);

INVx2_ASAP7_75t_L g9729 ( 
.A(n_8990),
.Y(n_9729)
);

BUFx3_ASAP7_75t_L g9730 ( 
.A(n_8994),
.Y(n_9730)
);

NOR2xp33_ASAP7_75t_L g9731 ( 
.A(n_8813),
.B(n_307),
.Y(n_9731)
);

AOI22xp5_ASAP7_75t_L g9732 ( 
.A1(n_8734),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_9732)
);

NOR2xp33_ASAP7_75t_SL g9733 ( 
.A(n_9286),
.B(n_308),
.Y(n_9733)
);

NOR3xp33_ASAP7_75t_SL g9734 ( 
.A(n_8834),
.B(n_309),
.C(n_311),
.Y(n_9734)
);

NAND2xp5_ASAP7_75t_L g9735 ( 
.A(n_9267),
.B(n_311),
.Y(n_9735)
);

INVx2_ASAP7_75t_L g9736 ( 
.A(n_9000),
.Y(n_9736)
);

NAND2xp5_ASAP7_75t_L g9737 ( 
.A(n_9269),
.B(n_312),
.Y(n_9737)
);

NOR3xp33_ASAP7_75t_SL g9738 ( 
.A(n_8992),
.B(n_312),
.C(n_313),
.Y(n_9738)
);

AND3x1_ASAP7_75t_SL g9739 ( 
.A(n_9282),
.B(n_313),
.C(n_314),
.Y(n_9739)
);

AND2x6_ASAP7_75t_SL g9740 ( 
.A(n_9002),
.B(n_315),
.Y(n_9740)
);

CKINVDCx5p33_ASAP7_75t_R g9741 ( 
.A(n_8912),
.Y(n_9741)
);

INVx1_ASAP7_75t_L g9742 ( 
.A(n_9064),
.Y(n_9742)
);

NAND2xp5_ASAP7_75t_L g9743 ( 
.A(n_9270),
.B(n_315),
.Y(n_9743)
);

AND2x4_ASAP7_75t_L g9744 ( 
.A(n_9119),
.B(n_316),
.Y(n_9744)
);

INVx2_ASAP7_75t_SL g9745 ( 
.A(n_9239),
.Y(n_9745)
);

INVx2_ASAP7_75t_L g9746 ( 
.A(n_9125),
.Y(n_9746)
);

BUFx2_ASAP7_75t_L g9747 ( 
.A(n_9286),
.Y(n_9747)
);

INVx1_ASAP7_75t_L g9748 ( 
.A(n_9125),
.Y(n_9748)
);

NAND2xp5_ASAP7_75t_L g9749 ( 
.A(n_8766),
.B(n_316),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_9052),
.Y(n_9750)
);

INVx1_ASAP7_75t_L g9751 ( 
.A(n_9057),
.Y(n_9751)
);

AND2x2_ASAP7_75t_L g9752 ( 
.A(n_9195),
.B(n_9083),
.Y(n_9752)
);

INVx2_ASAP7_75t_SL g9753 ( 
.A(n_9034),
.Y(n_9753)
);

NAND2xp5_ASAP7_75t_L g9754 ( 
.A(n_8780),
.B(n_317),
.Y(n_9754)
);

INVx2_ASAP7_75t_L g9755 ( 
.A(n_9120),
.Y(n_9755)
);

INVx3_ASAP7_75t_SL g9756 ( 
.A(n_9162),
.Y(n_9756)
);

NAND2xp5_ASAP7_75t_L g9757 ( 
.A(n_8790),
.B(n_8794),
.Y(n_9757)
);

INVx1_ASAP7_75t_L g9758 ( 
.A(n_9082),
.Y(n_9758)
);

BUFx6f_ASAP7_75t_L g9759 ( 
.A(n_9116),
.Y(n_9759)
);

CKINVDCx11_ASAP7_75t_R g9760 ( 
.A(n_9119),
.Y(n_9760)
);

BUFx12f_ASAP7_75t_L g9761 ( 
.A(n_8835),
.Y(n_9761)
);

NAND2xp5_ASAP7_75t_L g9762 ( 
.A(n_8798),
.B(n_317),
.Y(n_9762)
);

NAND2xp5_ASAP7_75t_L g9763 ( 
.A(n_8800),
.B(n_318),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_9122),
.Y(n_9764)
);

INVx1_ASAP7_75t_L g9765 ( 
.A(n_9134),
.Y(n_9765)
);

CKINVDCx5p33_ASAP7_75t_R g9766 ( 
.A(n_9174),
.Y(n_9766)
);

INVx2_ASAP7_75t_L g9767 ( 
.A(n_9140),
.Y(n_9767)
);

NOR2xp33_ASAP7_75t_SL g9768 ( 
.A(n_9147),
.B(n_318),
.Y(n_9768)
);

INVx1_ASAP7_75t_L g9769 ( 
.A(n_9024),
.Y(n_9769)
);

NAND2xp5_ASAP7_75t_L g9770 ( 
.A(n_8807),
.B(n_8810),
.Y(n_9770)
);

AND2x4_ASAP7_75t_L g9771 ( 
.A(n_8867),
.B(n_319),
.Y(n_9771)
);

INVx2_ASAP7_75t_L g9772 ( 
.A(n_9041),
.Y(n_9772)
);

NOR2xp33_ASAP7_75t_L g9773 ( 
.A(n_8738),
.B(n_8977),
.Y(n_9773)
);

BUFx6f_ASAP7_75t_L g9774 ( 
.A(n_9127),
.Y(n_9774)
);

BUFx2_ASAP7_75t_L g9775 ( 
.A(n_9132),
.Y(n_9775)
);

NOR3xp33_ASAP7_75t_SL g9776 ( 
.A(n_9081),
.B(n_319),
.C(n_320),
.Y(n_9776)
);

INVx2_ASAP7_75t_L g9777 ( 
.A(n_9049),
.Y(n_9777)
);

A2O1A1Ixp33_ASAP7_75t_L g9778 ( 
.A1(n_9159),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_9778)
);

INVx1_ASAP7_75t_L g9779 ( 
.A(n_8726),
.Y(n_9779)
);

INVx1_ASAP7_75t_L g9780 ( 
.A(n_8947),
.Y(n_9780)
);

BUFx3_ASAP7_75t_L g9781 ( 
.A(n_8956),
.Y(n_9781)
);

NAND2xp5_ASAP7_75t_L g9782 ( 
.A(n_8768),
.B(n_321),
.Y(n_9782)
);

BUFx2_ASAP7_75t_SL g9783 ( 
.A(n_9251),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9025),
.Y(n_9784)
);

INVx2_ASAP7_75t_SL g9785 ( 
.A(n_8967),
.Y(n_9785)
);

INVx2_ASAP7_75t_L g9786 ( 
.A(n_9196),
.Y(n_9786)
);

NAND2xp5_ASAP7_75t_L g9787 ( 
.A(n_9047),
.B(n_322),
.Y(n_9787)
);

BUFx3_ASAP7_75t_L g9788 ( 
.A(n_8821),
.Y(n_9788)
);

BUFx3_ASAP7_75t_L g9789 ( 
.A(n_8828),
.Y(n_9789)
);

BUFx6f_ASAP7_75t_L g9790 ( 
.A(n_9129),
.Y(n_9790)
);

INVx2_ASAP7_75t_L g9791 ( 
.A(n_8921),
.Y(n_9791)
);

INVx1_ASAP7_75t_L g9792 ( 
.A(n_8822),
.Y(n_9792)
);

INVx2_ASAP7_75t_L g9793 ( 
.A(n_9051),
.Y(n_9793)
);

AND3x1_ASAP7_75t_SL g9794 ( 
.A(n_8951),
.B(n_323),
.C(n_324),
.Y(n_9794)
);

INVx4_ASAP7_75t_L g9795 ( 
.A(n_8872),
.Y(n_9795)
);

INVx2_ASAP7_75t_L g9796 ( 
.A(n_9115),
.Y(n_9796)
);

NAND2xp5_ASAP7_75t_L g9797 ( 
.A(n_8739),
.B(n_324),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_9204),
.Y(n_9798)
);

OAI21xp5_ASAP7_75t_L g9799 ( 
.A1(n_8842),
.A2(n_325),
.B(n_326),
.Y(n_9799)
);

NAND2xp5_ASAP7_75t_L g9800 ( 
.A(n_8922),
.B(n_325),
.Y(n_9800)
);

INVx1_ASAP7_75t_L g9801 ( 
.A(n_9085),
.Y(n_9801)
);

INVx1_ASAP7_75t_SL g9802 ( 
.A(n_8756),
.Y(n_9802)
);

NAND2xp5_ASAP7_75t_L g9803 ( 
.A(n_8933),
.B(n_326),
.Y(n_9803)
);

HB1xp67_ASAP7_75t_L g9804 ( 
.A(n_9148),
.Y(n_9804)
);

AND2x4_ASAP7_75t_L g9805 ( 
.A(n_9273),
.B(n_327),
.Y(n_9805)
);

BUFx2_ASAP7_75t_L g9806 ( 
.A(n_8872),
.Y(n_9806)
);

INVx4_ASAP7_75t_L g9807 ( 
.A(n_9208),
.Y(n_9807)
);

INVx2_ASAP7_75t_L g9808 ( 
.A(n_9123),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_9087),
.Y(n_9809)
);

NAND2xp5_ASAP7_75t_L g9810 ( 
.A(n_8745),
.B(n_327),
.Y(n_9810)
);

NAND2xp5_ASAP7_75t_L g9811 ( 
.A(n_8748),
.B(n_328),
.Y(n_9811)
);

INVx3_ASAP7_75t_L g9812 ( 
.A(n_8819),
.Y(n_9812)
);

CKINVDCx5p33_ASAP7_75t_R g9813 ( 
.A(n_8795),
.Y(n_9813)
);

HB1xp67_ASAP7_75t_L g9814 ( 
.A(n_9192),
.Y(n_9814)
);

INVx2_ASAP7_75t_L g9815 ( 
.A(n_9128),
.Y(n_9815)
);

INVx2_ASAP7_75t_SL g9816 ( 
.A(n_8847),
.Y(n_9816)
);

NOR2xp33_ASAP7_75t_L g9817 ( 
.A(n_9023),
.B(n_328),
.Y(n_9817)
);

AND2x2_ASAP7_75t_L g9818 ( 
.A(n_9188),
.B(n_329),
.Y(n_9818)
);

INVx2_ASAP7_75t_SL g9819 ( 
.A(n_8986),
.Y(n_9819)
);

INVx1_ASAP7_75t_L g9820 ( 
.A(n_9092),
.Y(n_9820)
);

BUFx4f_ASAP7_75t_L g9821 ( 
.A(n_9199),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_9108),
.Y(n_9822)
);

NAND2xp5_ASAP7_75t_L g9823 ( 
.A(n_8751),
.B(n_329),
.Y(n_9823)
);

NAND2xp5_ASAP7_75t_SL g9824 ( 
.A(n_9131),
.B(n_330),
.Y(n_9824)
);

INVx5_ASAP7_75t_L g9825 ( 
.A(n_9113),
.Y(n_9825)
);

AND2x2_ASAP7_75t_L g9826 ( 
.A(n_9133),
.B(n_332),
.Y(n_9826)
);

BUFx3_ASAP7_75t_L g9827 ( 
.A(n_9078),
.Y(n_9827)
);

NOR2xp33_ASAP7_75t_L g9828 ( 
.A(n_8836),
.B(n_332),
.Y(n_9828)
);

INVx2_ASAP7_75t_L g9829 ( 
.A(n_9136),
.Y(n_9829)
);

INVx2_ASAP7_75t_SL g9830 ( 
.A(n_8846),
.Y(n_9830)
);

BUFx12f_ASAP7_75t_L g9831 ( 
.A(n_9105),
.Y(n_9831)
);

NAND2xp5_ASAP7_75t_L g9832 ( 
.A(n_8773),
.B(n_333),
.Y(n_9832)
);

INVx2_ASAP7_75t_L g9833 ( 
.A(n_9141),
.Y(n_9833)
);

AOI22xp5_ASAP7_75t_L g9834 ( 
.A1(n_9013),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_9834)
);

NAND2xp5_ASAP7_75t_L g9835 ( 
.A(n_8879),
.B(n_334),
.Y(n_9835)
);

NOR2xp33_ASAP7_75t_L g9836 ( 
.A(n_9068),
.B(n_335),
.Y(n_9836)
);

BUFx2_ASAP7_75t_L g9837 ( 
.A(n_9176),
.Y(n_9837)
);

NAND2xp5_ASAP7_75t_SL g9838 ( 
.A(n_9160),
.B(n_336),
.Y(n_9838)
);

BUFx3_ASAP7_75t_L g9839 ( 
.A(n_9151),
.Y(n_9839)
);

INVx1_ASAP7_75t_L g9840 ( 
.A(n_9272),
.Y(n_9840)
);

NAND2xp5_ASAP7_75t_L g9841 ( 
.A(n_8891),
.B(n_336),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_9190),
.Y(n_9842)
);

NAND2xp5_ASAP7_75t_L g9843 ( 
.A(n_8905),
.B(n_337),
.Y(n_9843)
);

NOR2xp33_ASAP7_75t_L g9844 ( 
.A(n_8873),
.B(n_337),
.Y(n_9844)
);

NAND2xp33_ASAP7_75t_R g9845 ( 
.A(n_8945),
.B(n_338),
.Y(n_9845)
);

NAND2xp5_ASAP7_75t_L g9846 ( 
.A(n_8906),
.B(n_338),
.Y(n_9846)
);

NOR2xp33_ASAP7_75t_R g9847 ( 
.A(n_9007),
.B(n_9173),
.Y(n_9847)
);

BUFx6f_ASAP7_75t_L g9848 ( 
.A(n_9166),
.Y(n_9848)
);

NAND2xp5_ASAP7_75t_SL g9849 ( 
.A(n_8914),
.B(n_339),
.Y(n_9849)
);

NAND2xp5_ASAP7_75t_L g9850 ( 
.A(n_8833),
.B(n_339),
.Y(n_9850)
);

NAND2xp33_ASAP7_75t_L g9851 ( 
.A(n_9044),
.B(n_340),
.Y(n_9851)
);

INVx1_ASAP7_75t_L g9852 ( 
.A(n_8843),
.Y(n_9852)
);

NAND2xp5_ASAP7_75t_L g9853 ( 
.A(n_8844),
.B(n_341),
.Y(n_9853)
);

OR2x2_ASAP7_75t_L g9854 ( 
.A(n_8850),
.B(n_8957),
.Y(n_9854)
);

NAND2xp5_ASAP7_75t_L g9855 ( 
.A(n_9137),
.B(n_341),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_9037),
.Y(n_9856)
);

BUFx6f_ASAP7_75t_L g9857 ( 
.A(n_9066),
.Y(n_9857)
);

AND2x2_ASAP7_75t_L g9858 ( 
.A(n_8746),
.B(n_342),
.Y(n_9858)
);

NAND2xp33_ASAP7_75t_SL g9859 ( 
.A(n_8894),
.B(n_342),
.Y(n_9859)
);

HB1xp67_ASAP7_75t_L g9860 ( 
.A(n_8982),
.Y(n_9860)
);

NOR2xp33_ASAP7_75t_R g9861 ( 
.A(n_9035),
.B(n_343),
.Y(n_9861)
);

AND2x4_ASAP7_75t_L g9862 ( 
.A(n_8963),
.B(n_344),
.Y(n_9862)
);

BUFx6f_ASAP7_75t_L g9863 ( 
.A(n_8999),
.Y(n_9863)
);

BUFx2_ASAP7_75t_L g9864 ( 
.A(n_8845),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9143),
.Y(n_9865)
);

NAND2xp5_ASAP7_75t_SL g9866 ( 
.A(n_9048),
.B(n_344),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_8878),
.Y(n_9867)
);

BUFx2_ASAP7_75t_L g9868 ( 
.A(n_8814),
.Y(n_9868)
);

INVx3_ASAP7_75t_L g9869 ( 
.A(n_9088),
.Y(n_9869)
);

INVx1_ASAP7_75t_SL g9870 ( 
.A(n_8862),
.Y(n_9870)
);

BUFx6f_ASAP7_75t_L g9871 ( 
.A(n_8898),
.Y(n_9871)
);

NAND2xp5_ASAP7_75t_SL g9872 ( 
.A(n_9015),
.B(n_345),
.Y(n_9872)
);

BUFx6f_ASAP7_75t_L g9873 ( 
.A(n_8876),
.Y(n_9873)
);

AOI22xp5_ASAP7_75t_L g9874 ( 
.A1(n_9183),
.A2(n_349),
.B1(n_345),
.B2(n_346),
.Y(n_9874)
);

AND2x2_ASAP7_75t_L g9875 ( 
.A(n_8743),
.B(n_346),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_9124),
.Y(n_9876)
);

NAND2xp5_ASAP7_75t_L g9877 ( 
.A(n_8731),
.B(n_349),
.Y(n_9877)
);

BUFx2_ASAP7_75t_L g9878 ( 
.A(n_9117),
.Y(n_9878)
);

OR2x6_ASAP7_75t_L g9879 ( 
.A(n_9018),
.B(n_351),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_8857),
.Y(n_9880)
);

CKINVDCx20_ASAP7_75t_R g9881 ( 
.A(n_8997),
.Y(n_9881)
);

CKINVDCx5p33_ASAP7_75t_R g9882 ( 
.A(n_9165),
.Y(n_9882)
);

CKINVDCx5p33_ASAP7_75t_R g9883 ( 
.A(n_9274),
.Y(n_9883)
);

NAND2xp5_ASAP7_75t_L g9884 ( 
.A(n_9252),
.B(n_352),
.Y(n_9884)
);

BUFx3_ASAP7_75t_L g9885 ( 
.A(n_8971),
.Y(n_9885)
);

BUFx6f_ASAP7_75t_L g9886 ( 
.A(n_9257),
.Y(n_9886)
);

AND2x2_ASAP7_75t_L g9887 ( 
.A(n_9265),
.B(n_353),
.Y(n_9887)
);

INVx4_ASAP7_75t_L g9888 ( 
.A(n_8955),
.Y(n_9888)
);

INVxp67_ASAP7_75t_L g9889 ( 
.A(n_8841),
.Y(n_9889)
);

INVx1_ASAP7_75t_L g9890 ( 
.A(n_8926),
.Y(n_9890)
);

AND2x4_ASAP7_75t_L g9891 ( 
.A(n_9114),
.B(n_353),
.Y(n_9891)
);

NAND2xp5_ASAP7_75t_SL g9892 ( 
.A(n_9101),
.B(n_354),
.Y(n_9892)
);

INVx2_ASAP7_75t_L g9893 ( 
.A(n_9093),
.Y(n_9893)
);

INVx2_ASAP7_75t_L g9894 ( 
.A(n_8709),
.Y(n_9894)
);

BUFx2_ASAP7_75t_L g9895 ( 
.A(n_8754),
.Y(n_9895)
);

INVx1_ASAP7_75t_L g9896 ( 
.A(n_9059),
.Y(n_9896)
);

AND2x2_ASAP7_75t_L g9897 ( 
.A(n_8778),
.B(n_354),
.Y(n_9897)
);

NOR2xp33_ASAP7_75t_R g9898 ( 
.A(n_8715),
.B(n_355),
.Y(n_9898)
);

CKINVDCx5p33_ASAP7_75t_R g9899 ( 
.A(n_8853),
.Y(n_9899)
);

NAND2xp5_ASAP7_75t_L g9900 ( 
.A(n_8713),
.B(n_355),
.Y(n_9900)
);

NAND2xp5_ASAP7_75t_L g9901 ( 
.A(n_8713),
.B(n_356),
.Y(n_9901)
);

AND2x4_ASAP7_75t_L g9902 ( 
.A(n_8864),
.B(n_356),
.Y(n_9902)
);

INVx3_ASAP7_75t_L g9903 ( 
.A(n_8736),
.Y(n_9903)
);

BUFx4f_ASAP7_75t_L g9904 ( 
.A(n_8840),
.Y(n_9904)
);

NAND2xp5_ASAP7_75t_L g9905 ( 
.A(n_8713),
.B(n_357),
.Y(n_9905)
);

NOR2xp67_ASAP7_75t_L g9906 ( 
.A(n_9181),
.B(n_357),
.Y(n_9906)
);

NOR2xp67_ASAP7_75t_L g9907 ( 
.A(n_9181),
.B(n_358),
.Y(n_9907)
);

INVx1_ASAP7_75t_L g9908 ( 
.A(n_9059),
.Y(n_9908)
);

INVx2_ASAP7_75t_SL g9909 ( 
.A(n_8722),
.Y(n_9909)
);

NAND2xp5_ASAP7_75t_L g9910 ( 
.A(n_8713),
.B(n_360),
.Y(n_9910)
);

NOR3xp33_ASAP7_75t_L g9911 ( 
.A(n_8719),
.B(n_360),
.C(n_361),
.Y(n_9911)
);

INVx2_ASAP7_75t_SL g9912 ( 
.A(n_8722),
.Y(n_9912)
);

OR2x2_ASAP7_75t_SL g9913 ( 
.A(n_9017),
.B(n_362),
.Y(n_9913)
);

INVx2_ASAP7_75t_L g9914 ( 
.A(n_8709),
.Y(n_9914)
);

AOI22xp33_ASAP7_75t_L g9915 ( 
.A1(n_9193),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_9915)
);

AO22x1_ASAP7_75t_L g9916 ( 
.A1(n_8984),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_9916)
);

NOR3xp33_ASAP7_75t_SL g9917 ( 
.A(n_8719),
.B(n_365),
.C(n_366),
.Y(n_9917)
);

A2O1A1Ixp33_ASAP7_75t_L g9918 ( 
.A1(n_8719),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_9918)
);

AO22x1_ASAP7_75t_L g9919 ( 
.A1(n_8984),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_9059),
.Y(n_9920)
);

INVx1_ASAP7_75t_L g9921 ( 
.A(n_9059),
.Y(n_9921)
);

INVx2_ASAP7_75t_L g9922 ( 
.A(n_8709),
.Y(n_9922)
);

NOR3xp33_ASAP7_75t_SL g9923 ( 
.A(n_8719),
.B(n_371),
.C(n_372),
.Y(n_9923)
);

BUFx2_ASAP7_75t_L g9924 ( 
.A(n_8754),
.Y(n_9924)
);

INVx1_ASAP7_75t_L g9925 ( 
.A(n_9059),
.Y(n_9925)
);

OAI22xp33_ASAP7_75t_L g9926 ( 
.A1(n_8725),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_9926)
);

INVx2_ASAP7_75t_L g9927 ( 
.A(n_8709),
.Y(n_9927)
);

NAND2xp5_ASAP7_75t_L g9928 ( 
.A(n_8713),
.B(n_373),
.Y(n_9928)
);

BUFx2_ASAP7_75t_L g9929 ( 
.A(n_8754),
.Y(n_9929)
);

OR2x2_ASAP7_75t_L g9930 ( 
.A(n_8953),
.B(n_376),
.Y(n_9930)
);

INVx1_ASAP7_75t_L g9931 ( 
.A(n_9059),
.Y(n_9931)
);

INVx1_ASAP7_75t_L g9932 ( 
.A(n_9059),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_9059),
.Y(n_9933)
);

CKINVDCx5p33_ASAP7_75t_R g9934 ( 
.A(n_8853),
.Y(n_9934)
);

HB1xp67_ASAP7_75t_L g9935 ( 
.A(n_8856),
.Y(n_9935)
);

NAND2xp5_ASAP7_75t_L g9936 ( 
.A(n_8713),
.B(n_376),
.Y(n_9936)
);

NOR2xp33_ASAP7_75t_L g9937 ( 
.A(n_8719),
.B(n_377),
.Y(n_9937)
);

AOI22xp33_ASAP7_75t_L g9938 ( 
.A1(n_9193),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_9938)
);

INVx1_ASAP7_75t_L g9939 ( 
.A(n_9059),
.Y(n_9939)
);

NAND2xp5_ASAP7_75t_L g9940 ( 
.A(n_8713),
.B(n_378),
.Y(n_9940)
);

INVx1_ASAP7_75t_SL g9941 ( 
.A(n_8907),
.Y(n_9941)
);

CKINVDCx5p33_ASAP7_75t_R g9942 ( 
.A(n_8853),
.Y(n_9942)
);

NAND2xp5_ASAP7_75t_L g9943 ( 
.A(n_8713),
.B(n_379),
.Y(n_9943)
);

NAND2xp5_ASAP7_75t_L g9944 ( 
.A(n_8713),
.B(n_380),
.Y(n_9944)
);

AND2x6_ASAP7_75t_SL g9945 ( 
.A(n_8837),
.B(n_381),
.Y(n_9945)
);

OR2x6_ASAP7_75t_L g9946 ( 
.A(n_8865),
.B(n_382),
.Y(n_9946)
);

AND2x2_ASAP7_75t_L g9947 ( 
.A(n_8778),
.B(n_383),
.Y(n_9947)
);

BUFx4f_ASAP7_75t_L g9948 ( 
.A(n_8840),
.Y(n_9948)
);

INVx2_ASAP7_75t_L g9949 ( 
.A(n_8709),
.Y(n_9949)
);

AOI22xp5_ASAP7_75t_L g9950 ( 
.A1(n_9077),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_9950)
);

AND2x2_ASAP7_75t_L g9951 ( 
.A(n_8778),
.B(n_384),
.Y(n_9951)
);

AND2x2_ASAP7_75t_L g9952 ( 
.A(n_8778),
.B(n_385),
.Y(n_9952)
);

INVx2_ASAP7_75t_L g9953 ( 
.A(n_8709),
.Y(n_9953)
);

NAND2xp5_ASAP7_75t_L g9954 ( 
.A(n_8713),
.B(n_386),
.Y(n_9954)
);

AOI22xp5_ASAP7_75t_L g9955 ( 
.A1(n_9077),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_9955)
);

INVx4_ASAP7_75t_L g9956 ( 
.A(n_9245),
.Y(n_9956)
);

INVx1_ASAP7_75t_L g9957 ( 
.A(n_9059),
.Y(n_9957)
);

HB1xp67_ASAP7_75t_L g9958 ( 
.A(n_8856),
.Y(n_9958)
);

INVx1_ASAP7_75t_SL g9959 ( 
.A(n_8907),
.Y(n_9959)
);

BUFx8_ASAP7_75t_L g9960 ( 
.A(n_8840),
.Y(n_9960)
);

BUFx6f_ASAP7_75t_L g9961 ( 
.A(n_8722),
.Y(n_9961)
);

AND2x4_ASAP7_75t_L g9962 ( 
.A(n_8864),
.B(n_388),
.Y(n_9962)
);

BUFx3_ASAP7_75t_L g9963 ( 
.A(n_8716),
.Y(n_9963)
);

O2A1O1Ixp33_ASAP7_75t_L g9964 ( 
.A1(n_8719),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_9964)
);

NAND2xp5_ASAP7_75t_SL g9965 ( 
.A(n_8719),
.B(n_390),
.Y(n_9965)
);

BUFx4f_ASAP7_75t_L g9966 ( 
.A(n_8840),
.Y(n_9966)
);

INVx2_ASAP7_75t_L g9967 ( 
.A(n_8709),
.Y(n_9967)
);

AOI22xp5_ASAP7_75t_L g9968 ( 
.A1(n_9077),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_9968)
);

INVx3_ASAP7_75t_L g9969 ( 
.A(n_8736),
.Y(n_9969)
);

BUFx4f_ASAP7_75t_L g9970 ( 
.A(n_8840),
.Y(n_9970)
);

INVx1_ASAP7_75t_L g9971 ( 
.A(n_9059),
.Y(n_9971)
);

BUFx3_ASAP7_75t_L g9972 ( 
.A(n_8716),
.Y(n_9972)
);

HB1xp67_ASAP7_75t_L g9973 ( 
.A(n_8856),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_9059),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_9059),
.Y(n_9975)
);

NOR2xp33_ASAP7_75t_SL g9976 ( 
.A(n_8853),
.B(n_392),
.Y(n_9976)
);

AOI22xp33_ASAP7_75t_L g9977 ( 
.A1(n_9193),
.A2(n_396),
.B1(n_393),
.B2(n_394),
.Y(n_9977)
);

INVx2_ASAP7_75t_L g9978 ( 
.A(n_8709),
.Y(n_9978)
);

BUFx3_ASAP7_75t_L g9979 ( 
.A(n_8716),
.Y(n_9979)
);

NAND2xp5_ASAP7_75t_L g9980 ( 
.A(n_8713),
.B(n_394),
.Y(n_9980)
);

NAND2xp5_ASAP7_75t_L g9981 ( 
.A(n_8713),
.B(n_397),
.Y(n_9981)
);

HB1xp67_ASAP7_75t_L g9982 ( 
.A(n_8856),
.Y(n_9982)
);

NOR2x1p5_ASAP7_75t_L g9983 ( 
.A(n_9191),
.B(n_398),
.Y(n_9983)
);

BUFx3_ASAP7_75t_L g9984 ( 
.A(n_8716),
.Y(n_9984)
);

CKINVDCx16_ASAP7_75t_R g9985 ( 
.A(n_8840),
.Y(n_9985)
);

AND2x2_ASAP7_75t_L g9986 ( 
.A(n_8778),
.B(n_398),
.Y(n_9986)
);

NAND2xp5_ASAP7_75t_L g9987 ( 
.A(n_8713),
.B(n_399),
.Y(n_9987)
);

NAND2xp5_ASAP7_75t_L g9988 ( 
.A(n_8713),
.B(n_399),
.Y(n_9988)
);

NAND3xp33_ASAP7_75t_SL g9989 ( 
.A(n_8719),
.B(n_400),
.C(n_401),
.Y(n_9989)
);

NOR3xp33_ASAP7_75t_SL g9990 ( 
.A(n_8719),
.B(n_400),
.C(n_402),
.Y(n_9990)
);

INVx1_ASAP7_75t_L g9991 ( 
.A(n_9059),
.Y(n_9991)
);

NAND2xp5_ASAP7_75t_L g9992 ( 
.A(n_9464),
.B(n_402),
.Y(n_9992)
);

AOI21xp5_ASAP7_75t_L g9993 ( 
.A1(n_9641),
.A2(n_403),
.B(n_404),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_9542),
.Y(n_9994)
);

A2O1A1Ixp33_ASAP7_75t_L g9995 ( 
.A1(n_9535),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_9995)
);

INVx3_ASAP7_75t_L g9996 ( 
.A(n_9557),
.Y(n_9996)
);

AOI21xp5_ASAP7_75t_L g9997 ( 
.A1(n_9659),
.A2(n_405),
.B(n_406),
.Y(n_9997)
);

AO21x1_ASAP7_75t_L g9998 ( 
.A1(n_9937),
.A2(n_406),
.B(n_407),
.Y(n_9998)
);

BUFx3_ASAP7_75t_L g9999 ( 
.A(n_9417),
.Y(n_9999)
);

NAND2xp5_ASAP7_75t_L g10000 ( 
.A(n_9325),
.B(n_407),
.Y(n_10000)
);

NAND2xp5_ASAP7_75t_SL g10001 ( 
.A(n_9847),
.B(n_408),
.Y(n_10001)
);

AOI22xp5_ASAP7_75t_L g10002 ( 
.A1(n_9597),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_10002)
);

INVx1_ASAP7_75t_L g10003 ( 
.A(n_9301),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_9320),
.Y(n_10004)
);

NAND3xp33_ASAP7_75t_SL g10005 ( 
.A(n_9911),
.B(n_409),
.C(n_410),
.Y(n_10005)
);

BUFx2_ASAP7_75t_L g10006 ( 
.A(n_9459),
.Y(n_10006)
);

NAND2xp5_ASAP7_75t_L g10007 ( 
.A(n_9532),
.B(n_411),
.Y(n_10007)
);

O2A1O1Ixp33_ASAP7_75t_L g10008 ( 
.A1(n_9778),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_10008)
);

CKINVDCx5p33_ASAP7_75t_R g10009 ( 
.A(n_9303),
.Y(n_10009)
);

AOI22xp5_ASAP7_75t_L g10010 ( 
.A1(n_9559),
.A2(n_415),
.B1(n_412),
.B2(n_414),
.Y(n_10010)
);

CKINVDCx20_ASAP7_75t_R g10011 ( 
.A(n_9606),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_9896),
.Y(n_10012)
);

O2A1O1Ixp33_ASAP7_75t_L g10013 ( 
.A1(n_9312),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_10013)
);

HB1xp67_ASAP7_75t_L g10014 ( 
.A(n_9302),
.Y(n_10014)
);

INVx1_ASAP7_75t_L g10015 ( 
.A(n_9908),
.Y(n_10015)
);

AOI21xp5_ASAP7_75t_L g10016 ( 
.A1(n_9634),
.A2(n_416),
.B(n_417),
.Y(n_10016)
);

O2A1O1Ixp33_ASAP7_75t_L g10017 ( 
.A1(n_9918),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_10017)
);

AND2x2_ASAP7_75t_L g10018 ( 
.A(n_9752),
.B(n_418),
.Y(n_10018)
);

NOR2xp33_ASAP7_75t_L g10019 ( 
.A(n_9773),
.B(n_419),
.Y(n_10019)
);

BUFx4f_ASAP7_75t_L g10020 ( 
.A(n_9336),
.Y(n_10020)
);

O2A1O1Ixp33_ASAP7_75t_L g10021 ( 
.A1(n_9965),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_10021)
);

A2O1A1Ixp33_ASAP7_75t_L g10022 ( 
.A1(n_9964),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_10022)
);

NAND2xp5_ASAP7_75t_SL g10023 ( 
.A(n_9587),
.B(n_423),
.Y(n_10023)
);

OAI21xp33_ASAP7_75t_L g10024 ( 
.A1(n_9917),
.A2(n_424),
.B(n_425),
.Y(n_10024)
);

NOR2xp33_ASAP7_75t_L g10025 ( 
.A(n_9310),
.B(n_425),
.Y(n_10025)
);

AOI21xp5_ASAP7_75t_L g10026 ( 
.A1(n_9503),
.A2(n_426),
.B(n_427),
.Y(n_10026)
);

AOI21xp5_ASAP7_75t_L g10027 ( 
.A1(n_9733),
.A2(n_426),
.B(n_427),
.Y(n_10027)
);

AND2x2_ASAP7_75t_L g10028 ( 
.A(n_9305),
.B(n_428),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_9920),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_9921),
.Y(n_10030)
);

NAND2xp5_ASAP7_75t_L g10031 ( 
.A(n_9536),
.B(n_428),
.Y(n_10031)
);

AOI21x1_ASAP7_75t_L g10032 ( 
.A1(n_9498),
.A2(n_429),
.B(n_430),
.Y(n_10032)
);

A2O1A1Ixp33_ASAP7_75t_L g10033 ( 
.A1(n_9923),
.A2(n_432),
.B(n_429),
.C(n_431),
.Y(n_10033)
);

OAI22xp5_ASAP7_75t_L g10034 ( 
.A1(n_9365),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_9545),
.Y(n_10035)
);

NOR2xp33_ASAP7_75t_R g10036 ( 
.A(n_9388),
.B(n_433),
.Y(n_10036)
);

OAI22xp5_ASAP7_75t_L g10037 ( 
.A1(n_9950),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_10037)
);

BUFx2_ASAP7_75t_L g10038 ( 
.A(n_9334),
.Y(n_10038)
);

NAND3xp33_ASAP7_75t_SL g10039 ( 
.A(n_9768),
.B(n_435),
.C(n_436),
.Y(n_10039)
);

NAND2xp5_ASAP7_75t_L g10040 ( 
.A(n_9772),
.B(n_437),
.Y(n_10040)
);

BUFx2_ASAP7_75t_L g10041 ( 
.A(n_9448),
.Y(n_10041)
);

INVx2_ASAP7_75t_L g10042 ( 
.A(n_9652),
.Y(n_10042)
);

BUFx12f_ASAP7_75t_L g10043 ( 
.A(n_9960),
.Y(n_10043)
);

HB1xp67_ASAP7_75t_L g10044 ( 
.A(n_9935),
.Y(n_10044)
);

NOR2xp33_ASAP7_75t_L g10045 ( 
.A(n_9941),
.B(n_438),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_9925),
.Y(n_10046)
);

AO21x1_ASAP7_75t_L g10047 ( 
.A1(n_9845),
.A2(n_439),
.B(n_440),
.Y(n_10047)
);

AOI21xp5_ASAP7_75t_L g10048 ( 
.A1(n_9821),
.A2(n_9668),
.B(n_9667),
.Y(n_10048)
);

NOR2xp33_ASAP7_75t_L g10049 ( 
.A(n_9959),
.B(n_439),
.Y(n_10049)
);

NOR2xp33_ASAP7_75t_R g10050 ( 
.A(n_9577),
.B(n_441),
.Y(n_10050)
);

INVx1_ASAP7_75t_L g10051 ( 
.A(n_9931),
.Y(n_10051)
);

OR2x6_ASAP7_75t_L g10052 ( 
.A(n_9795),
.B(n_442),
.Y(n_10052)
);

OAI22xp5_ASAP7_75t_L g10053 ( 
.A1(n_9955),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_10053)
);

O2A1O1Ixp33_ASAP7_75t_L g10054 ( 
.A1(n_9561),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_10054)
);

A2O1A1Ixp33_ASAP7_75t_L g10055 ( 
.A1(n_9990),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_SL g10056 ( 
.A(n_9587),
.B(n_449),
.Y(n_10056)
);

NOR3xp33_ASAP7_75t_SL g10057 ( 
.A(n_9813),
.B(n_449),
.C(n_450),
.Y(n_10057)
);

OR2x6_ASAP7_75t_L g10058 ( 
.A(n_9666),
.B(n_450),
.Y(n_10058)
);

NAND2xp5_ASAP7_75t_L g10059 ( 
.A(n_9777),
.B(n_451),
.Y(n_10059)
);

INVx3_ASAP7_75t_L g10060 ( 
.A(n_9307),
.Y(n_10060)
);

NOR2xp33_ASAP7_75t_L g10061 ( 
.A(n_9741),
.B(n_451),
.Y(n_10061)
);

INVx1_ASAP7_75t_L g10062 ( 
.A(n_9932),
.Y(n_10062)
);

BUFx12f_ASAP7_75t_L g10063 ( 
.A(n_9308),
.Y(n_10063)
);

AOI22xp5_ASAP7_75t_L g10064 ( 
.A1(n_9844),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_10064)
);

BUFx24_ASAP7_75t_L g10065 ( 
.A(n_9615),
.Y(n_10065)
);

NAND2xp5_ASAP7_75t_L g10066 ( 
.A(n_9322),
.B(n_453),
.Y(n_10066)
);

NAND3xp33_ASAP7_75t_L g10067 ( 
.A(n_9628),
.B(n_454),
.C(n_455),
.Y(n_10067)
);

AOI21xp5_ASAP7_75t_L g10068 ( 
.A1(n_9560),
.A2(n_9720),
.B(n_9866),
.Y(n_10068)
);

INVx2_ASAP7_75t_L g10069 ( 
.A(n_9572),
.Y(n_10069)
);

AOI21xp5_ASAP7_75t_L g10070 ( 
.A1(n_9851),
.A2(n_455),
.B(n_457),
.Y(n_10070)
);

NOR2xp33_ASAP7_75t_L g10071 ( 
.A(n_9340),
.B(n_457),
.Y(n_10071)
);

BUFx6f_ASAP7_75t_L g10072 ( 
.A(n_9468),
.Y(n_10072)
);

O2A1O1Ixp33_ASAP7_75t_L g10073 ( 
.A1(n_9989),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_10073)
);

INVx1_ASAP7_75t_L g10074 ( 
.A(n_9933),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_9573),
.Y(n_10075)
);

NAND2xp5_ASAP7_75t_SL g10076 ( 
.A(n_9555),
.B(n_458),
.Y(n_10076)
);

INVxp67_ASAP7_75t_SL g10077 ( 
.A(n_9814),
.Y(n_10077)
);

AND2x2_ASAP7_75t_L g10078 ( 
.A(n_9958),
.B(n_459),
.Y(n_10078)
);

AOI21xp5_ASAP7_75t_L g10079 ( 
.A1(n_9719),
.A2(n_460),
.B(n_461),
.Y(n_10079)
);

AOI21x1_ASAP7_75t_L g10080 ( 
.A1(n_9701),
.A2(n_461),
.B(n_462),
.Y(n_10080)
);

AOI22xp33_ASAP7_75t_L g10081 ( 
.A1(n_9888),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_10081)
);

NOR2xp33_ASAP7_75t_L g10082 ( 
.A(n_9756),
.B(n_463),
.Y(n_10082)
);

BUFx6f_ASAP7_75t_L g10083 ( 
.A(n_9417),
.Y(n_10083)
);

NOR2xp33_ASAP7_75t_L g10084 ( 
.A(n_9489),
.B(n_465),
.Y(n_10084)
);

AND2x2_ASAP7_75t_L g10085 ( 
.A(n_9973),
.B(n_465),
.Y(n_10085)
);

CKINVDCx10_ASAP7_75t_R g10086 ( 
.A(n_9985),
.Y(n_10086)
);

OAI22xp5_ASAP7_75t_L g10087 ( 
.A1(n_9968),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9584),
.Y(n_10088)
);

INVx4_ASAP7_75t_L g10089 ( 
.A(n_9419),
.Y(n_10089)
);

NAND2xp5_ASAP7_75t_L g10090 ( 
.A(n_9627),
.B(n_466),
.Y(n_10090)
);

O2A1O1Ixp33_ASAP7_75t_L g10091 ( 
.A1(n_9407),
.A2(n_469),
.B(n_467),
.C(n_468),
.Y(n_10091)
);

OAI21xp33_ASAP7_75t_L g10092 ( 
.A1(n_9515),
.A2(n_470),
.B(n_471),
.Y(n_10092)
);

A2O1A1Ixp33_ASAP7_75t_L g10093 ( 
.A1(n_9368),
.A2(n_472),
.B(n_470),
.C(n_471),
.Y(n_10093)
);

NOR2xp33_ASAP7_75t_L g10094 ( 
.A(n_9510),
.B(n_472),
.Y(n_10094)
);

AOI22xp5_ASAP7_75t_L g10095 ( 
.A1(n_9817),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_10095)
);

INVx6_ASAP7_75t_L g10096 ( 
.A(n_9311),
.Y(n_10096)
);

NAND2xp5_ASAP7_75t_L g10097 ( 
.A(n_9982),
.B(n_473),
.Y(n_10097)
);

A2O1A1Ixp33_ASAP7_75t_L g10098 ( 
.A1(n_9391),
.A2(n_477),
.B(n_475),
.C(n_476),
.Y(n_10098)
);

O2A1O1Ixp33_ASAP7_75t_L g10099 ( 
.A1(n_9824),
.A2(n_479),
.B(n_476),
.C(n_478),
.Y(n_10099)
);

AOI21xp5_ASAP7_75t_L g10100 ( 
.A1(n_9475),
.A2(n_479),
.B(n_480),
.Y(n_10100)
);

NAND2xp5_ASAP7_75t_SL g10101 ( 
.A(n_9555),
.B(n_480),
.Y(n_10101)
);

CKINVDCx20_ASAP7_75t_R g10102 ( 
.A(n_9328),
.Y(n_10102)
);

INVx1_ASAP7_75t_L g10103 ( 
.A(n_9939),
.Y(n_10103)
);

INVx2_ASAP7_75t_L g10104 ( 
.A(n_9585),
.Y(n_10104)
);

NOR2xp33_ASAP7_75t_R g10105 ( 
.A(n_9581),
.B(n_481),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_9592),
.Y(n_10106)
);

AOI21xp5_ASAP7_75t_L g10107 ( 
.A1(n_9441),
.A2(n_481),
.B(n_483),
.Y(n_10107)
);

AO32x1_ASAP7_75t_L g10108 ( 
.A1(n_9780),
.A2(n_485),
.A3(n_483),
.B1(n_484),
.B2(n_486),
.Y(n_10108)
);

A2O1A1Ixp33_ASAP7_75t_L g10109 ( 
.A1(n_9672),
.A2(n_487),
.B(n_484),
.C(n_486),
.Y(n_10109)
);

NOR2xp33_ASAP7_75t_L g10110 ( 
.A(n_9450),
.B(n_487),
.Y(n_10110)
);

O2A1O1Ixp33_ASAP7_75t_SL g10111 ( 
.A1(n_9926),
.A2(n_490),
.B(n_488),
.C(n_489),
.Y(n_10111)
);

INVx2_ASAP7_75t_L g10112 ( 
.A(n_9607),
.Y(n_10112)
);

NAND2xp5_ASAP7_75t_L g10113 ( 
.A(n_9314),
.B(n_489),
.Y(n_10113)
);

INVx1_ASAP7_75t_L g10114 ( 
.A(n_9957),
.Y(n_10114)
);

BUFx6f_ASAP7_75t_L g10115 ( 
.A(n_9422),
.Y(n_10115)
);

NAND2xp5_ASAP7_75t_L g10116 ( 
.A(n_9895),
.B(n_490),
.Y(n_10116)
);

NAND2xp5_ASAP7_75t_L g10117 ( 
.A(n_9924),
.B(n_491),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9971),
.Y(n_10118)
);

AOI21xp5_ASAP7_75t_L g10119 ( 
.A1(n_9666),
.A2(n_491),
.B(n_492),
.Y(n_10119)
);

OAI21xp33_ASAP7_75t_L g10120 ( 
.A1(n_9471),
.A2(n_492),
.B(n_493),
.Y(n_10120)
);

INVx2_ASAP7_75t_L g10121 ( 
.A(n_9609),
.Y(n_10121)
);

HB1xp67_ASAP7_75t_L g10122 ( 
.A(n_9929),
.Y(n_10122)
);

OR2x6_ASAP7_75t_SL g10123 ( 
.A(n_9379),
.B(n_495),
.Y(n_10123)
);

INVx1_ASAP7_75t_L g10124 ( 
.A(n_9974),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_9975),
.Y(n_10125)
);

AOI21xp5_ASAP7_75t_L g10126 ( 
.A1(n_9838),
.A2(n_495),
.B(n_496),
.Y(n_10126)
);

NOR2xp33_ASAP7_75t_L g10127 ( 
.A(n_9766),
.B(n_497),
.Y(n_10127)
);

INVx2_ASAP7_75t_L g10128 ( 
.A(n_9610),
.Y(n_10128)
);

NAND2xp5_ASAP7_75t_L g10129 ( 
.A(n_9802),
.B(n_498),
.Y(n_10129)
);

INVx2_ASAP7_75t_L g10130 ( 
.A(n_9619),
.Y(n_10130)
);

NAND2xp5_ASAP7_75t_L g10131 ( 
.A(n_9779),
.B(n_498),
.Y(n_10131)
);

A2O1A1Ixp33_ASAP7_75t_L g10132 ( 
.A1(n_9731),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_10132)
);

CKINVDCx16_ASAP7_75t_R g10133 ( 
.A(n_9371),
.Y(n_10133)
);

AOI22xp5_ASAP7_75t_L g10134 ( 
.A1(n_9883),
.A2(n_9657),
.B1(n_9882),
.B2(n_9869),
.Y(n_10134)
);

NAND2xp5_ASAP7_75t_SL g10135 ( 
.A(n_9493),
.B(n_500),
.Y(n_10135)
);

NAND2xp5_ASAP7_75t_SL g10136 ( 
.A(n_9493),
.B(n_501),
.Y(n_10136)
);

AOI21xp5_ASAP7_75t_L g10137 ( 
.A1(n_9747),
.A2(n_503),
.B(n_504),
.Y(n_10137)
);

AOI21xp5_ASAP7_75t_L g10138 ( 
.A1(n_9872),
.A2(n_504),
.B(n_505),
.Y(n_10138)
);

INVx1_ASAP7_75t_L g10139 ( 
.A(n_9991),
.Y(n_10139)
);

A2O1A1Ixp33_ASAP7_75t_L g10140 ( 
.A1(n_9580),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_10140)
);

A2O1A1Ixp33_ASAP7_75t_L g10141 ( 
.A1(n_9653),
.A2(n_9859),
.B(n_9529),
.C(n_9697),
.Y(n_10141)
);

NAND2x1p5_ASAP7_75t_L g10142 ( 
.A(n_9807),
.B(n_506),
.Y(n_10142)
);

NAND2xp5_ASAP7_75t_SL g10143 ( 
.A(n_9493),
.B(n_507),
.Y(n_10143)
);

BUFx6f_ASAP7_75t_L g10144 ( 
.A(n_9422),
.Y(n_10144)
);

INVx2_ASAP7_75t_L g10145 ( 
.A(n_9621),
.Y(n_10145)
);

AOI21xp5_ASAP7_75t_L g10146 ( 
.A1(n_9878),
.A2(n_508),
.B(n_509),
.Y(n_10146)
);

NOR2xp33_ASAP7_75t_L g10147 ( 
.A(n_9469),
.B(n_509),
.Y(n_10147)
);

NAND2xp5_ASAP7_75t_SL g10148 ( 
.A(n_9806),
.B(n_510),
.Y(n_10148)
);

INVx1_ASAP7_75t_L g10149 ( 
.A(n_9323),
.Y(n_10149)
);

BUFx3_ASAP7_75t_L g10150 ( 
.A(n_9449),
.Y(n_10150)
);

NAND2xp5_ASAP7_75t_SL g10151 ( 
.A(n_9825),
.B(n_510),
.Y(n_10151)
);

AOI21x1_ASAP7_75t_L g10152 ( 
.A1(n_9840),
.A2(n_511),
.B(n_512),
.Y(n_10152)
);

OAI22xp5_ASAP7_75t_L g10153 ( 
.A1(n_9617),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_10153)
);

A2O1A1Ixp33_ASAP7_75t_L g10154 ( 
.A1(n_9438),
.A2(n_516),
.B(n_513),
.C(n_515),
.Y(n_10154)
);

BUFx2_ASAP7_75t_L g10155 ( 
.A(n_9356),
.Y(n_10155)
);

NOR2xp33_ASAP7_75t_L g10156 ( 
.A(n_9579),
.B(n_515),
.Y(n_10156)
);

A2O1A1Ixp33_ASAP7_75t_L g10157 ( 
.A1(n_9799),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_10157)
);

BUFx2_ASAP7_75t_L g10158 ( 
.A(n_9363),
.Y(n_10158)
);

NOR2xp33_ASAP7_75t_L g10159 ( 
.A(n_9337),
.B(n_517),
.Y(n_10159)
);

BUFx2_ASAP7_75t_L g10160 ( 
.A(n_9685),
.Y(n_10160)
);

AOI21x1_ASAP7_75t_L g10161 ( 
.A1(n_9804),
.A2(n_518),
.B(n_519),
.Y(n_10161)
);

NAND2xp5_ASAP7_75t_SL g10162 ( 
.A(n_9825),
.B(n_520),
.Y(n_10162)
);

HB1xp67_ASAP7_75t_L g10163 ( 
.A(n_9474),
.Y(n_10163)
);

AOI22xp33_ASAP7_75t_L g10164 ( 
.A1(n_9886),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_10164)
);

NAND2xp5_ASAP7_75t_L g10165 ( 
.A(n_9643),
.B(n_521),
.Y(n_10165)
);

AOI21xp5_ASAP7_75t_L g10166 ( 
.A1(n_9636),
.A2(n_522),
.B(n_523),
.Y(n_10166)
);

NOR2xp33_ASAP7_75t_L g10167 ( 
.A(n_9716),
.B(n_524),
.Y(n_10167)
);

NOR2xp33_ASAP7_75t_L g10168 ( 
.A(n_9708),
.B(n_525),
.Y(n_10168)
);

AND2x4_ASAP7_75t_L g10169 ( 
.A(n_9727),
.B(n_525),
.Y(n_10169)
);

AOI21xp5_ASAP7_75t_L g10170 ( 
.A1(n_9642),
.A2(n_526),
.B(n_527),
.Y(n_10170)
);

OAI22xp5_ASAP7_75t_L g10171 ( 
.A1(n_9383),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_10171)
);

CKINVDCx16_ASAP7_75t_R g10172 ( 
.A(n_9496),
.Y(n_10172)
);

INVx2_ASAP7_75t_L g10173 ( 
.A(n_9329),
.Y(n_10173)
);

AOI21xp5_ASAP7_75t_L g10174 ( 
.A1(n_9404),
.A2(n_528),
.B(n_529),
.Y(n_10174)
);

O2A1O1Ixp5_ASAP7_75t_L g10175 ( 
.A1(n_9916),
.A2(n_532),
.B(n_530),
.C(n_531),
.Y(n_10175)
);

BUFx3_ASAP7_75t_L g10176 ( 
.A(n_9449),
.Y(n_10176)
);

BUFx6f_ASAP7_75t_L g10177 ( 
.A(n_9452),
.Y(n_10177)
);

OAI21xp5_ASAP7_75t_L g10178 ( 
.A1(n_9711),
.A2(n_530),
.B(n_532),
.Y(n_10178)
);

AOI21xp5_ASAP7_75t_L g10179 ( 
.A1(n_9404),
.A2(n_533),
.B(n_534),
.Y(n_10179)
);

A2O1A1Ixp33_ASAP7_75t_L g10180 ( 
.A1(n_9544),
.A2(n_536),
.B(n_534),
.C(n_535),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_SL g10181 ( 
.A(n_9848),
.B(n_9871),
.Y(n_10181)
);

NOR2xp33_ASAP7_75t_L g10182 ( 
.A(n_9695),
.B(n_535),
.Y(n_10182)
);

INVx3_ASAP7_75t_L g10183 ( 
.A(n_9307),
.Y(n_10183)
);

HB1xp67_ASAP7_75t_L g10184 ( 
.A(n_9508),
.Y(n_10184)
);

NOR2xp33_ASAP7_75t_L g10185 ( 
.A(n_9457),
.B(n_536),
.Y(n_10185)
);

OAI21x1_ASAP7_75t_L g10186 ( 
.A1(n_9786),
.A2(n_537),
.B(n_538),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_9343),
.Y(n_10187)
);

O2A1O1Ixp33_ASAP7_75t_L g10188 ( 
.A1(n_9506),
.A2(n_540),
.B(n_537),
.C(n_539),
.Y(n_10188)
);

INVx2_ASAP7_75t_L g10189 ( 
.A(n_9346),
.Y(n_10189)
);

NAND2xp5_ASAP7_75t_SL g10190 ( 
.A(n_9848),
.B(n_539),
.Y(n_10190)
);

OAI22xp5_ASAP7_75t_L g10191 ( 
.A1(n_9528),
.A2(n_9881),
.B1(n_9433),
.B2(n_9696),
.Y(n_10191)
);

OAI22xp5_ASAP7_75t_L g10192 ( 
.A1(n_9533),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_10192)
);

OAI22xp5_ASAP7_75t_L g10193 ( 
.A1(n_9874),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_10193)
);

AOI21xp5_ASAP7_75t_L g10194 ( 
.A1(n_9405),
.A2(n_543),
.B(n_544),
.Y(n_10194)
);

AOI22xp33_ASAP7_75t_L g10195 ( 
.A1(n_9886),
.A2(n_546),
.B1(n_544),
.B2(n_545),
.Y(n_10195)
);

INVx2_ASAP7_75t_L g10196 ( 
.A(n_9355),
.Y(n_10196)
);

NAND2xp5_ASAP7_75t_L g10197 ( 
.A(n_9769),
.B(n_545),
.Y(n_10197)
);

OA21x2_ASAP7_75t_L g10198 ( 
.A1(n_9798),
.A2(n_546),
.B(n_547),
.Y(n_10198)
);

INVx1_ASAP7_75t_L g10199 ( 
.A(n_9358),
.Y(n_10199)
);

HB1xp67_ASAP7_75t_L g10200 ( 
.A(n_9605),
.Y(n_10200)
);

NAND2xp5_ASAP7_75t_L g10201 ( 
.A(n_9702),
.B(n_548),
.Y(n_10201)
);

AOI21xp5_ASAP7_75t_L g10202 ( 
.A1(n_9405),
.A2(n_548),
.B(n_549),
.Y(n_10202)
);

OAI22xp5_ASAP7_75t_L g10203 ( 
.A1(n_9946),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_10203)
);

BUFx6f_ASAP7_75t_L g10204 ( 
.A(n_9452),
.Y(n_10204)
);

INVxp67_ASAP7_75t_SL g10205 ( 
.A(n_9631),
.Y(n_10205)
);

A2O1A1Ixp33_ASAP7_75t_L g10206 ( 
.A1(n_9399),
.A2(n_553),
.B(n_550),
.C(n_552),
.Y(n_10206)
);

NAND2xp5_ASAP7_75t_SL g10207 ( 
.A(n_9871),
.B(n_552),
.Y(n_10207)
);

AOI21xp5_ASAP7_75t_L g10208 ( 
.A1(n_9524),
.A2(n_553),
.B(n_554),
.Y(n_10208)
);

OAI22xp5_ASAP7_75t_L g10209 ( 
.A1(n_9946),
.A2(n_9434),
.B1(n_9638),
.B2(n_9734),
.Y(n_10209)
);

INVx3_ASAP7_75t_L g10210 ( 
.A(n_9316),
.Y(n_10210)
);

INVx1_ASAP7_75t_L g10211 ( 
.A(n_9366),
.Y(n_10211)
);

NAND2xp5_ASAP7_75t_SL g10212 ( 
.A(n_9863),
.B(n_554),
.Y(n_10212)
);

INVx2_ASAP7_75t_L g10213 ( 
.A(n_9382),
.Y(n_10213)
);

NOR2xp33_ASAP7_75t_L g10214 ( 
.A(n_9690),
.B(n_9715),
.Y(n_10214)
);

O2A1O1Ixp5_ASAP7_75t_L g10215 ( 
.A1(n_9919),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_10215)
);

O2A1O1Ixp33_ASAP7_75t_SL g10216 ( 
.A1(n_9526),
.A2(n_558),
.B(n_555),
.C(n_556),
.Y(n_10216)
);

NAND2xp5_ASAP7_75t_L g10217 ( 
.A(n_9319),
.B(n_559),
.Y(n_10217)
);

INVx1_ASAP7_75t_L g10218 ( 
.A(n_9385),
.Y(n_10218)
);

NAND2xp5_ASAP7_75t_L g10219 ( 
.A(n_9793),
.B(n_559),
.Y(n_10219)
);

AOI21xp5_ASAP7_75t_L g10220 ( 
.A1(n_9524),
.A2(n_561),
.B(n_562),
.Y(n_10220)
);

INVx1_ASAP7_75t_SL g10221 ( 
.A(n_9416),
.Y(n_10221)
);

NAND2xp5_ASAP7_75t_L g10222 ( 
.A(n_9750),
.B(n_561),
.Y(n_10222)
);

INVx1_ASAP7_75t_SL g10223 ( 
.A(n_9461),
.Y(n_10223)
);

OAI22xp5_ASAP7_75t_L g10224 ( 
.A1(n_9738),
.A2(n_565),
.B1(n_562),
.B2(n_563),
.Y(n_10224)
);

BUFx8_ASAP7_75t_L g10225 ( 
.A(n_9546),
.Y(n_10225)
);

NAND2xp5_ASAP7_75t_L g10226 ( 
.A(n_9751),
.B(n_563),
.Y(n_10226)
);

INVx1_ASAP7_75t_L g10227 ( 
.A(n_9394),
.Y(n_10227)
);

OR2x6_ASAP7_75t_L g10228 ( 
.A(n_9616),
.B(n_565),
.Y(n_10228)
);

INVx2_ASAP7_75t_SL g10229 ( 
.A(n_9473),
.Y(n_10229)
);

NAND3xp33_ASAP7_75t_L g10230 ( 
.A(n_9551),
.B(n_566),
.C(n_567),
.Y(n_10230)
);

OAI22xp5_ASAP7_75t_L g10231 ( 
.A1(n_9776),
.A2(n_569),
.B1(n_566),
.B2(n_568),
.Y(n_10231)
);

INVx1_ASAP7_75t_L g10232 ( 
.A(n_9395),
.Y(n_10232)
);

AOI22xp5_ASAP7_75t_L g10233 ( 
.A1(n_9873),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.Y(n_10233)
);

AOI21xp5_ASAP7_75t_L g10234 ( 
.A1(n_9556),
.A2(n_571),
.B(n_572),
.Y(n_10234)
);

INVx1_ASAP7_75t_L g10235 ( 
.A(n_9398),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9400),
.Y(n_10236)
);

O2A1O1Ixp33_ASAP7_75t_L g10237 ( 
.A1(n_9608),
.A2(n_9674),
.B(n_9692),
.C(n_9849),
.Y(n_10237)
);

INVx2_ASAP7_75t_L g10238 ( 
.A(n_9406),
.Y(n_10238)
);

INVx1_ASAP7_75t_L g10239 ( 
.A(n_9411),
.Y(n_10239)
);

BUFx6f_ASAP7_75t_L g10240 ( 
.A(n_9473),
.Y(n_10240)
);

NAND2xp5_ASAP7_75t_L g10241 ( 
.A(n_9758),
.B(n_571),
.Y(n_10241)
);

INVx2_ASAP7_75t_L g10242 ( 
.A(n_9414),
.Y(n_10242)
);

NOR2xp67_ASAP7_75t_L g10243 ( 
.A(n_9333),
.B(n_573),
.Y(n_10243)
);

NAND2xp33_ASAP7_75t_R g10244 ( 
.A(n_9423),
.B(n_573),
.Y(n_10244)
);

NOR2xp33_ASAP7_75t_L g10245 ( 
.A(n_9324),
.B(n_574),
.Y(n_10245)
);

NAND2xp5_ASAP7_75t_L g10246 ( 
.A(n_9837),
.B(n_575),
.Y(n_10246)
);

CKINVDCx5p33_ASAP7_75t_R g10247 ( 
.A(n_9899),
.Y(n_10247)
);

HB1xp67_ASAP7_75t_L g10248 ( 
.A(n_9420),
.Y(n_10248)
);

OAI22xp5_ASAP7_75t_L g10249 ( 
.A1(n_9454),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_10249)
);

OAI22xp5_ASAP7_75t_L g10250 ( 
.A1(n_9732),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_10250)
);

AOI22xp5_ASAP7_75t_L g10251 ( 
.A1(n_9873),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_10251)
);

BUFx12f_ASAP7_75t_L g10252 ( 
.A(n_9357),
.Y(n_10252)
);

BUFx6f_ASAP7_75t_L g10253 ( 
.A(n_9478),
.Y(n_10253)
);

AOI21xp5_ASAP7_75t_L g10254 ( 
.A1(n_9556),
.A2(n_579),
.B(n_580),
.Y(n_10254)
);

AOI21xp5_ASAP7_75t_L g10255 ( 
.A1(n_9483),
.A2(n_581),
.B(n_582),
.Y(n_10255)
);

AOI21xp5_ASAP7_75t_L g10256 ( 
.A1(n_9616),
.A2(n_582),
.B(n_583),
.Y(n_10256)
);

AOI21xp5_ASAP7_75t_L g10257 ( 
.A1(n_9645),
.A2(n_583),
.B(n_585),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_9425),
.Y(n_10258)
);

BUFx6f_ASAP7_75t_SL g10259 ( 
.A(n_9902),
.Y(n_10259)
);

INVx4_ASAP7_75t_L g10260 ( 
.A(n_9419),
.Y(n_10260)
);

OAI21xp5_ASAP7_75t_L g10261 ( 
.A1(n_9836),
.A2(n_587),
.B(n_588),
.Y(n_10261)
);

AO21x2_ASAP7_75t_L g10262 ( 
.A1(n_9675),
.A2(n_587),
.B(n_588),
.Y(n_10262)
);

OAI21xp5_ASAP7_75t_L g10263 ( 
.A1(n_9889),
.A2(n_9601),
.B(n_9864),
.Y(n_10263)
);

NOR2xp67_ASAP7_75t_L g10264 ( 
.A(n_9351),
.B(n_589),
.Y(n_10264)
);

OAI21x1_ASAP7_75t_L g10265 ( 
.A1(n_9677),
.A2(n_590),
.B(n_591),
.Y(n_10265)
);

AND2x2_ASAP7_75t_L g10266 ( 
.A(n_9812),
.B(n_592),
.Y(n_10266)
);

BUFx6f_ASAP7_75t_L g10267 ( 
.A(n_9478),
.Y(n_10267)
);

BUFx6f_ASAP7_75t_L g10268 ( 
.A(n_9316),
.Y(n_10268)
);

AOI21xp5_ASAP7_75t_L g10269 ( 
.A1(n_9645),
.A2(n_592),
.B(n_593),
.Y(n_10269)
);

INVx2_ASAP7_75t_L g10270 ( 
.A(n_9436),
.Y(n_10270)
);

INVx2_ASAP7_75t_L g10271 ( 
.A(n_9437),
.Y(n_10271)
);

AND2x4_ASAP7_75t_L g10272 ( 
.A(n_9456),
.B(n_594),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9440),
.Y(n_10273)
);

NAND2xp5_ASAP7_75t_L g10274 ( 
.A(n_9339),
.B(n_595),
.Y(n_10274)
);

BUFx3_ASAP7_75t_L g10275 ( 
.A(n_9963),
.Y(n_10275)
);

AND2x4_ASAP7_75t_L g10276 ( 
.A(n_9362),
.B(n_595),
.Y(n_10276)
);

CKINVDCx6p67_ASAP7_75t_R g10277 ( 
.A(n_9311),
.Y(n_10277)
);

AOI21xp5_ASAP7_75t_L g10278 ( 
.A1(n_9892),
.A2(n_596),
.B(n_597),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_9442),
.Y(n_10279)
);

NAND2xp5_ASAP7_75t_L g10280 ( 
.A(n_9451),
.B(n_596),
.Y(n_10280)
);

HB1xp67_ASAP7_75t_L g10281 ( 
.A(n_9455),
.Y(n_10281)
);

INVx2_ASAP7_75t_L g10282 ( 
.A(n_9465),
.Y(n_10282)
);

A2O1A1Ixp33_ASAP7_75t_L g10283 ( 
.A1(n_9671),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_10283)
);

NAND2xp5_ASAP7_75t_L g10284 ( 
.A(n_9796),
.B(n_598),
.Y(n_10284)
);

CKINVDCx5p33_ASAP7_75t_R g10285 ( 
.A(n_9934),
.Y(n_10285)
);

CKINVDCx14_ASAP7_75t_R g10286 ( 
.A(n_9898),
.Y(n_10286)
);

OAI22xp5_ASAP7_75t_L g10287 ( 
.A1(n_9870),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_10287)
);

AO22x1_ASAP7_75t_L g10288 ( 
.A1(n_9868),
.A2(n_9629),
.B1(n_9403),
.B2(n_9805),
.Y(n_10288)
);

INVx1_ASAP7_75t_L g10289 ( 
.A(n_9480),
.Y(n_10289)
);

AOI21xp5_ASAP7_75t_L g10290 ( 
.A1(n_9596),
.A2(n_601),
.B(n_602),
.Y(n_10290)
);

AND2x2_ASAP7_75t_L g10291 ( 
.A(n_9745),
.B(n_603),
.Y(n_10291)
);

NOR2xp33_ASAP7_75t_L g10292 ( 
.A(n_9827),
.B(n_604),
.Y(n_10292)
);

O2A1O1Ixp33_ASAP7_75t_L g10293 ( 
.A1(n_9884),
.A2(n_606),
.B(n_604),
.C(n_605),
.Y(n_10293)
);

NAND2xp5_ASAP7_75t_L g10294 ( 
.A(n_9808),
.B(n_605),
.Y(n_10294)
);

INVx1_ASAP7_75t_L g10295 ( 
.A(n_9482),
.Y(n_10295)
);

NAND2xp5_ASAP7_75t_L g10296 ( 
.A(n_9815),
.B(n_607),
.Y(n_10296)
);

INVx3_ASAP7_75t_L g10297 ( 
.A(n_9373),
.Y(n_10297)
);

NOR2x1_ASAP7_75t_R g10298 ( 
.A(n_9761),
.B(n_607),
.Y(n_10298)
);

INVx1_ASAP7_75t_L g10299 ( 
.A(n_9484),
.Y(n_10299)
);

BUFx12f_ASAP7_75t_L g10300 ( 
.A(n_9396),
.Y(n_10300)
);

INVx1_ASAP7_75t_L g10301 ( 
.A(n_9485),
.Y(n_10301)
);

INVx2_ASAP7_75t_L g10302 ( 
.A(n_9488),
.Y(n_10302)
);

A2O1A1Ixp33_ASAP7_75t_L g10303 ( 
.A1(n_9361),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_10303)
);

OAI21xp5_ASAP7_75t_L g10304 ( 
.A1(n_9834),
.A2(n_9681),
.B(n_9832),
.Y(n_10304)
);

NOR2xp33_ASAP7_75t_L g10305 ( 
.A(n_9839),
.B(n_9639),
.Y(n_10305)
);

O2A1O1Ixp5_ASAP7_75t_L g10306 ( 
.A1(n_9700),
.A2(n_611),
.B(n_608),
.C(n_610),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_9490),
.Y(n_10307)
);

OAI22xp5_ASAP7_75t_L g10308 ( 
.A1(n_9913),
.A2(n_9879),
.B1(n_9678),
.B2(n_9315),
.Y(n_10308)
);

NOR2xp33_ASAP7_75t_L g10309 ( 
.A(n_9640),
.B(n_611),
.Y(n_10309)
);

OAI22xp5_ASAP7_75t_L g10310 ( 
.A1(n_9879),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_10310)
);

NOR2xp33_ASAP7_75t_SL g10311 ( 
.A(n_9309),
.B(n_612),
.Y(n_10311)
);

NOR2xp33_ASAP7_75t_L g10312 ( 
.A(n_9781),
.B(n_9788),
.Y(n_10312)
);

INVxp67_ASAP7_75t_L g10313 ( 
.A(n_9374),
.Y(n_10313)
);

A2O1A1Ixp33_ASAP7_75t_L g10314 ( 
.A1(n_9445),
.A2(n_615),
.B(n_613),
.C(n_614),
.Y(n_10314)
);

AOI21xp5_ASAP7_75t_L g10315 ( 
.A1(n_9582),
.A2(n_615),
.B(n_616),
.Y(n_10315)
);

INVxp67_ASAP7_75t_L g10316 ( 
.A(n_9614),
.Y(n_10316)
);

NOR2xp33_ASAP7_75t_R g10317 ( 
.A(n_9942),
.B(n_617),
.Y(n_10317)
);

BUFx12f_ASAP7_75t_L g10318 ( 
.A(n_9603),
.Y(n_10318)
);

AOI22x1_ASAP7_75t_L g10319 ( 
.A1(n_9983),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.Y(n_10319)
);

O2A1O1Ixp5_ASAP7_75t_SL g10320 ( 
.A1(n_9865),
.A2(n_620),
.B(n_618),
.C(n_619),
.Y(n_10320)
);

A2O1A1Ixp33_ASAP7_75t_L g10321 ( 
.A1(n_9828),
.A2(n_622),
.B(n_620),
.C(n_621),
.Y(n_10321)
);

O2A1O1Ixp33_ASAP7_75t_L g10322 ( 
.A1(n_9877),
.A2(n_624),
.B(n_621),
.C(n_623),
.Y(n_10322)
);

NAND2xp5_ASAP7_75t_L g10323 ( 
.A(n_9829),
.B(n_623),
.Y(n_10323)
);

CKINVDCx5p33_ASAP7_75t_R g10324 ( 
.A(n_9569),
.Y(n_10324)
);

AOI21xp5_ASAP7_75t_L g10325 ( 
.A1(n_9791),
.A2(n_624),
.B(n_625),
.Y(n_10325)
);

A2O1A1Ixp33_ASAP7_75t_L g10326 ( 
.A1(n_9885),
.A2(n_628),
.B(n_626),
.C(n_627),
.Y(n_10326)
);

NAND2xp5_ASAP7_75t_L g10327 ( 
.A(n_9833),
.B(n_9842),
.Y(n_10327)
);

AND2x2_ASAP7_75t_L g10328 ( 
.A(n_9753),
.B(n_626),
.Y(n_10328)
);

AOI21xp5_ASAP7_75t_L g10329 ( 
.A1(n_9537),
.A2(n_627),
.B(n_628),
.Y(n_10329)
);

OAI22xp33_ASAP7_75t_L g10330 ( 
.A1(n_9976),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_10330)
);

NAND2xp5_ASAP7_75t_L g10331 ( 
.A(n_9543),
.B(n_630),
.Y(n_10331)
);

AOI21xp5_ASAP7_75t_L g10332 ( 
.A1(n_9547),
.A2(n_9876),
.B(n_9512),
.Y(n_10332)
);

NOR2xp33_ASAP7_75t_R g10333 ( 
.A(n_9904),
.B(n_631),
.Y(n_10333)
);

INVxp67_ASAP7_75t_SL g10334 ( 
.A(n_9552),
.Y(n_10334)
);

O2A1O1Ixp33_ASAP7_75t_L g10335 ( 
.A1(n_9782),
.A2(n_634),
.B(n_632),
.C(n_633),
.Y(n_10335)
);

CKINVDCx5p33_ASAP7_75t_R g10336 ( 
.A(n_9562),
.Y(n_10336)
);

INVx1_ASAP7_75t_L g10337 ( 
.A(n_9492),
.Y(n_10337)
);

NAND2xp5_ASAP7_75t_L g10338 ( 
.A(n_9852),
.B(n_632),
.Y(n_10338)
);

BUFx2_ASAP7_75t_L g10339 ( 
.A(n_9530),
.Y(n_10339)
);

AOI21xp5_ASAP7_75t_L g10340 ( 
.A1(n_9501),
.A2(n_633),
.B(n_634),
.Y(n_10340)
);

A2O1A1Ixp33_ASAP7_75t_SL g10341 ( 
.A1(n_9586),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_10341)
);

NAND2xp5_ASAP7_75t_L g10342 ( 
.A(n_9801),
.B(n_635),
.Y(n_10342)
);

BUFx2_ASAP7_75t_L g10343 ( 
.A(n_9746),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_9505),
.Y(n_10344)
);

INVx1_ASAP7_75t_L g10345 ( 
.A(n_9507),
.Y(n_10345)
);

OR2x2_ASAP7_75t_L g10346 ( 
.A(n_9816),
.B(n_636),
.Y(n_10346)
);

NOR2xp33_ASAP7_75t_L g10347 ( 
.A(n_9789),
.B(n_637),
.Y(n_10347)
);

INVx1_ASAP7_75t_L g10348 ( 
.A(n_9514),
.Y(n_10348)
);

NAND2xp5_ASAP7_75t_SL g10349 ( 
.A(n_9863),
.B(n_638),
.Y(n_10349)
);

OAI22xp5_ASAP7_75t_L g10350 ( 
.A1(n_9678),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_10350)
);

INVx2_ASAP7_75t_L g10351 ( 
.A(n_9520),
.Y(n_10351)
);

NAND3xp33_ASAP7_75t_SL g10352 ( 
.A(n_9694),
.B(n_639),
.C(n_640),
.Y(n_10352)
);

BUFx6f_ASAP7_75t_L g10353 ( 
.A(n_9373),
.Y(n_10353)
);

INVx1_ASAP7_75t_L g10354 ( 
.A(n_9525),
.Y(n_10354)
);

AOI21xp5_ASAP7_75t_L g10355 ( 
.A1(n_9491),
.A2(n_641),
.B(n_642),
.Y(n_10355)
);

INVx2_ASAP7_75t_L g10356 ( 
.A(n_9531),
.Y(n_10356)
);

CKINVDCx5p33_ASAP7_75t_R g10357 ( 
.A(n_9376),
.Y(n_10357)
);

AOI21xp5_ASAP7_75t_L g10358 ( 
.A1(n_9495),
.A2(n_641),
.B(n_642),
.Y(n_10358)
);

NAND2x1p5_ASAP7_75t_L g10359 ( 
.A(n_9564),
.B(n_643),
.Y(n_10359)
);

O2A1O1Ixp33_ASAP7_75t_L g10360 ( 
.A1(n_9688),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_10360)
);

AOI21xp5_ASAP7_75t_L g10361 ( 
.A1(n_9757),
.A2(n_644),
.B(n_645),
.Y(n_10361)
);

NAND2xp5_ASAP7_75t_L g10362 ( 
.A(n_9809),
.B(n_646),
.Y(n_10362)
);

AND2x2_ASAP7_75t_L g10363 ( 
.A(n_9534),
.B(n_646),
.Y(n_10363)
);

INVx1_ASAP7_75t_L g10364 ( 
.A(n_9540),
.Y(n_10364)
);

INVx2_ASAP7_75t_SL g10365 ( 
.A(n_9517),
.Y(n_10365)
);

O2A1O1Ixp33_ASAP7_75t_L g10366 ( 
.A1(n_9754),
.A2(n_649),
.B(n_647),
.C(n_648),
.Y(n_10366)
);

NAND2xp5_ASAP7_75t_L g10367 ( 
.A(n_9820),
.B(n_647),
.Y(n_10367)
);

BUFx3_ASAP7_75t_L g10368 ( 
.A(n_9972),
.Y(n_10368)
);

AOI21xp5_ASAP7_75t_L g10369 ( 
.A1(n_9770),
.A2(n_648),
.B(n_649),
.Y(n_10369)
);

NOR2xp33_ASAP7_75t_L g10370 ( 
.A(n_9611),
.B(n_650),
.Y(n_10370)
);

HB1xp67_ASAP7_75t_L g10371 ( 
.A(n_9775),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9654),
.Y(n_10372)
);

INVx2_ASAP7_75t_SL g10373 ( 
.A(n_9517),
.Y(n_10373)
);

O2A1O1Ixp33_ASAP7_75t_L g10374 ( 
.A1(n_9797),
.A2(n_652),
.B(n_650),
.C(n_651),
.Y(n_10374)
);

NOR3xp33_ASAP7_75t_SL g10375 ( 
.A(n_9463),
.B(n_651),
.C(n_653),
.Y(n_10375)
);

A2O1A1Ixp33_ASAP7_75t_L g10376 ( 
.A1(n_9891),
.A2(n_655),
.B(n_653),
.C(n_654),
.Y(n_10376)
);

AND2x2_ASAP7_75t_L g10377 ( 
.A(n_9725),
.B(n_654),
.Y(n_10377)
);

INVx2_ASAP7_75t_L g10378 ( 
.A(n_9656),
.Y(n_10378)
);

NOR3xp33_ASAP7_75t_SL g10379 ( 
.A(n_9401),
.B(n_655),
.C(n_657),
.Y(n_10379)
);

AOI21xp5_ASAP7_75t_L g10380 ( 
.A1(n_9682),
.A2(n_9822),
.B(n_9890),
.Y(n_10380)
);

INVx2_ASAP7_75t_L g10381 ( 
.A(n_9661),
.Y(n_10381)
);

NAND2xp5_ASAP7_75t_L g10382 ( 
.A(n_9714),
.B(n_657),
.Y(n_10382)
);

OAI21xp33_ASAP7_75t_L g10383 ( 
.A1(n_9915),
.A2(n_658),
.B(n_659),
.Y(n_10383)
);

AOI21xp5_ASAP7_75t_L g10384 ( 
.A1(n_9893),
.A2(n_658),
.B(n_659),
.Y(n_10384)
);

INVx1_ASAP7_75t_L g10385 ( 
.A(n_9665),
.Y(n_10385)
);

HB1xp67_ASAP7_75t_L g10386 ( 
.A(n_9730),
.Y(n_10386)
);

NAND2xp5_ASAP7_75t_L g10387 ( 
.A(n_9819),
.B(n_660),
.Y(n_10387)
);

INVx3_ASAP7_75t_L g10388 ( 
.A(n_9408),
.Y(n_10388)
);

NAND2xp5_ASAP7_75t_L g10389 ( 
.A(n_9726),
.B(n_660),
.Y(n_10389)
);

NAND2xp5_ASAP7_75t_L g10390 ( 
.A(n_9686),
.B(n_661),
.Y(n_10390)
);

OAI21xp5_ASAP7_75t_L g10391 ( 
.A1(n_9938),
.A2(n_661),
.B(n_662),
.Y(n_10391)
);

NOR2x1_ASAP7_75t_SL g10392 ( 
.A(n_9783),
.B(n_662),
.Y(n_10392)
);

AOI22xp33_ASAP7_75t_L g10393 ( 
.A1(n_9403),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_10393)
);

AOI21xp5_ASAP7_75t_L g10394 ( 
.A1(n_9669),
.A2(n_9856),
.B(n_9318),
.Y(n_10394)
);

NAND2xp5_ASAP7_75t_L g10395 ( 
.A(n_9687),
.B(n_663),
.Y(n_10395)
);

OR2x6_ASAP7_75t_L g10396 ( 
.A(n_9709),
.B(n_664),
.Y(n_10396)
);

INVx2_ASAP7_75t_SL g10397 ( 
.A(n_9519),
.Y(n_10397)
);

NAND2xp5_ASAP7_75t_L g10398 ( 
.A(n_9698),
.B(n_666),
.Y(n_10398)
);

INVx1_ASAP7_75t_L g10399 ( 
.A(n_9699),
.Y(n_10399)
);

AOI22xp33_ASAP7_75t_L g10400 ( 
.A1(n_9403),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_10400)
);

CKINVDCx5p33_ASAP7_75t_R g10401 ( 
.A(n_9566),
.Y(n_10401)
);

INVx2_ASAP7_75t_L g10402 ( 
.A(n_9344),
.Y(n_10402)
);

NAND2xp5_ASAP7_75t_SL g10403 ( 
.A(n_9857),
.B(n_667),
.Y(n_10403)
);

A2O1A1Ixp33_ASAP7_75t_L g10404 ( 
.A1(n_9880),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_10404)
);

OR2x6_ASAP7_75t_L g10405 ( 
.A(n_9831),
.B(n_9707),
.Y(n_10405)
);

BUFx6f_ASAP7_75t_L g10406 ( 
.A(n_9408),
.Y(n_10406)
);

O2A1O1Ixp33_ASAP7_75t_L g10407 ( 
.A1(n_9332),
.A2(n_9787),
.B(n_9811),
.C(n_9810),
.Y(n_10407)
);

AOI21xp5_ASAP7_75t_L g10408 ( 
.A1(n_9784),
.A2(n_669),
.B(n_670),
.Y(n_10408)
);

NAND2xp5_ASAP7_75t_L g10409 ( 
.A(n_9706),
.B(n_671),
.Y(n_10409)
);

INVx1_ASAP7_75t_L g10410 ( 
.A(n_9722),
.Y(n_10410)
);

AOI22xp33_ASAP7_75t_L g10411 ( 
.A1(n_9887),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_10411)
);

OR2x6_ASAP7_75t_L g10412 ( 
.A(n_9553),
.B(n_672),
.Y(n_10412)
);

AND2x4_ASAP7_75t_L g10413 ( 
.A(n_9527),
.B(n_673),
.Y(n_10413)
);

NAND2xp5_ASAP7_75t_L g10414 ( 
.A(n_9742),
.B(n_674),
.Y(n_10414)
);

BUFx2_ASAP7_75t_L g10415 ( 
.A(n_9516),
.Y(n_10415)
);

AND2x2_ASAP7_75t_L g10416 ( 
.A(n_9785),
.B(n_675),
.Y(n_10416)
);

AOI22xp33_ASAP7_75t_L g10417 ( 
.A1(n_9875),
.A2(n_678),
.B1(n_675),
.B2(n_677),
.Y(n_10417)
);

AND2x4_ASAP7_75t_L g10418 ( 
.A(n_9472),
.B(n_677),
.Y(n_10418)
);

O2A1O1Ixp33_ASAP7_75t_SL g10419 ( 
.A1(n_9749),
.A2(n_680),
.B(n_678),
.C(n_679),
.Y(n_10419)
);

AND2x4_ASAP7_75t_L g10420 ( 
.A(n_9494),
.B(n_680),
.Y(n_10420)
);

NAND2x1p5_ASAP7_75t_L g10421 ( 
.A(n_9574),
.B(n_681),
.Y(n_10421)
);

INVx1_ASAP7_75t_L g10422 ( 
.A(n_9765),
.Y(n_10422)
);

INVxp67_ASAP7_75t_L g10423 ( 
.A(n_9578),
.Y(n_10423)
);

O2A1O1Ixp33_ASAP7_75t_L g10424 ( 
.A1(n_9823),
.A2(n_683),
.B(n_681),
.C(n_682),
.Y(n_10424)
);

O2A1O1Ixp33_ASAP7_75t_L g10425 ( 
.A1(n_9735),
.A2(n_685),
.B(n_683),
.C(n_684),
.Y(n_10425)
);

NAND2xp5_ASAP7_75t_L g10426 ( 
.A(n_9347),
.B(n_9367),
.Y(n_10426)
);

NAND2xp5_ASAP7_75t_SL g10427 ( 
.A(n_9857),
.B(n_684),
.Y(n_10427)
);

O2A1O1Ixp5_ASAP7_75t_L g10428 ( 
.A1(n_9867),
.A2(n_688),
.B(n_685),
.C(n_686),
.Y(n_10428)
);

OAI22xp5_ASAP7_75t_L g10429 ( 
.A1(n_9977),
.A2(n_689),
.B1(n_686),
.B2(n_688),
.Y(n_10429)
);

INVx3_ASAP7_75t_L g10430 ( 
.A(n_9961),
.Y(n_10430)
);

BUFx6f_ASAP7_75t_L g10431 ( 
.A(n_9961),
.Y(n_10431)
);

BUFx2_ASAP7_75t_L g10432 ( 
.A(n_9748),
.Y(n_10432)
);

NAND2xp5_ASAP7_75t_L g10433 ( 
.A(n_9369),
.B(n_689),
.Y(n_10433)
);

OAI22xp5_ASAP7_75t_L g10434 ( 
.A1(n_9854),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.Y(n_10434)
);

BUFx2_ASAP7_75t_L g10435 ( 
.A(n_9583),
.Y(n_10435)
);

AND2x6_ASAP7_75t_L g10436 ( 
.A(n_9744),
.B(n_690),
.Y(n_10436)
);

INVx2_ASAP7_75t_L g10437 ( 
.A(n_9372),
.Y(n_10437)
);

HB1xp67_ASAP7_75t_L g10438 ( 
.A(n_9755),
.Y(n_10438)
);

AND2x2_ASAP7_75t_L g10439 ( 
.A(n_9549),
.B(n_691),
.Y(n_10439)
);

NOR2xp33_ASAP7_75t_L g10440 ( 
.A(n_9623),
.B(n_693),
.Y(n_10440)
);

BUFx2_ASAP7_75t_L g10441 ( 
.A(n_9342),
.Y(n_10441)
);

NAND2xp5_ASAP7_75t_SL g10442 ( 
.A(n_9759),
.B(n_694),
.Y(n_10442)
);

AND2x2_ASAP7_75t_L g10443 ( 
.A(n_9897),
.B(n_694),
.Y(n_10443)
);

INVx1_ASAP7_75t_L g10444 ( 
.A(n_9377),
.Y(n_10444)
);

INVx1_ASAP7_75t_L g10445 ( 
.A(n_9392),
.Y(n_10445)
);

INVx1_ASAP7_75t_L g10446 ( 
.A(n_9393),
.Y(n_10446)
);

INVx1_ASAP7_75t_L g10447 ( 
.A(n_9397),
.Y(n_10447)
);

NAND2xp5_ASAP7_75t_L g10448 ( 
.A(n_9402),
.B(n_695),
.Y(n_10448)
);

AO32x1_ASAP7_75t_L g10449 ( 
.A1(n_9830),
.A2(n_697),
.A3(n_695),
.B1(n_696),
.B2(n_698),
.Y(n_10449)
);

INVx1_ASAP7_75t_L g10450 ( 
.A(n_9415),
.Y(n_10450)
);

INVx1_ASAP7_75t_L g10451 ( 
.A(n_9421),
.Y(n_10451)
);

NOR2xp33_ASAP7_75t_L g10452 ( 
.A(n_9623),
.B(n_696),
.Y(n_10452)
);

BUFx3_ASAP7_75t_L g10453 ( 
.A(n_9979),
.Y(n_10453)
);

OAI22xp5_ASAP7_75t_L g10454 ( 
.A1(n_9860),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.Y(n_10454)
);

NOR2xp67_ASAP7_75t_L g10455 ( 
.A(n_9956),
.B(n_699),
.Y(n_10455)
);

NAND2xp5_ASAP7_75t_SL g10456 ( 
.A(n_9759),
.B(n_9774),
.Y(n_10456)
);

BUFx2_ASAP7_75t_L g10457 ( 
.A(n_9522),
.Y(n_10457)
);

NAND3xp33_ASAP7_75t_SL g10458 ( 
.A(n_9861),
.B(n_700),
.C(n_701),
.Y(n_10458)
);

AOI21xp5_ASAP7_75t_L g10459 ( 
.A1(n_9792),
.A2(n_702),
.B(n_703),
.Y(n_10459)
);

BUFx6f_ASAP7_75t_L g10460 ( 
.A(n_9519),
.Y(n_10460)
);

NOR2xp33_ASAP7_75t_L g10461 ( 
.A(n_9625),
.B(n_703),
.Y(n_10461)
);

HB1xp67_ASAP7_75t_L g10462 ( 
.A(n_9764),
.Y(n_10462)
);

NAND2xp5_ASAP7_75t_L g10463 ( 
.A(n_9428),
.B(n_704),
.Y(n_10463)
);

BUFx3_ASAP7_75t_L g10464 ( 
.A(n_9984),
.Y(n_10464)
);

NOR2xp33_ASAP7_75t_R g10465 ( 
.A(n_9948),
.B(n_704),
.Y(n_10465)
);

BUFx6f_ASAP7_75t_L g10466 ( 
.A(n_9444),
.Y(n_10466)
);

AOI21xp5_ASAP7_75t_L g10467 ( 
.A1(n_9717),
.A2(n_705),
.B(n_706),
.Y(n_10467)
);

AND2x2_ASAP7_75t_L g10468 ( 
.A(n_9947),
.B(n_705),
.Y(n_10468)
);

BUFx3_ASAP7_75t_L g10469 ( 
.A(n_9509),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_9430),
.B(n_706),
.Y(n_10470)
);

BUFx6f_ASAP7_75t_L g10471 ( 
.A(n_9635),
.Y(n_10471)
);

INVx2_ASAP7_75t_L g10472 ( 
.A(n_9443),
.Y(n_10472)
);

INVxp67_ASAP7_75t_SL g10473 ( 
.A(n_9767),
.Y(n_10473)
);

NAND2xp5_ASAP7_75t_L g10474 ( 
.A(n_9447),
.B(n_707),
.Y(n_10474)
);

OAI21xp33_ASAP7_75t_SL g10475 ( 
.A1(n_9327),
.A2(n_707),
.B(n_708),
.Y(n_10475)
);

INVx2_ASAP7_75t_SL g10476 ( 
.A(n_9635),
.Y(n_10476)
);

CKINVDCx16_ASAP7_75t_R g10477 ( 
.A(n_9710),
.Y(n_10477)
);

NAND2xp5_ASAP7_75t_L g10478 ( 
.A(n_9453),
.B(n_708),
.Y(n_10478)
);

AOI21x1_ASAP7_75t_L g10479 ( 
.A1(n_9679),
.A2(n_709),
.B(n_710),
.Y(n_10479)
);

INVxp67_ASAP7_75t_L g10480 ( 
.A(n_9604),
.Y(n_10480)
);

INVx2_ASAP7_75t_L g10481 ( 
.A(n_9479),
.Y(n_10481)
);

AOI21xp5_ASAP7_75t_L g10482 ( 
.A1(n_9651),
.A2(n_709),
.B(n_711),
.Y(n_10482)
);

AOI21xp5_ASAP7_75t_L g10483 ( 
.A1(n_9649),
.A2(n_712),
.B(n_713),
.Y(n_10483)
);

AOI21xp5_ASAP7_75t_L g10484 ( 
.A1(n_9637),
.A2(n_714),
.B(n_715),
.Y(n_10484)
);

NAND2xp5_ASAP7_75t_SL g10485 ( 
.A(n_9774),
.B(n_714),
.Y(n_10485)
);

A2O1A1Ixp33_ASAP7_75t_L g10486 ( 
.A1(n_9571),
.A2(n_9595),
.B(n_9907),
.C(n_9906),
.Y(n_10486)
);

BUFx6f_ASAP7_75t_L g10487 ( 
.A(n_9625),
.Y(n_10487)
);

AOI21xp5_ASAP7_75t_L g10488 ( 
.A1(n_9341),
.A2(n_715),
.B(n_716),
.Y(n_10488)
);

INVx1_ASAP7_75t_L g10489 ( 
.A(n_9481),
.Y(n_10489)
);

AOI22xp33_ASAP7_75t_L g10490 ( 
.A1(n_9858),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_10490)
);

NAND2xp5_ASAP7_75t_SL g10491 ( 
.A(n_9790),
.B(n_718),
.Y(n_10491)
);

A2O1A1Ixp33_ASAP7_75t_L g10492 ( 
.A1(n_9704),
.A2(n_721),
.B(n_719),
.C(n_720),
.Y(n_10492)
);

NAND2xp5_ASAP7_75t_SL g10493 ( 
.A(n_9790),
.B(n_719),
.Y(n_10493)
);

HB1xp67_ASAP7_75t_L g10494 ( 
.A(n_9724),
.Y(n_10494)
);

OAI21xp33_ASAP7_75t_L g10495 ( 
.A1(n_9737),
.A2(n_721),
.B(n_722),
.Y(n_10495)
);

CKINVDCx5p33_ASAP7_75t_R g10496 ( 
.A(n_9966),
.Y(n_10496)
);

AO21x1_ASAP7_75t_L g10497 ( 
.A1(n_9743),
.A2(n_722),
.B(n_723),
.Y(n_10497)
);

AOI22xp33_ASAP7_75t_SL g10498 ( 
.A1(n_9446),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_10498)
);

A2O1A1Ixp33_ASAP7_75t_L g10499 ( 
.A1(n_9835),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_10499)
);

AOI22xp5_ASAP7_75t_L g10500 ( 
.A1(n_9387),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_10500)
);

INVx2_ASAP7_75t_L g10501 ( 
.A(n_9486),
.Y(n_10501)
);

NAND2xp5_ASAP7_75t_L g10502 ( 
.A(n_9513),
.B(n_728),
.Y(n_10502)
);

NAND2xp5_ASAP7_75t_SL g10503 ( 
.A(n_9724),
.B(n_729),
.Y(n_10503)
);

AOI22xp5_ASAP7_75t_L g10504 ( 
.A1(n_9548),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_10504)
);

AOI21xp5_ASAP7_75t_L g10505 ( 
.A1(n_9321),
.A2(n_730),
.B(n_731),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_9521),
.Y(n_10506)
);

NOR2xp67_ASAP7_75t_L g10507 ( 
.A(n_9511),
.B(n_9705),
.Y(n_10507)
);

OR2x2_ASAP7_75t_L g10508 ( 
.A(n_9588),
.B(n_732),
.Y(n_10508)
);

NAND2xp33_ASAP7_75t_L g10509 ( 
.A(n_9306),
.B(n_733),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9538),
.Y(n_10510)
);

NAND2xp5_ASAP7_75t_L g10511 ( 
.A(n_9550),
.B(n_734),
.Y(n_10511)
);

INVx2_ASAP7_75t_L g10512 ( 
.A(n_9554),
.Y(n_10512)
);

OAI21xp33_ASAP7_75t_SL g10513 ( 
.A1(n_9350),
.A2(n_735),
.B(n_736),
.Y(n_10513)
);

AOI21xp5_ASAP7_75t_L g10514 ( 
.A1(n_9676),
.A2(n_735),
.B(n_737),
.Y(n_10514)
);

NAND2xp5_ASAP7_75t_SL g10515 ( 
.A(n_9728),
.B(n_738),
.Y(n_10515)
);

NOR3xp33_ASAP7_75t_SL g10516 ( 
.A(n_9349),
.B(n_738),
.C(n_739),
.Y(n_10516)
);

BUFx6f_ASAP7_75t_L g10517 ( 
.A(n_9684),
.Y(n_10517)
);

NAND2xp5_ASAP7_75t_SL g10518 ( 
.A(n_9728),
.B(n_740),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_L g10519 ( 
.A(n_9568),
.B(n_741),
.Y(n_10519)
);

AOI22xp5_ASAP7_75t_L g10520 ( 
.A1(n_9760),
.A2(n_9703),
.B1(n_9862),
.B2(n_9794),
.Y(n_10520)
);

NAND2xp5_ASAP7_75t_L g10521 ( 
.A(n_9599),
.B(n_741),
.Y(n_10521)
);

A2O1A1Ixp33_ASAP7_75t_L g10522 ( 
.A1(n_9841),
.A2(n_744),
.B(n_742),
.C(n_743),
.Y(n_10522)
);

CKINVDCx5p33_ASAP7_75t_R g10523 ( 
.A(n_9970),
.Y(n_10523)
);

NAND2xp5_ASAP7_75t_SL g10524 ( 
.A(n_9684),
.B(n_742),
.Y(n_10524)
);

INVx2_ASAP7_75t_L g10525 ( 
.A(n_9620),
.Y(n_10525)
);

NOR2xp33_ASAP7_75t_L g10526 ( 
.A(n_9632),
.B(n_743),
.Y(n_10526)
);

OAI22xp5_ASAP7_75t_L g10527 ( 
.A1(n_9313),
.A2(n_746),
.B1(n_744),
.B2(n_745),
.Y(n_10527)
);

NAND2xp5_ASAP7_75t_L g10528 ( 
.A(n_9624),
.B(n_9626),
.Y(n_10528)
);

AOI21xp5_ASAP7_75t_L g10529 ( 
.A1(n_9576),
.A2(n_9613),
.B(n_9591),
.Y(n_10529)
);

INVx3_ASAP7_75t_L g10530 ( 
.A(n_9460),
.Y(n_10530)
);

BUFx3_ASAP7_75t_L g10531 ( 
.A(n_9466),
.Y(n_10531)
);

NOR2xp33_ASAP7_75t_L g10532 ( 
.A(n_9655),
.B(n_746),
.Y(n_10532)
);

INVx2_ASAP7_75t_L g10533 ( 
.A(n_9633),
.Y(n_10533)
);

NOR2xp33_ASAP7_75t_R g10534 ( 
.A(n_9670),
.B(n_747),
.Y(n_10534)
);

NOR2xp33_ASAP7_75t_L g10535 ( 
.A(n_9622),
.B(n_747),
.Y(n_10535)
);

NAND2xp5_ASAP7_75t_L g10536 ( 
.A(n_9650),
.B(n_748),
.Y(n_10536)
);

AOI21xp5_ASAP7_75t_L g10537 ( 
.A1(n_9326),
.A2(n_748),
.B(n_750),
.Y(n_10537)
);

BUFx8_ASAP7_75t_SL g10538 ( 
.A(n_9723),
.Y(n_10538)
);

A2O1A1Ixp33_ASAP7_75t_L g10539 ( 
.A1(n_9843),
.A2(n_752),
.B(n_750),
.C(n_751),
.Y(n_10539)
);

NOR2xp33_ASAP7_75t_L g10540 ( 
.A(n_9646),
.B(n_751),
.Y(n_10540)
);

INVx2_ASAP7_75t_L g10541 ( 
.A(n_9658),
.Y(n_10541)
);

O2A1O1Ixp33_ASAP7_75t_L g10542 ( 
.A1(n_9846),
.A2(n_754),
.B(n_752),
.C(n_753),
.Y(n_10542)
);

NAND2xp5_ASAP7_75t_L g10543 ( 
.A(n_9662),
.B(n_754),
.Y(n_10543)
);

NAND2xp5_ASAP7_75t_SL g10544 ( 
.A(n_9353),
.B(n_755),
.Y(n_10544)
);

AOI21xp5_ASAP7_75t_L g10545 ( 
.A1(n_9304),
.A2(n_755),
.B(n_756),
.Y(n_10545)
);

NOR2xp33_ASAP7_75t_L g10546 ( 
.A(n_9409),
.B(n_756),
.Y(n_10546)
);

NAND2xp5_ASAP7_75t_L g10547 ( 
.A(n_9673),
.B(n_757),
.Y(n_10547)
);

AND2x2_ASAP7_75t_L g10548 ( 
.A(n_9951),
.B(n_758),
.Y(n_10548)
);

BUFx4f_ASAP7_75t_L g10549 ( 
.A(n_9648),
.Y(n_10549)
);

INVx3_ASAP7_75t_L g10550 ( 
.A(n_9504),
.Y(n_10550)
);

NAND2xp5_ASAP7_75t_L g10551 ( 
.A(n_9894),
.B(n_758),
.Y(n_10551)
);

AOI21xp5_ASAP7_75t_L g10552 ( 
.A1(n_9900),
.A2(n_759),
.B(n_760),
.Y(n_10552)
);

INVx1_ASAP7_75t_L g10553 ( 
.A(n_9914),
.Y(n_10553)
);

NAND2xp5_ASAP7_75t_L g10554 ( 
.A(n_9922),
.B(n_759),
.Y(n_10554)
);

INVx1_ASAP7_75t_L g10555 ( 
.A(n_9927),
.Y(n_10555)
);

BUFx2_ASAP7_75t_L g10556 ( 
.A(n_9691),
.Y(n_10556)
);

BUFx2_ASAP7_75t_L g10557 ( 
.A(n_9345),
.Y(n_10557)
);

BUFx2_ASAP7_75t_L g10558 ( 
.A(n_9903),
.Y(n_10558)
);

NOR2xp33_ASAP7_75t_R g10559 ( 
.A(n_9693),
.B(n_760),
.Y(n_10559)
);

A2O1A1Ixp33_ASAP7_75t_L g10560 ( 
.A1(n_9800),
.A2(n_764),
.B(n_761),
.C(n_763),
.Y(n_10560)
);

NAND2xp5_ASAP7_75t_SL g10561 ( 
.A(n_9424),
.B(n_761),
.Y(n_10561)
);

AOI22x1_ASAP7_75t_L g10562 ( 
.A1(n_9713),
.A2(n_9771),
.B1(n_9589),
.B2(n_9818),
.Y(n_10562)
);

AOI21xp5_ASAP7_75t_L g10563 ( 
.A1(n_9901),
.A2(n_765),
.B(n_766),
.Y(n_10563)
);

O2A1O1Ixp33_ASAP7_75t_L g10564 ( 
.A1(n_9803),
.A2(n_767),
.B(n_765),
.C(n_766),
.Y(n_10564)
);

AOI22xp5_ASAP7_75t_L g10565 ( 
.A1(n_9439),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.Y(n_10565)
);

AOI21xp5_ASAP7_75t_L g10566 ( 
.A1(n_9905),
.A2(n_771),
.B(n_772),
.Y(n_10566)
);

AOI21xp5_ASAP7_75t_L g10567 ( 
.A1(n_9910),
.A2(n_771),
.B(n_772),
.Y(n_10567)
);

INVx2_ASAP7_75t_L g10568 ( 
.A(n_9949),
.Y(n_10568)
);

NOR2xp33_ASAP7_75t_SL g10569 ( 
.A(n_9476),
.B(n_773),
.Y(n_10569)
);

BUFx6f_ASAP7_75t_L g10570 ( 
.A(n_9497),
.Y(n_10570)
);

INVx2_ASAP7_75t_L g10571 ( 
.A(n_9953),
.Y(n_10571)
);

INVx5_ASAP7_75t_L g10572 ( 
.A(n_9594),
.Y(n_10572)
);

NOR2xp33_ASAP7_75t_R g10573 ( 
.A(n_9575),
.B(n_773),
.Y(n_10573)
);

INVx2_ASAP7_75t_L g10574 ( 
.A(n_9967),
.Y(n_10574)
);

INVx2_ASAP7_75t_L g10575 ( 
.A(n_9978),
.Y(n_10575)
);

AND2x4_ASAP7_75t_L g10576 ( 
.A(n_9969),
.B(n_774),
.Y(n_10576)
);

AOI21xp33_ASAP7_75t_L g10577 ( 
.A1(n_9850),
.A2(n_774),
.B(n_775),
.Y(n_10577)
);

A2O1A1Ixp33_ASAP7_75t_L g10578 ( 
.A1(n_9853),
.A2(n_778),
.B(n_775),
.C(n_776),
.Y(n_10578)
);

CKINVDCx5p33_ASAP7_75t_R g10579 ( 
.A(n_9502),
.Y(n_10579)
);

O2A1O1Ixp33_ASAP7_75t_L g10580 ( 
.A1(n_9762),
.A2(n_779),
.B(n_776),
.C(n_778),
.Y(n_10580)
);

OAI22xp5_ASAP7_75t_L g10581 ( 
.A1(n_9664),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_10581)
);

INVx2_ASAP7_75t_L g10582 ( 
.A(n_9683),
.Y(n_10582)
);

NOR2xp33_ASAP7_75t_L g10583 ( 
.A(n_9648),
.B(n_780),
.Y(n_10583)
);

INVx2_ASAP7_75t_L g10584 ( 
.A(n_9689),
.Y(n_10584)
);

INVx1_ASAP7_75t_L g10585 ( 
.A(n_9729),
.Y(n_10585)
);

NAND2xp5_ASAP7_75t_L g10586 ( 
.A(n_9736),
.B(n_781),
.Y(n_10586)
);

AOI21xp5_ASAP7_75t_L g10587 ( 
.A1(n_9928),
.A2(n_784),
.B(n_785),
.Y(n_10587)
);

NAND2xp5_ASAP7_75t_SL g10588 ( 
.A(n_9594),
.B(n_784),
.Y(n_10588)
);

INVx1_ASAP7_75t_L g10589 ( 
.A(n_9354),
.Y(n_10589)
);

OAI21x1_ASAP7_75t_L g10590 ( 
.A1(n_9359),
.A2(n_786),
.B(n_787),
.Y(n_10590)
);

NAND2xp5_ASAP7_75t_L g10591 ( 
.A(n_9660),
.B(n_786),
.Y(n_10591)
);

NAND2xp5_ASAP7_75t_L g10592 ( 
.A(n_9936),
.B(n_787),
.Y(n_10592)
);

INVx1_ASAP7_75t_L g10593 ( 
.A(n_9360),
.Y(n_10593)
);

AOI22xp5_ASAP7_75t_L g10594 ( 
.A1(n_9565),
.A2(n_791),
.B1(n_788),
.B2(n_789),
.Y(n_10594)
);

A2O1A1Ixp33_ASAP7_75t_L g10595 ( 
.A1(n_9763),
.A2(n_793),
.B(n_788),
.C(n_792),
.Y(n_10595)
);

INVx1_ASAP7_75t_L g10596 ( 
.A(n_9370),
.Y(n_10596)
);

INVx1_ASAP7_75t_SL g10597 ( 
.A(n_9602),
.Y(n_10597)
);

AOI21xp5_ASAP7_75t_L g10598 ( 
.A1(n_9940),
.A2(n_792),
.B(n_793),
.Y(n_10598)
);

OR2x2_ASAP7_75t_L g10599 ( 
.A(n_9467),
.B(n_794),
.Y(n_10599)
);

INVx3_ASAP7_75t_L g10600 ( 
.A(n_9352),
.Y(n_10600)
);

NAND2xp5_ASAP7_75t_SL g10601 ( 
.A(n_9563),
.B(n_794),
.Y(n_10601)
);

NAND2xp5_ASAP7_75t_L g10602 ( 
.A(n_9943),
.B(n_9944),
.Y(n_10602)
);

O2A1O1Ixp33_ASAP7_75t_L g10603 ( 
.A1(n_9855),
.A2(n_797),
.B(n_795),
.C(n_796),
.Y(n_10603)
);

BUFx6f_ASAP7_75t_L g10604 ( 
.A(n_9600),
.Y(n_10604)
);

OAI22xp5_ASAP7_75t_L g10605 ( 
.A1(n_9680),
.A2(n_800),
.B1(n_795),
.B2(n_799),
.Y(n_10605)
);

AOI21xp5_ASAP7_75t_L g10606 ( 
.A1(n_9954),
.A2(n_799),
.B(n_801),
.Y(n_10606)
);

AO32x1_ASAP7_75t_L g10607 ( 
.A1(n_9826),
.A2(n_804),
.A3(n_802),
.B1(n_803),
.B2(n_805),
.Y(n_10607)
);

AND2x2_ASAP7_75t_L g10608 ( 
.A(n_9952),
.B(n_802),
.Y(n_10608)
);

NOR2xp33_ASAP7_75t_L g10609 ( 
.A(n_9523),
.B(n_804),
.Y(n_10609)
);

AND2x4_ASAP7_75t_L g10610 ( 
.A(n_9663),
.B(n_806),
.Y(n_10610)
);

NAND2xp5_ASAP7_75t_SL g10611 ( 
.A(n_9600),
.B(n_806),
.Y(n_10611)
);

NAND2xp5_ASAP7_75t_L g10612 ( 
.A(n_9980),
.B(n_807),
.Y(n_10612)
);

OAI21x1_ASAP7_75t_SL g10613 ( 
.A1(n_9375),
.A2(n_807),
.B(n_808),
.Y(n_10613)
);

NOR2xp33_ASAP7_75t_L g10614 ( 
.A(n_9945),
.B(n_808),
.Y(n_10614)
);

AOI22xp33_ASAP7_75t_L g10615 ( 
.A1(n_9986),
.A2(n_811),
.B1(n_809),
.B2(n_810),
.Y(n_10615)
);

BUFx6f_ASAP7_75t_L g10616 ( 
.A(n_9364),
.Y(n_10616)
);

NAND2xp5_ASAP7_75t_SL g10617 ( 
.A(n_9981),
.B(n_809),
.Y(n_10617)
);

NAND2xp5_ASAP7_75t_L g10618 ( 
.A(n_9987),
.B(n_811),
.Y(n_10618)
);

BUFx8_ASAP7_75t_SL g10619 ( 
.A(n_9962),
.Y(n_10619)
);

INVx4_ASAP7_75t_L g10620 ( 
.A(n_9330),
.Y(n_10620)
);

NOR2xp33_ASAP7_75t_L g10621 ( 
.A(n_9647),
.B(n_812),
.Y(n_10621)
);

AND2x4_ASAP7_75t_L g10622 ( 
.A(n_9909),
.B(n_9912),
.Y(n_10622)
);

INVxp67_ASAP7_75t_SL g10623 ( 
.A(n_9378),
.Y(n_10623)
);

OAI21xp5_ASAP7_75t_L g10624 ( 
.A1(n_9988),
.A2(n_812),
.B(n_813),
.Y(n_10624)
);

A2O1A1Ixp33_ASAP7_75t_L g10625 ( 
.A1(n_9590),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_10625)
);

BUFx4f_ASAP7_75t_L g10626 ( 
.A(n_9317),
.Y(n_10626)
);

NAND2xp5_ASAP7_75t_L g10627 ( 
.A(n_9644),
.B(n_814),
.Y(n_10627)
);

NAND2x1p5_ASAP7_75t_L g10628 ( 
.A(n_9539),
.B(n_815),
.Y(n_10628)
);

NAND2xp5_ASAP7_75t_SL g10629 ( 
.A(n_9593),
.B(n_816),
.Y(n_10629)
);

AOI22xp5_ASAP7_75t_L g10630 ( 
.A1(n_9331),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_10630)
);

CKINVDCx6p67_ASAP7_75t_R g10631 ( 
.A(n_9470),
.Y(n_10631)
);

A2O1A1Ixp33_ASAP7_75t_L g10632 ( 
.A1(n_9598),
.A2(n_820),
.B(n_817),
.C(n_819),
.Y(n_10632)
);

CKINVDCx5p33_ASAP7_75t_R g10633 ( 
.A(n_10009),
.Y(n_10633)
);

INVx2_ASAP7_75t_L g10634 ( 
.A(n_10173),
.Y(n_10634)
);

OAI21x1_ASAP7_75t_L g10635 ( 
.A1(n_10380),
.A2(n_9381),
.B(n_9380),
.Y(n_10635)
);

AOI21xp5_ASAP7_75t_L g10636 ( 
.A1(n_9997),
.A2(n_9390),
.B(n_9389),
.Y(n_10636)
);

NAND2xp5_ASAP7_75t_L g10637 ( 
.A(n_10200),
.B(n_9612),
.Y(n_10637)
);

OAI21x1_ASAP7_75t_L g10638 ( 
.A1(n_10016),
.A2(n_9418),
.B(n_9410),
.Y(n_10638)
);

NAND2xp5_ASAP7_75t_L g10639 ( 
.A(n_10623),
.B(n_10205),
.Y(n_10639)
);

BUFx10_ASAP7_75t_L g10640 ( 
.A(n_10466),
.Y(n_10640)
);

CKINVDCx5p33_ASAP7_75t_R g10641 ( 
.A(n_10247),
.Y(n_10641)
);

AOI21xp5_ASAP7_75t_L g10642 ( 
.A1(n_10026),
.A2(n_9435),
.B(n_9429),
.Y(n_10642)
);

OR2x2_ASAP7_75t_L g10643 ( 
.A(n_10014),
.B(n_9930),
.Y(n_10643)
);

INVx4_ASAP7_75t_L g10644 ( 
.A(n_10579),
.Y(n_10644)
);

AO31x2_ASAP7_75t_L g10645 ( 
.A1(n_9998),
.A2(n_9499),
.A3(n_9518),
.B(n_9477),
.Y(n_10645)
);

INVx1_ASAP7_75t_L g10646 ( 
.A(n_10248),
.Y(n_10646)
);

NOR2xp33_ASAP7_75t_L g10647 ( 
.A(n_10214),
.B(n_9740),
.Y(n_10647)
);

INVx2_ASAP7_75t_SL g10648 ( 
.A(n_10275),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_10281),
.Y(n_10649)
);

OAI21xp5_ASAP7_75t_L g10650 ( 
.A1(n_10067),
.A2(n_9630),
.B(n_9567),
.Y(n_10650)
);

NAND2xp5_ASAP7_75t_L g10651 ( 
.A(n_10044),
.B(n_9558),
.Y(n_10651)
);

INVx1_ASAP7_75t_L g10652 ( 
.A(n_10149),
.Y(n_10652)
);

NAND2xp5_ASAP7_75t_L g10653 ( 
.A(n_10158),
.B(n_9718),
.Y(n_10653)
);

INVx1_ASAP7_75t_L g10654 ( 
.A(n_10199),
.Y(n_10654)
);

BUFx6f_ASAP7_75t_L g10655 ( 
.A(n_10083),
.Y(n_10655)
);

INVx2_ASAP7_75t_SL g10656 ( 
.A(n_10368),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_10211),
.Y(n_10657)
);

NAND2xp5_ASAP7_75t_L g10658 ( 
.A(n_10163),
.B(n_9712),
.Y(n_10658)
);

AO31x2_ASAP7_75t_L g10659 ( 
.A1(n_10055),
.A2(n_9739),
.A3(n_822),
.B(n_820),
.Y(n_10659)
);

INVx1_ASAP7_75t_L g10660 ( 
.A(n_10218),
.Y(n_10660)
);

BUFx3_ASAP7_75t_L g10661 ( 
.A(n_10020),
.Y(n_10661)
);

AOI21xp5_ASAP7_75t_L g10662 ( 
.A1(n_10048),
.A2(n_9426),
.B(n_9412),
.Y(n_10662)
);

OAI21x1_ASAP7_75t_L g10663 ( 
.A1(n_10332),
.A2(n_9570),
.B(n_9338),
.Y(n_10663)
);

NAND2xp5_ASAP7_75t_SL g10664 ( 
.A(n_10394),
.B(n_9618),
.Y(n_10664)
);

INVx2_ASAP7_75t_SL g10665 ( 
.A(n_10453),
.Y(n_10665)
);

CKINVDCx11_ASAP7_75t_R g10666 ( 
.A(n_10043),
.Y(n_10666)
);

NAND2xp5_ASAP7_75t_L g10667 ( 
.A(n_10184),
.B(n_9721),
.Y(n_10667)
);

OAI21x1_ASAP7_75t_L g10668 ( 
.A1(n_10186),
.A2(n_9348),
.B(n_9335),
.Y(n_10668)
);

OAI21xp5_ASAP7_75t_L g10669 ( 
.A1(n_10141),
.A2(n_10134),
.B(n_10098),
.Y(n_10669)
);

NAND2xp5_ASAP7_75t_L g10670 ( 
.A(n_10122),
.B(n_9431),
.Y(n_10670)
);

INVx1_ASAP7_75t_SL g10671 ( 
.A(n_10221),
.Y(n_10671)
);

AND2x4_ASAP7_75t_L g10672 ( 
.A(n_10041),
.B(n_9386),
.Y(n_10672)
);

INVx2_ASAP7_75t_SL g10673 ( 
.A(n_10464),
.Y(n_10673)
);

NAND2xp5_ASAP7_75t_L g10674 ( 
.A(n_10077),
.B(n_9413),
.Y(n_10674)
);

NAND2xp5_ASAP7_75t_L g10675 ( 
.A(n_10038),
.B(n_9427),
.Y(n_10675)
);

OR2x6_ASAP7_75t_L g10676 ( 
.A(n_10288),
.B(n_9384),
.Y(n_10676)
);

BUFx6f_ASAP7_75t_L g10677 ( 
.A(n_10083),
.Y(n_10677)
);

BUFx3_ASAP7_75t_L g10678 ( 
.A(n_10115),
.Y(n_10678)
);

NOR2xp33_ASAP7_75t_R g10679 ( 
.A(n_10244),
.B(n_9432),
.Y(n_10679)
);

OAI21x1_ASAP7_75t_L g10680 ( 
.A1(n_10529),
.A2(n_9462),
.B(n_9458),
.Y(n_10680)
);

OAI21x1_ASAP7_75t_L g10681 ( 
.A1(n_10161),
.A2(n_9500),
.B(n_9487),
.Y(n_10681)
);

NAND2xp5_ASAP7_75t_L g10682 ( 
.A(n_9994),
.B(n_9541),
.Y(n_10682)
);

OAI21x1_ASAP7_75t_L g10683 ( 
.A1(n_10265),
.A2(n_821),
.B(n_822),
.Y(n_10683)
);

AND2x2_ASAP7_75t_L g10684 ( 
.A(n_10006),
.B(n_823),
.Y(n_10684)
);

A2O1A1Ixp33_ASAP7_75t_L g10685 ( 
.A1(n_10024),
.A2(n_825),
.B(n_823),
.C(n_824),
.Y(n_10685)
);

CKINVDCx14_ASAP7_75t_R g10686 ( 
.A(n_10286),
.Y(n_10686)
);

O2A1O1Ixp33_ASAP7_75t_L g10687 ( 
.A1(n_10093),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_10687)
);

NAND3x1_ASAP7_75t_L g10688 ( 
.A(n_10614),
.B(n_826),
.C(n_827),
.Y(n_10688)
);

AND2x2_ASAP7_75t_L g10689 ( 
.A(n_10155),
.B(n_827),
.Y(n_10689)
);

O2A1O1Ixp33_ASAP7_75t_SL g10690 ( 
.A1(n_10033),
.A2(n_830),
.B(n_828),
.C(n_829),
.Y(n_10690)
);

INVx2_ASAP7_75t_SL g10691 ( 
.A(n_10469),
.Y(n_10691)
);

NOR2xp67_ASAP7_75t_L g10692 ( 
.A(n_10003),
.B(n_828),
.Y(n_10692)
);

A2O1A1Ixp33_ASAP7_75t_L g10693 ( 
.A1(n_10237),
.A2(n_831),
.B(n_829),
.C(n_830),
.Y(n_10693)
);

OAI21x1_ASAP7_75t_L g10694 ( 
.A1(n_10152),
.A2(n_10080),
.B(n_10320),
.Y(n_10694)
);

NAND2xp5_ASAP7_75t_SL g10695 ( 
.A(n_10172),
.B(n_831),
.Y(n_10695)
);

INVx1_ASAP7_75t_L g10696 ( 
.A(n_10227),
.Y(n_10696)
);

OAI21x1_ASAP7_75t_L g10697 ( 
.A1(n_10166),
.A2(n_832),
.B(n_833),
.Y(n_10697)
);

AOI21xp5_ASAP7_75t_L g10698 ( 
.A1(n_10005),
.A2(n_832),
.B(n_833),
.Y(n_10698)
);

AOI21xp5_ASAP7_75t_L g10699 ( 
.A1(n_10070),
.A2(n_834),
.B(n_835),
.Y(n_10699)
);

NOR2xp33_ASAP7_75t_SL g10700 ( 
.A(n_10133),
.B(n_836),
.Y(n_10700)
);

INVx1_ASAP7_75t_L g10701 ( 
.A(n_10232),
.Y(n_10701)
);

OAI21x1_ASAP7_75t_L g10702 ( 
.A1(n_10170),
.A2(n_836),
.B(n_837),
.Y(n_10702)
);

BUFx2_ASAP7_75t_L g10703 ( 
.A(n_10160),
.Y(n_10703)
);

OR2x2_ASAP7_75t_L g10704 ( 
.A(n_10004),
.B(n_837),
.Y(n_10704)
);

AND2x2_ASAP7_75t_L g10705 ( 
.A(n_10371),
.B(n_838),
.Y(n_10705)
);

AOI21xp5_ASAP7_75t_L g10706 ( 
.A1(n_10008),
.A2(n_839),
.B(n_840),
.Y(n_10706)
);

AOI21xp5_ASAP7_75t_SL g10707 ( 
.A1(n_9995),
.A2(n_839),
.B(n_840),
.Y(n_10707)
);

NAND2xp5_ASAP7_75t_L g10708 ( 
.A(n_10035),
.B(n_10042),
.Y(n_10708)
);

OAI22xp5_ASAP7_75t_L g10709 ( 
.A1(n_10010),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_10235),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_L g10711 ( 
.A(n_10438),
.B(n_842),
.Y(n_10711)
);

AND2x4_ASAP7_75t_L g10712 ( 
.A(n_10435),
.B(n_844),
.Y(n_10712)
);

OAI21x1_ASAP7_75t_L g10713 ( 
.A1(n_10590),
.A2(n_844),
.B(n_845),
.Y(n_10713)
);

INVx3_ASAP7_75t_L g10714 ( 
.A(n_10096),
.Y(n_10714)
);

O2A1O1Ixp5_ASAP7_75t_L g10715 ( 
.A1(n_10047),
.A2(n_847),
.B(n_845),
.C(n_846),
.Y(n_10715)
);

AOI221xp5_ASAP7_75t_L g10716 ( 
.A1(n_10261),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.C(n_849),
.Y(n_10716)
);

NAND2xp5_ASAP7_75t_L g10717 ( 
.A(n_10462),
.B(n_850),
.Y(n_10717)
);

O2A1O1Ixp5_ASAP7_75t_L g10718 ( 
.A1(n_10171),
.A2(n_10178),
.B(n_10027),
.C(n_10146),
.Y(n_10718)
);

AND2x2_ASAP7_75t_L g10719 ( 
.A(n_10223),
.B(n_10313),
.Y(n_10719)
);

OAI21x1_ASAP7_75t_L g10720 ( 
.A1(n_10327),
.A2(n_850),
.B(n_851),
.Y(n_10720)
);

NOR2x1_ASAP7_75t_SL g10721 ( 
.A(n_10151),
.B(n_852),
.Y(n_10721)
);

INVx2_ASAP7_75t_L g10722 ( 
.A(n_10187),
.Y(n_10722)
);

OAI21x1_ASAP7_75t_L g10723 ( 
.A1(n_10032),
.A2(n_853),
.B(n_854),
.Y(n_10723)
);

INVx5_ASAP7_75t_L g10724 ( 
.A(n_10300),
.Y(n_10724)
);

AO31x2_ASAP7_75t_L g10725 ( 
.A1(n_10022),
.A2(n_856),
.A3(n_854),
.B(n_855),
.Y(n_10725)
);

NAND3x1_ASAP7_75t_L g10726 ( 
.A(n_10535),
.B(n_855),
.C(n_856),
.Y(n_10726)
);

NAND2xp5_ASAP7_75t_L g10727 ( 
.A(n_10012),
.B(n_857),
.Y(n_10727)
);

NAND2xp5_ASAP7_75t_SL g10728 ( 
.A(n_10068),
.B(n_857),
.Y(n_10728)
);

INVx1_ASAP7_75t_L g10729 ( 
.A(n_10236),
.Y(n_10729)
);

NAND2xp33_ASAP7_75t_L g10730 ( 
.A(n_10375),
.B(n_858),
.Y(n_10730)
);

OAI21xp5_ASAP7_75t_L g10731 ( 
.A1(n_10100),
.A2(n_858),
.B(n_859),
.Y(n_10731)
);

INVx8_ASAP7_75t_L g10732 ( 
.A(n_10466),
.Y(n_10732)
);

OAI21xp5_ASAP7_75t_L g10733 ( 
.A1(n_10329),
.A2(n_859),
.B(n_861),
.Y(n_10733)
);

OAI21xp5_ASAP7_75t_L g10734 ( 
.A1(n_10361),
.A2(n_862),
.B(n_863),
.Y(n_10734)
);

AOI21xp5_ASAP7_75t_L g10735 ( 
.A1(n_10013),
.A2(n_862),
.B(n_864),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_10239),
.Y(n_10736)
);

NAND2xp5_ASAP7_75t_SL g10737 ( 
.A(n_10312),
.B(n_865),
.Y(n_10737)
);

NOR2xp33_ASAP7_75t_L g10738 ( 
.A(n_10602),
.B(n_866),
.Y(n_10738)
);

AOI21xp5_ASAP7_75t_L g10739 ( 
.A1(n_10017),
.A2(n_866),
.B(n_867),
.Y(n_10739)
);

OA21x2_ASAP7_75t_L g10740 ( 
.A1(n_10428),
.A2(n_868),
.B(n_869),
.Y(n_10740)
);

AOI21xp5_ASAP7_75t_L g10741 ( 
.A1(n_10054),
.A2(n_868),
.B(n_870),
.Y(n_10741)
);

OAI21x1_ASAP7_75t_L g10742 ( 
.A1(n_10426),
.A2(n_870),
.B(n_871),
.Y(n_10742)
);

BUFx2_ASAP7_75t_L g10743 ( 
.A(n_10415),
.Y(n_10743)
);

INVx1_ASAP7_75t_SL g10744 ( 
.A(n_10597),
.Y(n_10744)
);

INVx1_ASAP7_75t_SL g10745 ( 
.A(n_10457),
.Y(n_10745)
);

NAND2xp5_ASAP7_75t_L g10746 ( 
.A(n_10015),
.B(n_871),
.Y(n_10746)
);

OR2x2_ASAP7_75t_L g10747 ( 
.A(n_10029),
.B(n_872),
.Y(n_10747)
);

NAND2x1p5_ASAP7_75t_L g10748 ( 
.A(n_10557),
.B(n_872),
.Y(n_10748)
);

A2O1A1Ixp33_ASAP7_75t_L g10749 ( 
.A1(n_10120),
.A2(n_875),
.B(n_873),
.C(n_874),
.Y(n_10749)
);

AOI221xp5_ASAP7_75t_L g10750 ( 
.A1(n_10424),
.A2(n_875),
.B1(n_873),
.B2(n_874),
.C(n_876),
.Y(n_10750)
);

INVx1_ASAP7_75t_L g10751 ( 
.A(n_10258),
.Y(n_10751)
);

AOI21xp5_ASAP7_75t_L g10752 ( 
.A1(n_10304),
.A2(n_877),
.B(n_878),
.Y(n_10752)
);

AOI221x1_ASAP7_75t_L g10753 ( 
.A1(n_10079),
.A2(n_880),
.B1(n_877),
.B2(n_879),
.C(n_881),
.Y(n_10753)
);

NOR4xp25_ASAP7_75t_L g10754 ( 
.A(n_10425),
.B(n_881),
.C(n_879),
.D(n_880),
.Y(n_10754)
);

INVxp67_ASAP7_75t_L g10755 ( 
.A(n_10386),
.Y(n_10755)
);

OAI21x1_ASAP7_75t_L g10756 ( 
.A1(n_10528),
.A2(n_882),
.B(n_883),
.Y(n_10756)
);

AOI31xp67_ASAP7_75t_L g10757 ( 
.A1(n_10594),
.A2(n_10136),
.A3(n_10143),
.B(n_10135),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_SL g10758 ( 
.A(n_10305),
.B(n_882),
.Y(n_10758)
);

OAI22xp5_ASAP7_75t_L g10759 ( 
.A1(n_10206),
.A2(n_10500),
.B1(n_10504),
.B2(n_10140),
.Y(n_10759)
);

CKINVDCx11_ASAP7_75t_R g10760 ( 
.A(n_10011),
.Y(n_10760)
);

AOI21xp5_ASAP7_75t_L g10761 ( 
.A1(n_10073),
.A2(n_10091),
.B(n_10509),
.Y(n_10761)
);

AOI22xp5_ASAP7_75t_L g10762 ( 
.A1(n_10092),
.A2(n_885),
.B1(n_883),
.B2(n_884),
.Y(n_10762)
);

BUFx6f_ASAP7_75t_L g10763 ( 
.A(n_10115),
.Y(n_10763)
);

NAND2xp5_ASAP7_75t_SL g10764 ( 
.A(n_10600),
.B(n_884),
.Y(n_10764)
);

NAND2xp5_ASAP7_75t_SL g10765 ( 
.A(n_10486),
.B(n_885),
.Y(n_10765)
);

INVx1_ASAP7_75t_L g10766 ( 
.A(n_10273),
.Y(n_10766)
);

NAND2xp5_ASAP7_75t_L g10767 ( 
.A(n_10030),
.B(n_886),
.Y(n_10767)
);

BUFx2_ASAP7_75t_L g10768 ( 
.A(n_10339),
.Y(n_10768)
);

BUFx2_ASAP7_75t_L g10769 ( 
.A(n_10343),
.Y(n_10769)
);

INVx2_ASAP7_75t_L g10770 ( 
.A(n_10189),
.Y(n_10770)
);

AOI21xp5_ASAP7_75t_L g10771 ( 
.A1(n_10191),
.A2(n_886),
.B(n_887),
.Y(n_10771)
);

OAI21xp5_ASAP7_75t_L g10772 ( 
.A1(n_10369),
.A2(n_887),
.B(n_888),
.Y(n_10772)
);

BUFx2_ASAP7_75t_L g10773 ( 
.A(n_10432),
.Y(n_10773)
);

OA21x2_ASAP7_75t_L g10774 ( 
.A1(n_10334),
.A2(n_888),
.B(n_889),
.Y(n_10774)
);

OAI21x1_ASAP7_75t_L g10775 ( 
.A1(n_10408),
.A2(n_889),
.B(n_890),
.Y(n_10775)
);

CKINVDCx14_ASAP7_75t_R g10776 ( 
.A(n_10534),
.Y(n_10776)
);

HB1xp67_ASAP7_75t_L g10777 ( 
.A(n_10046),
.Y(n_10777)
);

AOI21xp5_ASAP7_75t_L g10778 ( 
.A1(n_10263),
.A2(n_890),
.B(n_891),
.Y(n_10778)
);

NAND3xp33_ASAP7_75t_L g10779 ( 
.A(n_10542),
.B(n_892),
.C(n_893),
.Y(n_10779)
);

INVx3_ASAP7_75t_L g10780 ( 
.A(n_10096),
.Y(n_10780)
);

AND2x2_ASAP7_75t_L g10781 ( 
.A(n_10558),
.B(n_10441),
.Y(n_10781)
);

O2A1O1Ixp5_ASAP7_75t_SL g10782 ( 
.A1(n_10162),
.A2(n_894),
.B(n_892),
.C(n_893),
.Y(n_10782)
);

OAI21xp5_ASAP7_75t_L g10783 ( 
.A1(n_10384),
.A2(n_894),
.B(n_895),
.Y(n_10783)
);

INVx5_ASAP7_75t_L g10784 ( 
.A(n_10538),
.Y(n_10784)
);

OAI21xp5_ASAP7_75t_L g10785 ( 
.A1(n_10505),
.A2(n_10545),
.B(n_10537),
.Y(n_10785)
);

INVx2_ASAP7_75t_L g10786 ( 
.A(n_10196),
.Y(n_10786)
);

BUFx3_ASAP7_75t_L g10787 ( 
.A(n_10144),
.Y(n_10787)
);

INVx2_ASAP7_75t_L g10788 ( 
.A(n_10213),
.Y(n_10788)
);

AO21x1_ASAP7_75t_L g10789 ( 
.A1(n_10209),
.A2(n_10001),
.B(n_10224),
.Y(n_10789)
);

NAND2xp5_ASAP7_75t_L g10790 ( 
.A(n_10051),
.B(n_895),
.Y(n_10790)
);

INVx3_ASAP7_75t_L g10791 ( 
.A(n_10531),
.Y(n_10791)
);

NAND2xp5_ASAP7_75t_L g10792 ( 
.A(n_10062),
.B(n_896),
.Y(n_10792)
);

AO32x2_ASAP7_75t_L g10793 ( 
.A1(n_10231),
.A2(n_899),
.A3(n_897),
.B1(n_898),
.B2(n_900),
.Y(n_10793)
);

BUFx10_ASAP7_75t_L g10794 ( 
.A(n_10072),
.Y(n_10794)
);

AOI21xp5_ASAP7_75t_L g10795 ( 
.A1(n_10157),
.A2(n_897),
.B(n_898),
.Y(n_10795)
);

OAI21xp5_ASAP7_75t_L g10796 ( 
.A1(n_10552),
.A2(n_899),
.B(n_900),
.Y(n_10796)
);

AOI21xp33_ASAP7_75t_L g10797 ( 
.A1(n_10293),
.A2(n_901),
.B(n_902),
.Y(n_10797)
);

INVxp67_ASAP7_75t_SL g10798 ( 
.A(n_10473),
.Y(n_10798)
);

AOI21xp5_ASAP7_75t_L g10799 ( 
.A1(n_10341),
.A2(n_901),
.B(n_903),
.Y(n_10799)
);

NAND2xp5_ASAP7_75t_L g10800 ( 
.A(n_10074),
.B(n_904),
.Y(n_10800)
);

OA21x2_ASAP7_75t_L g10801 ( 
.A1(n_10279),
.A2(n_904),
.B(n_905),
.Y(n_10801)
);

NAND2x1_ASAP7_75t_L g10802 ( 
.A(n_10103),
.B(n_905),
.Y(n_10802)
);

OAI21xp5_ASAP7_75t_L g10803 ( 
.A1(n_10563),
.A2(n_906),
.B(n_907),
.Y(n_10803)
);

OAI21x1_ASAP7_75t_L g10804 ( 
.A1(n_10459),
.A2(n_910),
.B(n_911),
.Y(n_10804)
);

A2O1A1Ixp33_ASAP7_75t_L g10805 ( 
.A1(n_10322),
.A2(n_912),
.B(n_910),
.C(n_911),
.Y(n_10805)
);

INVxp67_ASAP7_75t_SL g10806 ( 
.A(n_10114),
.Y(n_10806)
);

OAI21x1_ASAP7_75t_L g10807 ( 
.A1(n_10255),
.A2(n_912),
.B(n_913),
.Y(n_10807)
);

BUFx6f_ASAP7_75t_L g10808 ( 
.A(n_10144),
.Y(n_10808)
);

OAI22xp5_ASAP7_75t_L g10809 ( 
.A1(n_10393),
.A2(n_915),
.B1(n_913),
.B2(n_914),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_10289),
.Y(n_10810)
);

AOI21xp33_ASAP7_75t_L g10811 ( 
.A1(n_10335),
.A2(n_914),
.B(n_915),
.Y(n_10811)
);

NAND2xp5_ASAP7_75t_L g10812 ( 
.A(n_10118),
.B(n_916),
.Y(n_10812)
);

OA21x2_ASAP7_75t_L g10813 ( 
.A1(n_10295),
.A2(n_916),
.B(n_917),
.Y(n_10813)
);

A2O1A1Ixp33_ASAP7_75t_L g10814 ( 
.A1(n_10564),
.A2(n_919),
.B(n_917),
.C(n_918),
.Y(n_10814)
);

CKINVDCx20_ASAP7_75t_R g10815 ( 
.A(n_10102),
.Y(n_10815)
);

AO32x2_ASAP7_75t_L g10816 ( 
.A1(n_10034),
.A2(n_921),
.A3(n_919),
.B1(n_920),
.B2(n_922),
.Y(n_10816)
);

AND2x2_ASAP7_75t_L g10817 ( 
.A(n_10124),
.B(n_921),
.Y(n_10817)
);

OAI21xp5_ASAP7_75t_L g10818 ( 
.A1(n_10566),
.A2(n_922),
.B(n_923),
.Y(n_10818)
);

INVx2_ASAP7_75t_L g10819 ( 
.A(n_10238),
.Y(n_10819)
);

NOR2xp33_ASAP7_75t_L g10820 ( 
.A(n_10019),
.B(n_923),
.Y(n_10820)
);

NAND2xp5_ASAP7_75t_L g10821 ( 
.A(n_10125),
.B(n_924),
.Y(n_10821)
);

AND2x4_ASAP7_75t_L g10822 ( 
.A(n_10378),
.B(n_924),
.Y(n_10822)
);

AOI21x1_ASAP7_75t_L g10823 ( 
.A1(n_10479),
.A2(n_925),
.B(n_926),
.Y(n_10823)
);

OA21x2_ASAP7_75t_L g10824 ( 
.A1(n_10299),
.A2(n_925),
.B(n_927),
.Y(n_10824)
);

AOI221x1_ASAP7_75t_L g10825 ( 
.A1(n_10137),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.C(n_930),
.Y(n_10825)
);

AOI21xp5_ASAP7_75t_L g10826 ( 
.A1(n_10626),
.A2(n_928),
.B(n_929),
.Y(n_10826)
);

INVx2_ASAP7_75t_L g10827 ( 
.A(n_10242),
.Y(n_10827)
);

OR2x2_ASAP7_75t_L g10828 ( 
.A(n_10139),
.B(n_930),
.Y(n_10828)
);

NAND3xp33_ASAP7_75t_L g10829 ( 
.A(n_10580),
.B(n_10366),
.C(n_10360),
.Y(n_10829)
);

AOI21xp5_ASAP7_75t_L g10830 ( 
.A1(n_10230),
.A2(n_931),
.B(n_932),
.Y(n_10830)
);

NOR2xp33_ASAP7_75t_L g10831 ( 
.A(n_10147),
.B(n_10159),
.Y(n_10831)
);

NAND2xp5_ASAP7_75t_L g10832 ( 
.A(n_10381),
.B(n_10372),
.Y(n_10832)
);

OAI21x1_ASAP7_75t_L g10833 ( 
.A1(n_10198),
.A2(n_931),
.B(n_933),
.Y(n_10833)
);

INVx1_ASAP7_75t_L g10834 ( 
.A(n_10301),
.Y(n_10834)
);

OA21x2_ASAP7_75t_L g10835 ( 
.A1(n_10307),
.A2(n_933),
.B(n_935),
.Y(n_10835)
);

AND2x4_ASAP7_75t_L g10836 ( 
.A(n_10556),
.B(n_936),
.Y(n_10836)
);

AO31x2_ASAP7_75t_L g10837 ( 
.A1(n_10497),
.A2(n_938),
.A3(n_936),
.B(n_937),
.Y(n_10837)
);

CKINVDCx20_ASAP7_75t_R g10838 ( 
.A(n_10225),
.Y(n_10838)
);

CKINVDCx20_ASAP7_75t_R g10839 ( 
.A(n_10357),
.Y(n_10839)
);

OAI21xp5_ASAP7_75t_L g10840 ( 
.A1(n_10567),
.A2(n_937),
.B(n_938),
.Y(n_10840)
);

AOI21xp5_ASAP7_75t_L g10841 ( 
.A1(n_10391),
.A2(n_939),
.B(n_941),
.Y(n_10841)
);

INVx1_ASAP7_75t_L g10842 ( 
.A(n_10337),
.Y(n_10842)
);

OAI21x1_ASAP7_75t_L g10843 ( 
.A1(n_10355),
.A2(n_939),
.B(n_941),
.Y(n_10843)
);

OAI21xp5_ASAP7_75t_L g10844 ( 
.A1(n_10587),
.A2(n_942),
.B(n_943),
.Y(n_10844)
);

AOI21xp5_ASAP7_75t_L g10845 ( 
.A1(n_10228),
.A2(n_943),
.B(n_944),
.Y(n_10845)
);

OAI21xp5_ASAP7_75t_L g10846 ( 
.A1(n_10598),
.A2(n_945),
.B(n_946),
.Y(n_10846)
);

OAI22xp5_ASAP7_75t_L g10847 ( 
.A1(n_10400),
.A2(n_10303),
.B1(n_10180),
.B2(n_10283),
.Y(n_10847)
);

AND2x4_ASAP7_75t_L g10848 ( 
.A(n_10494),
.B(n_945),
.Y(n_10848)
);

INVx1_ASAP7_75t_L g10849 ( 
.A(n_10345),
.Y(n_10849)
);

CKINVDCx20_ASAP7_75t_R g10850 ( 
.A(n_10336),
.Y(n_10850)
);

NAND2xp5_ASAP7_75t_L g10851 ( 
.A(n_10385),
.B(n_946),
.Y(n_10851)
);

HB1xp67_ASAP7_75t_L g10852 ( 
.A(n_10270),
.Y(n_10852)
);

HB1xp67_ASAP7_75t_L g10853 ( 
.A(n_10271),
.Y(n_10853)
);

NAND2xp5_ASAP7_75t_L g10854 ( 
.A(n_10399),
.B(n_947),
.Y(n_10854)
);

OA21x2_ASAP7_75t_L g10855 ( 
.A1(n_10348),
.A2(n_947),
.B(n_948),
.Y(n_10855)
);

OAI21xp5_ASAP7_75t_L g10856 ( 
.A1(n_10606),
.A2(n_948),
.B(n_949),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_10354),
.Y(n_10857)
);

INVxp67_ASAP7_75t_L g10858 ( 
.A(n_10589),
.Y(n_10858)
);

OAI21x1_ASAP7_75t_L g10859 ( 
.A1(n_10358),
.A2(n_950),
.B(n_951),
.Y(n_10859)
);

NAND2xp5_ASAP7_75t_L g10860 ( 
.A(n_10410),
.B(n_950),
.Y(n_10860)
);

OAI21x1_ASAP7_75t_L g10861 ( 
.A1(n_10290),
.A2(n_951),
.B(n_952),
.Y(n_10861)
);

AND2x2_ASAP7_75t_L g10862 ( 
.A(n_10282),
.B(n_952),
.Y(n_10862)
);

INVx1_ASAP7_75t_L g10863 ( 
.A(n_10364),
.Y(n_10863)
);

AO31x2_ASAP7_75t_L g10864 ( 
.A1(n_10154),
.A2(n_956),
.A3(n_953),
.B(n_955),
.Y(n_10864)
);

AND2x2_ASAP7_75t_L g10865 ( 
.A(n_10302),
.B(n_953),
.Y(n_10865)
);

OAI21x1_ASAP7_75t_L g10866 ( 
.A1(n_10325),
.A2(n_955),
.B(n_957),
.Y(n_10866)
);

AOI22xp5_ASAP7_75t_L g10867 ( 
.A1(n_10249),
.A2(n_959),
.B1(n_957),
.B2(n_958),
.Y(n_10867)
);

CKINVDCx5p33_ASAP7_75t_R g10868 ( 
.A(n_10285),
.Y(n_10868)
);

OAI21x1_ASAP7_75t_L g10869 ( 
.A1(n_10390),
.A2(n_958),
.B(n_959),
.Y(n_10869)
);

AND2x2_ASAP7_75t_L g10870 ( 
.A(n_10344),
.B(n_960),
.Y(n_10870)
);

OAI22xp33_ASAP7_75t_L g10871 ( 
.A1(n_10228),
.A2(n_962),
.B1(n_960),
.B2(n_961),
.Y(n_10871)
);

NAND2xp5_ASAP7_75t_L g10872 ( 
.A(n_10351),
.B(n_961),
.Y(n_10872)
);

CKINVDCx11_ASAP7_75t_R g10873 ( 
.A(n_10123),
.Y(n_10873)
);

INVx2_ASAP7_75t_L g10874 ( 
.A(n_10356),
.Y(n_10874)
);

OAI21xp5_ASAP7_75t_L g10875 ( 
.A1(n_10340),
.A2(n_962),
.B(n_963),
.Y(n_10875)
);

INVx2_ASAP7_75t_SL g10876 ( 
.A(n_10570),
.Y(n_10876)
);

AO32x2_ASAP7_75t_L g10877 ( 
.A1(n_10037),
.A2(n_966),
.A3(n_964),
.B1(n_965),
.B2(n_967),
.Y(n_10877)
);

NAND2xp5_ASAP7_75t_L g10878 ( 
.A(n_10069),
.B(n_964),
.Y(n_10878)
);

OAI21x1_ASAP7_75t_L g10879 ( 
.A1(n_10395),
.A2(n_965),
.B(n_966),
.Y(n_10879)
);

BUFx10_ASAP7_75t_L g10880 ( 
.A(n_10072),
.Y(n_10880)
);

AOI21xp5_ASAP7_75t_L g10881 ( 
.A1(n_10188),
.A2(n_967),
.B(n_968),
.Y(n_10881)
);

OAI21x1_ASAP7_75t_L g10882 ( 
.A1(n_10398),
.A2(n_969),
.B(n_970),
.Y(n_10882)
);

OAI21xp33_ASAP7_75t_L g10883 ( 
.A1(n_10132),
.A2(n_969),
.B(n_970),
.Y(n_10883)
);

AOI21x1_ASAP7_75t_L g10884 ( 
.A1(n_10148),
.A2(n_971),
.B(n_972),
.Y(n_10884)
);

INVx1_ASAP7_75t_SL g10885 ( 
.A(n_10570),
.Y(n_10885)
);

INVx1_ASAP7_75t_L g10886 ( 
.A(n_10075),
.Y(n_10886)
);

OAI21x1_ASAP7_75t_L g10887 ( 
.A1(n_10409),
.A2(n_971),
.B(n_972),
.Y(n_10887)
);

O2A1O1Ixp5_ASAP7_75t_SL g10888 ( 
.A1(n_10076),
.A2(n_975),
.B(n_973),
.C(n_974),
.Y(n_10888)
);

NOR4xp25_ASAP7_75t_L g10889 ( 
.A(n_10603),
.B(n_977),
.C(n_973),
.D(n_976),
.Y(n_10889)
);

NAND2xp5_ASAP7_75t_L g10890 ( 
.A(n_10088),
.B(n_978),
.Y(n_10890)
);

OAI21x1_ASAP7_75t_L g10891 ( 
.A1(n_10414),
.A2(n_978),
.B(n_979),
.Y(n_10891)
);

BUFx6f_ASAP7_75t_L g10892 ( 
.A(n_10177),
.Y(n_10892)
);

NAND2xp5_ASAP7_75t_L g10893 ( 
.A(n_10104),
.B(n_979),
.Y(n_10893)
);

OAI21x1_ASAP7_75t_L g10894 ( 
.A1(n_10402),
.A2(n_980),
.B(n_981),
.Y(n_10894)
);

AOI21xp5_ASAP7_75t_L g10895 ( 
.A1(n_10108),
.A2(n_980),
.B(n_982),
.Y(n_10895)
);

AND2x4_ASAP7_75t_L g10896 ( 
.A(n_10106),
.B(n_982),
.Y(n_10896)
);

OAI22xp5_ASAP7_75t_L g10897 ( 
.A1(n_10109),
.A2(n_986),
.B1(n_983),
.B2(n_985),
.Y(n_10897)
);

AOI21xp5_ASAP7_75t_L g10898 ( 
.A1(n_10108),
.A2(n_983),
.B(n_986),
.Y(n_10898)
);

A2O1A1Ixp33_ASAP7_75t_L g10899 ( 
.A1(n_10021),
.A2(n_989),
.B(n_987),
.C(n_988),
.Y(n_10899)
);

AOI21xp5_ASAP7_75t_L g10900 ( 
.A1(n_10607),
.A2(n_987),
.B(n_988),
.Y(n_10900)
);

AND2x2_ASAP7_75t_L g10901 ( 
.A(n_10112),
.B(n_989),
.Y(n_10901)
);

NAND2xp5_ASAP7_75t_L g10902 ( 
.A(n_10121),
.B(n_10128),
.Y(n_10902)
);

NOR3xp33_ASAP7_75t_SL g10903 ( 
.A(n_10352),
.B(n_990),
.C(n_991),
.Y(n_10903)
);

AOI21xp33_ASAP7_75t_L g10904 ( 
.A1(n_10374),
.A2(n_992),
.B(n_993),
.Y(n_10904)
);

OAI21x1_ASAP7_75t_L g10905 ( 
.A1(n_10437),
.A2(n_992),
.B(n_994),
.Y(n_10905)
);

NAND2xp5_ASAP7_75t_L g10906 ( 
.A(n_10130),
.B(n_994),
.Y(n_10906)
);

HB1xp67_ASAP7_75t_L g10907 ( 
.A(n_10145),
.Y(n_10907)
);

AO21x1_ASAP7_75t_L g10908 ( 
.A1(n_10569),
.A2(n_995),
.B(n_996),
.Y(n_10908)
);

AND2x4_ASAP7_75t_L g10909 ( 
.A(n_10444),
.B(n_995),
.Y(n_10909)
);

AOI21xp5_ASAP7_75t_L g10910 ( 
.A1(n_10607),
.A2(n_996),
.B(n_997),
.Y(n_10910)
);

INVx1_ASAP7_75t_SL g10911 ( 
.A(n_9999),
.Y(n_10911)
);

OAI21x1_ASAP7_75t_L g10912 ( 
.A1(n_10472),
.A2(n_997),
.B(n_998),
.Y(n_10912)
);

NAND2xp5_ASAP7_75t_L g10913 ( 
.A(n_10593),
.B(n_998),
.Y(n_10913)
);

AO21x2_ASAP7_75t_L g10914 ( 
.A1(n_10624),
.A2(n_9992),
.B(n_10262),
.Y(n_10914)
);

NAND2xp5_ASAP7_75t_L g10915 ( 
.A(n_10596),
.B(n_1000),
.Y(n_10915)
);

OA21x2_ASAP7_75t_L g10916 ( 
.A1(n_10175),
.A2(n_1000),
.B(n_1001),
.Y(n_10916)
);

INVx3_ASAP7_75t_L g10917 ( 
.A(n_10471),
.Y(n_10917)
);

NAND3x1_ASAP7_75t_L g10918 ( 
.A(n_10168),
.B(n_1001),
.C(n_1002),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_10422),
.Y(n_10919)
);

OAI21x1_ASAP7_75t_L g10920 ( 
.A1(n_10481),
.A2(n_1002),
.B(n_1003),
.Y(n_10920)
);

AOI21x1_ASAP7_75t_L g10921 ( 
.A1(n_10101),
.A2(n_10190),
.B(n_10207),
.Y(n_10921)
);

OAI22xp33_ASAP7_75t_L g10922 ( 
.A1(n_10064),
.A2(n_1006),
.B1(n_1004),
.B2(n_1005),
.Y(n_10922)
);

INVx1_ASAP7_75t_L g10923 ( 
.A(n_10445),
.Y(n_10923)
);

NAND2xp5_ASAP7_75t_L g10924 ( 
.A(n_10446),
.B(n_1005),
.Y(n_10924)
);

OA21x2_ASAP7_75t_L g10925 ( 
.A1(n_10215),
.A2(n_1006),
.B(n_1007),
.Y(n_10925)
);

AOI21xp5_ASAP7_75t_L g10926 ( 
.A1(n_10449),
.A2(n_1008),
.B(n_1009),
.Y(n_10926)
);

INVx2_ASAP7_75t_L g10927 ( 
.A(n_10447),
.Y(n_10927)
);

INVx1_ASAP7_75t_L g10928 ( 
.A(n_10450),
.Y(n_10928)
);

AO21x2_ASAP7_75t_L g10929 ( 
.A1(n_10131),
.A2(n_1008),
.B(n_1009),
.Y(n_10929)
);

OAI21x1_ASAP7_75t_L g10930 ( 
.A1(n_10501),
.A2(n_1010),
.B(n_1011),
.Y(n_10930)
);

AND2x2_ASAP7_75t_L g10931 ( 
.A(n_10631),
.B(n_1010),
.Y(n_10931)
);

INVxp67_ASAP7_75t_SL g10932 ( 
.A(n_10451),
.Y(n_10932)
);

AND2x4_ASAP7_75t_L g10933 ( 
.A(n_10489),
.B(n_1011),
.Y(n_10933)
);

AOI21xp33_ASAP7_75t_L g10934 ( 
.A1(n_10407),
.A2(n_1012),
.B(n_1013),
.Y(n_10934)
);

BUFx8_ASAP7_75t_L g10935 ( 
.A(n_10063),
.Y(n_10935)
);

CKINVDCx14_ASAP7_75t_R g10936 ( 
.A(n_10105),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_10510),
.Y(n_10937)
);

NAND3xp33_ASAP7_75t_L g10938 ( 
.A(n_10379),
.B(n_1012),
.C(n_1013),
.Y(n_10938)
);

OAI21xp5_ASAP7_75t_L g10939 ( 
.A1(n_9993),
.A2(n_1014),
.B(n_1015),
.Y(n_10939)
);

AND2x2_ASAP7_75t_L g10940 ( 
.A(n_10316),
.B(n_1014),
.Y(n_10940)
);

NAND3xp33_ASAP7_75t_L g10941 ( 
.A(n_10516),
.B(n_1015),
.C(n_1016),
.Y(n_10941)
);

AOI21xp5_ASAP7_75t_L g10942 ( 
.A1(n_10449),
.A2(n_1017),
.B(n_1018),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_10553),
.B(n_1017),
.Y(n_10943)
);

INVx3_ASAP7_75t_L g10944 ( 
.A(n_10471),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_10555),
.Y(n_10945)
);

AOI22xp5_ASAP7_75t_L g10946 ( 
.A1(n_10053),
.A2(n_1021),
.B1(n_1019),
.B2(n_1020),
.Y(n_10946)
);

A2O1A1Ixp33_ASAP7_75t_L g10947 ( 
.A1(n_10383),
.A2(n_10099),
.B(n_10179),
.C(n_10174),
.Y(n_10947)
);

NAND2xp5_ASAP7_75t_L g10948 ( 
.A(n_10585),
.B(n_1019),
.Y(n_10948)
);

AND2x4_ASAP7_75t_L g10949 ( 
.A(n_10506),
.B(n_1022),
.Y(n_10949)
);

INVx1_ASAP7_75t_L g10950 ( 
.A(n_10512),
.Y(n_10950)
);

NAND2xp5_ASAP7_75t_L g10951 ( 
.A(n_10525),
.B(n_1022),
.Y(n_10951)
);

AOI21xp5_ASAP7_75t_L g10952 ( 
.A1(n_10111),
.A2(n_1023),
.B(n_1024),
.Y(n_10952)
);

OAI21x1_ASAP7_75t_SL g10953 ( 
.A1(n_10392),
.A2(n_1023),
.B(n_1024),
.Y(n_10953)
);

NAND2xp5_ASAP7_75t_L g10954 ( 
.A(n_10533),
.B(n_1025),
.Y(n_10954)
);

AOI21xp5_ASAP7_75t_L g10955 ( 
.A1(n_10216),
.A2(n_1025),
.B(n_1026),
.Y(n_10955)
);

A2O1A1Ixp33_ASAP7_75t_L g10956 ( 
.A1(n_10194),
.A2(n_10208),
.B(n_10220),
.C(n_10202),
.Y(n_10956)
);

BUFx2_ASAP7_75t_L g10957 ( 
.A(n_10405),
.Y(n_10957)
);

AOI21xp5_ASAP7_75t_L g10958 ( 
.A1(n_10308),
.A2(n_1026),
.B(n_1027),
.Y(n_10958)
);

NOR2xp33_ASAP7_75t_L g10959 ( 
.A(n_10084),
.B(n_1027),
.Y(n_10959)
);

INVx1_ASAP7_75t_SL g10960 ( 
.A(n_10150),
.Y(n_10960)
);

INVx2_ASAP7_75t_L g10961 ( 
.A(n_10541),
.Y(n_10961)
);

OAI21x1_ASAP7_75t_L g10962 ( 
.A1(n_10568),
.A2(n_1028),
.B(n_1029),
.Y(n_10962)
);

OAI21x1_ASAP7_75t_L g10963 ( 
.A1(n_10571),
.A2(n_1030),
.B(n_1031),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_10574),
.Y(n_10964)
);

INVx2_ASAP7_75t_SL g10965 ( 
.A(n_10572),
.Y(n_10965)
);

OAI21x1_ASAP7_75t_L g10966 ( 
.A1(n_10575),
.A2(n_1030),
.B(n_1032),
.Y(n_10966)
);

AOI21xp5_ASAP7_75t_L g10967 ( 
.A1(n_10256),
.A2(n_1032),
.B(n_1033),
.Y(n_10967)
);

NOR2x1_ASAP7_75t_L g10968 ( 
.A(n_10181),
.B(n_1033),
.Y(n_10968)
);

INVxp67_ASAP7_75t_L g10969 ( 
.A(n_10382),
.Y(n_10969)
);

AO21x2_ASAP7_75t_L g10970 ( 
.A1(n_10097),
.A2(n_1034),
.B(n_1035),
.Y(n_10970)
);

AOI21xp5_ASAP7_75t_L g10971 ( 
.A1(n_10257),
.A2(n_1034),
.B(n_1035),
.Y(n_10971)
);

BUFx10_ASAP7_75t_L g10972 ( 
.A(n_10496),
.Y(n_10972)
);

BUFx6f_ASAP7_75t_L g10973 ( 
.A(n_10177),
.Y(n_10973)
);

NOR4xp25_ASAP7_75t_L g10974 ( 
.A(n_10458),
.B(n_1038),
.C(n_1036),
.D(n_1037),
.Y(n_10974)
);

AO22x2_ASAP7_75t_L g10975 ( 
.A1(n_10310),
.A2(n_1040),
.B1(n_1036),
.B2(n_1039),
.Y(n_10975)
);

AO31x2_ASAP7_75t_L g10976 ( 
.A1(n_10404),
.A2(n_1041),
.A3(n_1039),
.B(n_1040),
.Y(n_10976)
);

AOI21xp5_ASAP7_75t_L g10977 ( 
.A1(n_10269),
.A2(n_1042),
.B(n_1043),
.Y(n_10977)
);

A2O1A1Ixp33_ASAP7_75t_L g10978 ( 
.A1(n_10234),
.A2(n_1044),
.B(n_1042),
.C(n_1043),
.Y(n_10978)
);

OA21x2_ASAP7_75t_L g10979 ( 
.A1(n_10007),
.A2(n_1044),
.B(n_1045),
.Y(n_10979)
);

OAI21x1_ASAP7_75t_L g10980 ( 
.A1(n_10582),
.A2(n_1045),
.B(n_1046),
.Y(n_10980)
);

AND2x2_ASAP7_75t_L g10981 ( 
.A(n_10028),
.B(n_10078),
.Y(n_10981)
);

OAI21xp5_ASAP7_75t_SL g10982 ( 
.A1(n_10095),
.A2(n_1046),
.B(n_1047),
.Y(n_10982)
);

AND2x2_ASAP7_75t_L g10983 ( 
.A(n_10085),
.B(n_1047),
.Y(n_10983)
);

AO32x2_ASAP7_75t_L g10984 ( 
.A1(n_10087),
.A2(n_1050),
.A3(n_1048),
.B1(n_1049),
.B2(n_1051),
.Y(n_10984)
);

NAND3x1_ASAP7_75t_L g10985 ( 
.A(n_10082),
.B(n_1048),
.C(n_1049),
.Y(n_10985)
);

OAI21xp5_ASAP7_75t_L g10986 ( 
.A1(n_10138),
.A2(n_1050),
.B(n_1052),
.Y(n_10986)
);

AOI21xp5_ASAP7_75t_L g10987 ( 
.A1(n_10254),
.A2(n_1052),
.B(n_1053),
.Y(n_10987)
);

AOI21xp5_ASAP7_75t_L g10988 ( 
.A1(n_10107),
.A2(n_1053),
.B(n_1054),
.Y(n_10988)
);

BUFx2_ASAP7_75t_L g10989 ( 
.A(n_10405),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_10584),
.Y(n_10990)
);

AO31x2_ASAP7_75t_L g10991 ( 
.A1(n_10326),
.A2(n_1056),
.A3(n_1054),
.B(n_1055),
.Y(n_10991)
);

AOI21xp5_ASAP7_75t_L g10992 ( 
.A1(n_10495),
.A2(n_1055),
.B(n_1056),
.Y(n_10992)
);

AND2x2_ASAP7_75t_L g10993 ( 
.A(n_10018),
.B(n_1057),
.Y(n_10993)
);

AOI21xp5_ASAP7_75t_L g10994 ( 
.A1(n_10278),
.A2(n_1057),
.B(n_1058),
.Y(n_10994)
);

OAI21x1_ASAP7_75t_L g10995 ( 
.A1(n_10433),
.A2(n_1058),
.B(n_1059),
.Y(n_10995)
);

NOR4xp25_ASAP7_75t_L g10996 ( 
.A(n_10039),
.B(n_1061),
.C(n_1059),
.D(n_1060),
.Y(n_10996)
);

NAND3xp33_ASAP7_75t_SL g10997 ( 
.A(n_10573),
.B(n_1060),
.C(n_1061),
.Y(n_10997)
);

INVx2_ASAP7_75t_SL g10998 ( 
.A(n_10572),
.Y(n_10998)
);

OAI21x1_ASAP7_75t_L g10999 ( 
.A1(n_10448),
.A2(n_1062),
.B(n_1063),
.Y(n_10999)
);

AOI221x1_ASAP7_75t_L g11000 ( 
.A1(n_10613),
.A2(n_1064),
.B1(n_1062),
.B2(n_1063),
.C(n_1065),
.Y(n_11000)
);

NAND3xp33_ASAP7_75t_L g11001 ( 
.A(n_10321),
.B(n_1064),
.C(n_1065),
.Y(n_11001)
);

INVx1_ASAP7_75t_SL g11002 ( 
.A(n_10176),
.Y(n_11002)
);

OAI21xp5_ASAP7_75t_L g11003 ( 
.A1(n_10315),
.A2(n_1066),
.B(n_1067),
.Y(n_11003)
);

AOI211x1_ASAP7_75t_L g11004 ( 
.A1(n_10330),
.A2(n_1068),
.B(n_1066),
.C(n_1067),
.Y(n_11004)
);

NAND2xp5_ASAP7_75t_L g11005 ( 
.A(n_10031),
.B(n_1068),
.Y(n_11005)
);

CKINVDCx20_ASAP7_75t_R g11006 ( 
.A(n_10619),
.Y(n_11006)
);

NAND2xp5_ASAP7_75t_L g11007 ( 
.A(n_10165),
.B(n_1069),
.Y(n_11007)
);

NAND2xp5_ASAP7_75t_L g11008 ( 
.A(n_10331),
.B(n_1070),
.Y(n_11008)
);

AOI21xp5_ASAP7_75t_L g11009 ( 
.A1(n_10306),
.A2(n_1070),
.B(n_1072),
.Y(n_11009)
);

O2A1O1Ixp33_ASAP7_75t_L g11010 ( 
.A1(n_10314),
.A2(n_1075),
.B(n_1073),
.C(n_1074),
.Y(n_11010)
);

NAND2xp5_ASAP7_75t_L g11011 ( 
.A(n_10246),
.B(n_1073),
.Y(n_11011)
);

NAND2xp5_ASAP7_75t_L g11012 ( 
.A(n_10000),
.B(n_1074),
.Y(n_11012)
);

INVx2_ASAP7_75t_L g11013 ( 
.A(n_10363),
.Y(n_11013)
);

NAND2xp5_ASAP7_75t_L g11014 ( 
.A(n_10156),
.B(n_1075),
.Y(n_11014)
);

OAI21xp5_ASAP7_75t_L g11015 ( 
.A1(n_10126),
.A2(n_1076),
.B(n_1077),
.Y(n_11015)
);

INVx6_ASAP7_75t_L g11016 ( 
.A(n_10318),
.Y(n_11016)
);

NAND2xp5_ASAP7_75t_L g11017 ( 
.A(n_10201),
.B(n_1076),
.Y(n_11017)
);

NAND2xp5_ASAP7_75t_SL g11018 ( 
.A(n_10507),
.B(n_1078),
.Y(n_11018)
);

OAI21x1_ASAP7_75t_L g11019 ( 
.A1(n_10463),
.A2(n_1078),
.B(n_1079),
.Y(n_11019)
);

BUFx6f_ASAP7_75t_L g11020 ( 
.A(n_10204),
.Y(n_11020)
);

OAI21x1_ASAP7_75t_L g11021 ( 
.A1(n_10470),
.A2(n_1079),
.B(n_1080),
.Y(n_11021)
);

OAI21xp5_ASAP7_75t_L g11022 ( 
.A1(n_10499),
.A2(n_1081),
.B(n_1082),
.Y(n_11022)
);

HB1xp67_ASAP7_75t_L g11023 ( 
.A(n_10423),
.Y(n_11023)
);

BUFx2_ASAP7_75t_L g11024 ( 
.A(n_10277),
.Y(n_11024)
);

AOI21xp33_ASAP7_75t_L g11025 ( 
.A1(n_10475),
.A2(n_1081),
.B(n_1083),
.Y(n_11025)
);

A2O1A1Ixp33_ASAP7_75t_L g11026 ( 
.A1(n_10376),
.A2(n_1085),
.B(n_1083),
.C(n_1084),
.Y(n_11026)
);

INVx1_ASAP7_75t_L g11027 ( 
.A(n_10474),
.Y(n_11027)
);

O2A1O1Ixp5_ASAP7_75t_L g11028 ( 
.A1(n_10119),
.A2(n_1086),
.B(n_1084),
.C(n_1085),
.Y(n_11028)
);

AOI21xp5_ASAP7_75t_L g11029 ( 
.A1(n_10193),
.A2(n_10058),
.B(n_10419),
.Y(n_11029)
);

OAI21x1_ASAP7_75t_L g11030 ( 
.A1(n_10478),
.A2(n_1087),
.B(n_1088),
.Y(n_11030)
);

INVx2_ASAP7_75t_L g11031 ( 
.A(n_10480),
.Y(n_11031)
);

AND2x2_ASAP7_75t_L g11032 ( 
.A(n_10476),
.B(n_10266),
.Y(n_11032)
);

OAI21xp5_ASAP7_75t_L g11033 ( 
.A1(n_10522),
.A2(n_1087),
.B(n_1089),
.Y(n_11033)
);

INVx5_ASAP7_75t_L g11034 ( 
.A(n_10052),
.Y(n_11034)
);

AOI22xp33_ASAP7_75t_L g11035 ( 
.A1(n_10094),
.A2(n_1092),
.B1(n_1090),
.B2(n_1091),
.Y(n_11035)
);

INVx2_ASAP7_75t_L g11036 ( 
.A(n_10502),
.Y(n_11036)
);

AOI21xp5_ASAP7_75t_L g11037 ( 
.A1(n_10058),
.A2(n_1090),
.B(n_1092),
.Y(n_11037)
);

OR2x2_ASAP7_75t_L g11038 ( 
.A(n_10113),
.B(n_1093),
.Y(n_11038)
);

BUFx2_ASAP7_75t_L g11039 ( 
.A(n_10089),
.Y(n_11039)
);

OAI21xp5_ASAP7_75t_L g11040 ( 
.A1(n_10539),
.A2(n_1093),
.B(n_1094),
.Y(n_11040)
);

OAI22xp33_ASAP7_75t_L g11041 ( 
.A1(n_10565),
.A2(n_1096),
.B1(n_1094),
.B2(n_1095),
.Y(n_11041)
);

AOI21xp5_ASAP7_75t_L g11042 ( 
.A1(n_10625),
.A2(n_1096),
.B(n_1097),
.Y(n_11042)
);

NOR2xp33_ASAP7_75t_L g11043 ( 
.A(n_10185),
.B(n_1098),
.Y(n_11043)
);

BUFx12f_ASAP7_75t_L g11044 ( 
.A(n_10523),
.Y(n_11044)
);

AO21x1_ASAP7_75t_L g11045 ( 
.A1(n_10527),
.A2(n_10056),
.B(n_10023),
.Y(n_11045)
);

NAND2xp5_ASAP7_75t_L g11046 ( 
.A(n_10116),
.B(n_1098),
.Y(n_11046)
);

NAND2xp5_ASAP7_75t_L g11047 ( 
.A(n_10117),
.B(n_1099),
.Y(n_11047)
);

NAND2xp5_ASAP7_75t_L g11048 ( 
.A(n_10066),
.B(n_1099),
.Y(n_11048)
);

AOI21xp5_ASAP7_75t_L g11049 ( 
.A1(n_10632),
.A2(n_1100),
.B(n_1101),
.Y(n_11049)
);

NAND2xp5_ASAP7_75t_L g11050 ( 
.A(n_10090),
.B(n_1101),
.Y(n_11050)
);

OAI21xp33_ASAP7_75t_L g11051 ( 
.A1(n_10002),
.A2(n_1102),
.B(n_1103),
.Y(n_11051)
);

NAND2xp5_ASAP7_75t_L g11052 ( 
.A(n_10292),
.B(n_10347),
.Y(n_11052)
);

OAI22xp5_ASAP7_75t_L g11053 ( 
.A1(n_10520),
.A2(n_1106),
.B1(n_1104),
.B2(n_1105),
.Y(n_11053)
);

OAI21x1_ASAP7_75t_L g11054 ( 
.A1(n_10511),
.A2(n_1104),
.B(n_1106),
.Y(n_11054)
);

OA21x2_ASAP7_75t_L g11055 ( 
.A1(n_10519),
.A2(n_10536),
.B(n_10521),
.Y(n_11055)
);

INVx1_ASAP7_75t_SL g11056 ( 
.A(n_10460),
.Y(n_11056)
);

AND2x4_ASAP7_75t_L g11057 ( 
.A(n_9996),
.B(n_1107),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10543),
.Y(n_11058)
);

BUFx2_ASAP7_75t_L g11059 ( 
.A(n_10260),
.Y(n_11059)
);

BUFx3_ASAP7_75t_L g11060 ( 
.A(n_10604),
.Y(n_11060)
);

AOI221xp5_ASAP7_75t_L g11061 ( 
.A1(n_10577),
.A2(n_1110),
.B1(n_1108),
.B2(n_1109),
.C(n_1111),
.Y(n_11061)
);

AO21x2_ASAP7_75t_L g11062 ( 
.A1(n_10547),
.A2(n_10554),
.B(n_10551),
.Y(n_11062)
);

INVx1_ASAP7_75t_L g11063 ( 
.A(n_10586),
.Y(n_11063)
);

AO22x2_ASAP7_75t_L g11064 ( 
.A1(n_10203),
.A2(n_1111),
.B1(n_1108),
.B2(n_1109),
.Y(n_11064)
);

AO21x1_ASAP7_75t_L g11065 ( 
.A1(n_10350),
.A2(n_1112),
.B(n_1113),
.Y(n_11065)
);

AO31x2_ASAP7_75t_L g11066 ( 
.A1(n_10250),
.A2(n_1114),
.A3(n_1112),
.B(n_1113),
.Y(n_11066)
);

NOR2xp33_ASAP7_75t_SL g11067 ( 
.A(n_10324),
.B(n_1114),
.Y(n_11067)
);

A2O1A1Ixp33_ASAP7_75t_L g11068 ( 
.A1(n_10560),
.A2(n_1117),
.B(n_1115),
.C(n_1116),
.Y(n_11068)
);

OAI21x1_ASAP7_75t_L g11069 ( 
.A1(n_10467),
.A2(n_1115),
.B(n_1118),
.Y(n_11069)
);

AOI21xp5_ASAP7_75t_L g11070 ( 
.A1(n_10617),
.A2(n_1118),
.B(n_1119),
.Y(n_11070)
);

OAI21xp5_ASAP7_75t_L g11071 ( 
.A1(n_10578),
.A2(n_1119),
.B(n_1120),
.Y(n_11071)
);

OAI21x1_ASAP7_75t_L g11072 ( 
.A1(n_10040),
.A2(n_1121),
.B(n_1122),
.Y(n_11072)
);

OAI21x1_ASAP7_75t_SL g11073 ( 
.A1(n_10319),
.A2(n_1121),
.B(n_1123),
.Y(n_11073)
);

AOI21xp5_ASAP7_75t_SL g11074 ( 
.A1(n_10492),
.A2(n_1123),
.B(n_1124),
.Y(n_11074)
);

AO22x2_ASAP7_75t_L g11075 ( 
.A1(n_10192),
.A2(n_1126),
.B1(n_1124),
.B2(n_1125),
.Y(n_11075)
);

NAND2xp5_ASAP7_75t_SL g11076 ( 
.A(n_10620),
.B(n_1126),
.Y(n_11076)
);

INVx1_ASAP7_75t_L g11077 ( 
.A(n_10059),
.Y(n_11077)
);

OAI22xp5_ASAP7_75t_L g11078 ( 
.A1(n_10498),
.A2(n_1129),
.B1(n_1127),
.B2(n_1128),
.Y(n_11078)
);

NOR2x1_ASAP7_75t_R g11079 ( 
.A(n_10252),
.B(n_1128),
.Y(n_11079)
);

A2O1A1Ixp33_ASAP7_75t_L g11080 ( 
.A1(n_10595),
.A2(n_1132),
.B(n_1129),
.C(n_1131),
.Y(n_11080)
);

OAI22xp5_ASAP7_75t_L g11081 ( 
.A1(n_10081),
.A2(n_10052),
.B1(n_10195),
.B2(n_10164),
.Y(n_11081)
);

INVx1_ASAP7_75t_L g11082 ( 
.A(n_10219),
.Y(n_11082)
);

NAND2xp5_ASAP7_75t_L g11083 ( 
.A(n_10284),
.B(n_1131),
.Y(n_11083)
);

AO31x2_ASAP7_75t_L g11084 ( 
.A1(n_10434),
.A2(n_10454),
.A3(n_10429),
.B(n_10153),
.Y(n_11084)
);

OAI21xp5_ASAP7_75t_L g11085 ( 
.A1(n_10482),
.A2(n_1132),
.B(n_1133),
.Y(n_11085)
);

OA21x2_ASAP7_75t_L g11086 ( 
.A1(n_10197),
.A2(n_1134),
.B(n_1135),
.Y(n_11086)
);

OAI21xp5_ASAP7_75t_L g11087 ( 
.A1(n_10488),
.A2(n_1134),
.B(n_1135),
.Y(n_11087)
);

OAI21xp5_ASAP7_75t_L g11088 ( 
.A1(n_10514),
.A2(n_1136),
.B(n_1137),
.Y(n_11088)
);

CKINVDCx16_ASAP7_75t_R g11089 ( 
.A(n_10477),
.Y(n_11089)
);

INVx1_ASAP7_75t_L g11090 ( 
.A(n_10294),
.Y(n_11090)
);

AOI21xp5_ASAP7_75t_L g11091 ( 
.A1(n_10629),
.A2(n_1136),
.B(n_1137),
.Y(n_11091)
);

NOR2xp33_ASAP7_75t_R g11092 ( 
.A(n_10086),
.B(n_1138),
.Y(n_11092)
);

NAND3x1_ASAP7_75t_L g11093 ( 
.A(n_10167),
.B(n_1138),
.C(n_1139),
.Y(n_11093)
);

NAND2xp5_ASAP7_75t_L g11094 ( 
.A(n_10296),
.B(n_1139),
.Y(n_11094)
);

NOR2x1_ASAP7_75t_L g11095 ( 
.A(n_10338),
.B(n_1140),
.Y(n_11095)
);

INVx2_ASAP7_75t_L g11096 ( 
.A(n_10346),
.Y(n_11096)
);

OR2x2_ASAP7_75t_L g11097 ( 
.A(n_10274),
.B(n_1140),
.Y(n_11097)
);

OAI21xp5_ASAP7_75t_L g11098 ( 
.A1(n_10513),
.A2(n_1141),
.B(n_1142),
.Y(n_11098)
);

A2O1A1Ixp33_ASAP7_75t_L g11099 ( 
.A1(n_10484),
.A2(n_1144),
.B(n_1142),
.C(n_1143),
.Y(n_11099)
);

OAI22x1_ASAP7_75t_L g11100 ( 
.A1(n_10562),
.A2(n_10065),
.B1(n_10127),
.B2(n_10182),
.Y(n_11100)
);

OAI21x1_ASAP7_75t_L g11101 ( 
.A1(n_10323),
.A2(n_1143),
.B(n_1144),
.Y(n_11101)
);

AOI21xp5_ASAP7_75t_L g11102 ( 
.A1(n_10456),
.A2(n_1145),
.B(n_1146),
.Y(n_11102)
);

OAI21x1_ASAP7_75t_L g11103 ( 
.A1(n_10222),
.A2(n_1145),
.B(n_1146),
.Y(n_11103)
);

OAI22xp5_ASAP7_75t_L g11104 ( 
.A1(n_10411),
.A2(n_1149),
.B1(n_1147),
.B2(n_1148),
.Y(n_11104)
);

AOI21xp5_ASAP7_75t_SL g11105 ( 
.A1(n_10503),
.A2(n_10518),
.B(n_10515),
.Y(n_11105)
);

A2O1A1Ixp33_ASAP7_75t_L g11106 ( 
.A1(n_10483),
.A2(n_1149),
.B(n_1147),
.C(n_1148),
.Y(n_11106)
);

INVx3_ASAP7_75t_L g11107 ( 
.A(n_10517),
.Y(n_11107)
);

AO21x1_ASAP7_75t_L g11108 ( 
.A1(n_10311),
.A2(n_1150),
.B(n_1151),
.Y(n_11108)
);

AO31x2_ASAP7_75t_L g11109 ( 
.A1(n_10287),
.A2(n_1153),
.A3(n_1151),
.B(n_1152),
.Y(n_11109)
);

OAI21x1_ASAP7_75t_L g11110 ( 
.A1(n_10226),
.A2(n_1152),
.B(n_1153),
.Y(n_11110)
);

NOR2xp67_ASAP7_75t_SL g11111 ( 
.A(n_10212),
.B(n_1154),
.Y(n_11111)
);

AOI21xp5_ASAP7_75t_L g11112 ( 
.A1(n_10349),
.A2(n_1154),
.B(n_1156),
.Y(n_11112)
);

NAND2xp5_ASAP7_75t_L g11113 ( 
.A(n_10591),
.B(n_1156),
.Y(n_11113)
);

NAND2xp5_ASAP7_75t_SL g11114 ( 
.A(n_10487),
.B(n_1157),
.Y(n_11114)
);

OR2x6_ASAP7_75t_L g11115 ( 
.A(n_10396),
.B(n_1157),
.Y(n_11115)
);

NAND3xp33_ASAP7_75t_L g11116 ( 
.A(n_10233),
.B(n_10251),
.C(n_10630),
.Y(n_11116)
);

AOI21x1_ASAP7_75t_SL g11117 ( 
.A1(n_10627),
.A2(n_1158),
.B(n_1159),
.Y(n_11117)
);

OAI21x1_ASAP7_75t_L g11118 ( 
.A1(n_10241),
.A2(n_1159),
.B(n_1160),
.Y(n_11118)
);

NAND2xp5_ASAP7_75t_L g11119 ( 
.A(n_10592),
.B(n_1160),
.Y(n_11119)
);

CKINVDCx20_ASAP7_75t_R g11120 ( 
.A(n_10401),
.Y(n_11120)
);

INVx1_ASAP7_75t_L g11121 ( 
.A(n_10342),
.Y(n_11121)
);

NAND2xp5_ASAP7_75t_L g11122 ( 
.A(n_10612),
.B(n_1161),
.Y(n_11122)
);

AOI21xp5_ASAP7_75t_L g11123 ( 
.A1(n_10601),
.A2(n_10561),
.B(n_10544),
.Y(n_11123)
);

OAI21x1_ASAP7_75t_L g11124 ( 
.A1(n_10362),
.A2(n_1161),
.B(n_1162),
.Y(n_11124)
);

NAND2xp5_ASAP7_75t_SL g11125 ( 
.A(n_10487),
.B(n_1162),
.Y(n_11125)
);

NAND2xp5_ASAP7_75t_SL g11126 ( 
.A(n_10050),
.B(n_1163),
.Y(n_11126)
);

CKINVDCx5p33_ASAP7_75t_R g11127 ( 
.A(n_10036),
.Y(n_11127)
);

INVx1_ASAP7_75t_L g11128 ( 
.A(n_10367),
.Y(n_11128)
);

NAND2xp5_ASAP7_75t_L g11129 ( 
.A(n_10618),
.B(n_1164),
.Y(n_11129)
);

INVx2_ASAP7_75t_L g11130 ( 
.A(n_10517),
.Y(n_11130)
);

INVx1_ASAP7_75t_L g11131 ( 
.A(n_10806),
.Y(n_11131)
);

INVx2_ASAP7_75t_SL g11132 ( 
.A(n_10781),
.Y(n_11132)
);

INVx2_ASAP7_75t_L g11133 ( 
.A(n_10773),
.Y(n_11133)
);

INVx3_ASAP7_75t_L g11134 ( 
.A(n_10714),
.Y(n_11134)
);

NAND2x1p5_ASAP7_75t_L g11135 ( 
.A(n_11034),
.B(n_10745),
.Y(n_11135)
);

CKINVDCx5p33_ASAP7_75t_R g11136 ( 
.A(n_10760),
.Y(n_11136)
);

INVx1_ASAP7_75t_L g11137 ( 
.A(n_10777),
.Y(n_11137)
);

INVx3_ASAP7_75t_L g11138 ( 
.A(n_10780),
.Y(n_11138)
);

NAND2xp5_ASAP7_75t_L g11139 ( 
.A(n_10639),
.B(n_10110),
.Y(n_11139)
);

INVx1_ASAP7_75t_L g11140 ( 
.A(n_10652),
.Y(n_11140)
);

INVx1_ASAP7_75t_SL g11141 ( 
.A(n_10815),
.Y(n_11141)
);

NAND2xp5_ASAP7_75t_L g11142 ( 
.A(n_10858),
.B(n_10071),
.Y(n_11142)
);

NAND2xp5_ASAP7_75t_L g11143 ( 
.A(n_10637),
.B(n_10025),
.Y(n_11143)
);

AND2x2_ASAP7_75t_L g11144 ( 
.A(n_10743),
.B(n_10377),
.Y(n_11144)
);

A2O1A1Ixp33_ASAP7_75t_L g11145 ( 
.A1(n_10752),
.A2(n_10057),
.B(n_10061),
.C(n_10621),
.Y(n_11145)
);

AOI21xp5_ASAP7_75t_L g11146 ( 
.A1(n_10785),
.A2(n_10761),
.B(n_10664),
.Y(n_11146)
);

INVxp67_ASAP7_75t_L g11147 ( 
.A(n_11023),
.Y(n_11147)
);

BUFx6f_ASAP7_75t_L g11148 ( 
.A(n_10661),
.Y(n_11148)
);

INVx2_ASAP7_75t_L g11149 ( 
.A(n_10654),
.Y(n_11149)
);

INVx1_ASAP7_75t_L g11150 ( 
.A(n_10657),
.Y(n_11150)
);

NAND2xp33_ASAP7_75t_L g11151 ( 
.A(n_10784),
.B(n_10559),
.Y(n_11151)
);

OR2x2_ASAP7_75t_SL g11152 ( 
.A(n_11089),
.B(n_10599),
.Y(n_11152)
);

AOI211xp5_ASAP7_75t_L g11153 ( 
.A1(n_10669),
.A2(n_10298),
.B(n_10465),
.C(n_10333),
.Y(n_11153)
);

INVx2_ASAP7_75t_L g11154 ( 
.A(n_10660),
.Y(n_11154)
);

INVx1_ASAP7_75t_L g11155 ( 
.A(n_10696),
.Y(n_11155)
);

NAND2xp5_ASAP7_75t_L g11156 ( 
.A(n_10798),
.B(n_10646),
.Y(n_11156)
);

HB1xp67_ASAP7_75t_L g11157 ( 
.A(n_10852),
.Y(n_11157)
);

OAI21xp33_ASAP7_75t_L g11158 ( 
.A1(n_10754),
.A2(n_10490),
.B(n_10417),
.Y(n_11158)
);

BUFx2_ASAP7_75t_L g11159 ( 
.A(n_10769),
.Y(n_11159)
);

BUFx6f_ASAP7_75t_L g11160 ( 
.A(n_10666),
.Y(n_11160)
);

NOR2x1_ASAP7_75t_SL g11161 ( 
.A(n_10676),
.B(n_10412),
.Y(n_11161)
);

NAND2xp5_ASAP7_75t_SL g11162 ( 
.A(n_11034),
.B(n_10530),
.Y(n_11162)
);

OR2x2_ASAP7_75t_L g11163 ( 
.A(n_10649),
.B(n_10280),
.Y(n_11163)
);

NAND2xp5_ASAP7_75t_L g11164 ( 
.A(n_10755),
.B(n_10045),
.Y(n_11164)
);

INVx2_ASAP7_75t_L g11165 ( 
.A(n_10701),
.Y(n_11165)
);

INVx1_ASAP7_75t_L g11166 ( 
.A(n_10710),
.Y(n_11166)
);

NAND2xp5_ASAP7_75t_L g11167 ( 
.A(n_10651),
.B(n_10049),
.Y(n_11167)
);

AOI21xp5_ASAP7_75t_L g11168 ( 
.A1(n_10829),
.A2(n_10427),
.B(n_10403),
.Y(n_11168)
);

AOI222xp33_ASAP7_75t_L g11169 ( 
.A1(n_10716),
.A2(n_10615),
.B1(n_10581),
.B2(n_10605),
.C1(n_10588),
.C2(n_10611),
.Y(n_11169)
);

INVxp67_ASAP7_75t_L g11170 ( 
.A(n_10703),
.Y(n_11170)
);

NAND2x1p5_ASAP7_75t_L g11171 ( 
.A(n_10671),
.B(n_10550),
.Y(n_11171)
);

INVx2_ASAP7_75t_L g11172 ( 
.A(n_10729),
.Y(n_11172)
);

INVx1_ASAP7_75t_L g11173 ( 
.A(n_10736),
.Y(n_11173)
);

INVx1_ASAP7_75t_L g11174 ( 
.A(n_10751),
.Y(n_11174)
);

NOR2xp33_ASAP7_75t_L g11175 ( 
.A(n_10957),
.B(n_10989),
.Y(n_11175)
);

BUFx2_ASAP7_75t_L g11176 ( 
.A(n_10768),
.Y(n_11176)
);

BUFx12f_ASAP7_75t_L g11177 ( 
.A(n_10935),
.Y(n_11177)
);

AOI21xp5_ASAP7_75t_L g11178 ( 
.A1(n_10956),
.A2(n_10741),
.B(n_10706),
.Y(n_11178)
);

AND2x2_ASAP7_75t_SL g11179 ( 
.A(n_10889),
.B(n_10549),
.Y(n_11179)
);

INVxp67_ASAP7_75t_L g11180 ( 
.A(n_11121),
.Y(n_11180)
);

INVx2_ASAP7_75t_L g11181 ( 
.A(n_10766),
.Y(n_11181)
);

AND2x4_ASAP7_75t_L g11182 ( 
.A(n_10719),
.B(n_10365),
.Y(n_11182)
);

BUFx2_ASAP7_75t_L g11183 ( 
.A(n_11039),
.Y(n_11183)
);

AOI21xp5_ASAP7_75t_L g11184 ( 
.A1(n_10735),
.A2(n_10485),
.B(n_10442),
.Y(n_11184)
);

INVx1_ASAP7_75t_L g11185 ( 
.A(n_10810),
.Y(n_11185)
);

NAND2xp5_ASAP7_75t_L g11186 ( 
.A(n_11036),
.B(n_10508),
.Y(n_11186)
);

AND2x4_ASAP7_75t_L g11187 ( 
.A(n_11059),
.B(n_10373),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_10834),
.Y(n_11188)
);

INVx1_ASAP7_75t_SL g11189 ( 
.A(n_10744),
.Y(n_11189)
);

AND2x4_ASAP7_75t_L g11190 ( 
.A(n_11031),
.B(n_11096),
.Y(n_11190)
);

BUFx3_ASAP7_75t_L g11191 ( 
.A(n_10784),
.Y(n_11191)
);

INVx6_ASAP7_75t_SL g11192 ( 
.A(n_10972),
.Y(n_11192)
);

INVx2_ASAP7_75t_L g11193 ( 
.A(n_10842),
.Y(n_11193)
);

BUFx2_ASAP7_75t_L g11194 ( 
.A(n_10853),
.Y(n_11194)
);

AOI21xp5_ASAP7_75t_L g11195 ( 
.A1(n_10739),
.A2(n_10493),
.B(n_10491),
.Y(n_11195)
);

BUFx2_ASAP7_75t_R g11196 ( 
.A(n_10633),
.Y(n_11196)
);

INVx1_ASAP7_75t_L g11197 ( 
.A(n_10849),
.Y(n_11197)
);

INVx2_ASAP7_75t_L g11198 ( 
.A(n_10857),
.Y(n_11198)
);

AND2x4_ASAP7_75t_L g11199 ( 
.A(n_10932),
.B(n_10397),
.Y(n_11199)
);

INVx1_ASAP7_75t_L g11200 ( 
.A(n_10863),
.Y(n_11200)
);

OAI21x1_ASAP7_75t_L g11201 ( 
.A1(n_10663),
.A2(n_10635),
.B(n_10833),
.Y(n_11201)
);

BUFx2_ASAP7_75t_L g11202 ( 
.A(n_10907),
.Y(n_11202)
);

AOI21xp5_ASAP7_75t_L g11203 ( 
.A1(n_10642),
.A2(n_10524),
.B(n_10387),
.Y(n_11203)
);

OAI22xp5_ASAP7_75t_L g11204 ( 
.A1(n_11001),
.A2(n_10396),
.B1(n_10412),
.B2(n_10142),
.Y(n_11204)
);

AND2x4_ASAP7_75t_L g11205 ( 
.A(n_10927),
.B(n_10622),
.Y(n_11205)
);

INVx2_ASAP7_75t_L g11206 ( 
.A(n_10919),
.Y(n_11206)
);

AND2x4_ASAP7_75t_L g11207 ( 
.A(n_10886),
.B(n_10229),
.Y(n_11207)
);

INVx1_ASAP7_75t_L g11208 ( 
.A(n_10923),
.Y(n_11208)
);

INVx3_ASAP7_75t_L g11209 ( 
.A(n_10678),
.Y(n_11209)
);

CKINVDCx5p33_ASAP7_75t_R g11210 ( 
.A(n_10641),
.Y(n_11210)
);

NOR2xp33_ASAP7_75t_R g11211 ( 
.A(n_11006),
.B(n_10259),
.Y(n_11211)
);

AOI21xp5_ASAP7_75t_L g11212 ( 
.A1(n_10636),
.A2(n_10841),
.B(n_10811),
.Y(n_11212)
);

NAND2xp5_ASAP7_75t_L g11213 ( 
.A(n_11027),
.B(n_10217),
.Y(n_11213)
);

NOR2xp33_ASAP7_75t_L g11214 ( 
.A(n_10644),
.B(n_10604),
.Y(n_11214)
);

BUFx6f_ASAP7_75t_L g11215 ( 
.A(n_10655),
.Y(n_11215)
);

INVx1_ASAP7_75t_SL g11216 ( 
.A(n_10873),
.Y(n_11216)
);

AOI21x1_ASAP7_75t_L g11217 ( 
.A1(n_11100),
.A2(n_10129),
.B(n_10389),
.Y(n_11217)
);

INVx1_ASAP7_75t_L g11218 ( 
.A(n_10928),
.Y(n_11218)
);

INVx2_ASAP7_75t_L g11219 ( 
.A(n_10634),
.Y(n_11219)
);

INVx2_ASAP7_75t_L g11220 ( 
.A(n_10722),
.Y(n_11220)
);

INVx3_ASAP7_75t_L g11221 ( 
.A(n_10787),
.Y(n_11221)
);

AOI22xp5_ASAP7_75t_L g11222 ( 
.A1(n_10847),
.A2(n_10759),
.B1(n_10789),
.B2(n_10883),
.Y(n_11222)
);

OA21x2_ASAP7_75t_L g11223 ( 
.A1(n_10832),
.A2(n_10416),
.B(n_10309),
.Y(n_11223)
);

AOI21xp5_ASAP7_75t_L g11224 ( 
.A1(n_10904),
.A2(n_10609),
.B(n_10546),
.Y(n_11224)
);

OAI31xp33_ASAP7_75t_L g11225 ( 
.A1(n_10693),
.A2(n_10359),
.A3(n_10421),
.B(n_10628),
.Y(n_11225)
);

BUFx3_ASAP7_75t_L g11226 ( 
.A(n_10838),
.Y(n_11226)
);

BUFx3_ASAP7_75t_L g11227 ( 
.A(n_11044),
.Y(n_11227)
);

AOI21xp5_ASAP7_75t_L g11228 ( 
.A1(n_10797),
.A2(n_10264),
.B(n_10243),
.Y(n_11228)
);

BUFx6f_ASAP7_75t_L g11229 ( 
.A(n_10655),
.Y(n_11229)
);

AOI21xp5_ASAP7_75t_L g11230 ( 
.A1(n_10779),
.A2(n_10455),
.B(n_10532),
.Y(n_11230)
);

NAND2xp5_ASAP7_75t_L g11231 ( 
.A(n_11058),
.B(n_10291),
.Y(n_11231)
);

NAND2xp5_ASAP7_75t_L g11232 ( 
.A(n_11063),
.B(n_10328),
.Y(n_11232)
);

AND2x4_ASAP7_75t_L g11233 ( 
.A(n_10950),
.B(n_10060),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_10937),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_10945),
.Y(n_11235)
);

AOI21xp5_ASAP7_75t_L g11236 ( 
.A1(n_10947),
.A2(n_10169),
.B(n_10526),
.Y(n_11236)
);

NAND2xp5_ASAP7_75t_L g11237 ( 
.A(n_11055),
.B(n_10370),
.Y(n_11237)
);

OAI22xp5_ASAP7_75t_L g11238 ( 
.A1(n_11026),
.A2(n_10210),
.B1(n_10297),
.B2(n_10183),
.Y(n_11238)
);

NOR2xp33_ASAP7_75t_L g11239 ( 
.A(n_10969),
.B(n_10616),
.Y(n_11239)
);

INVx1_ASAP7_75t_L g11240 ( 
.A(n_10770),
.Y(n_11240)
);

AND2x4_ASAP7_75t_L g11241 ( 
.A(n_10964),
.B(n_10388),
.Y(n_11241)
);

OAI22xp5_ASAP7_75t_L g11242 ( 
.A1(n_11116),
.A2(n_10430),
.B1(n_10616),
.B2(n_10272),
.Y(n_11242)
);

AOI21xp5_ASAP7_75t_L g11243 ( 
.A1(n_10687),
.A2(n_10799),
.B(n_11009),
.Y(n_11243)
);

NAND2xp5_ASAP7_75t_L g11244 ( 
.A(n_11077),
.B(n_10443),
.Y(n_11244)
);

BUFx12f_ASAP7_75t_L g11245 ( 
.A(n_10724),
.Y(n_11245)
);

AO32x1_ASAP7_75t_L g11246 ( 
.A1(n_11053),
.A2(n_10439),
.A3(n_10548),
.B1(n_10608),
.B2(n_10468),
.Y(n_11246)
);

BUFx2_ASAP7_75t_L g11247 ( 
.A(n_10643),
.Y(n_11247)
);

OA21x2_ASAP7_75t_L g11248 ( 
.A1(n_10902),
.A2(n_10540),
.B(n_10245),
.Y(n_11248)
);

INVx1_ASAP7_75t_L g11249 ( 
.A(n_10786),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_L g11250 ( 
.A(n_11082),
.B(n_10276),
.Y(n_11250)
);

AO31x2_ASAP7_75t_L g11251 ( 
.A1(n_10908),
.A2(n_10583),
.A3(n_10452),
.B(n_10461),
.Y(n_11251)
);

OAI21x1_ASAP7_75t_L g11252 ( 
.A1(n_10668),
.A2(n_10440),
.B(n_10436),
.Y(n_11252)
);

BUFx6f_ASAP7_75t_L g11253 ( 
.A(n_10677),
.Y(n_11253)
);

INVx3_ASAP7_75t_L g11254 ( 
.A(n_11060),
.Y(n_11254)
);

NAND2xp5_ASAP7_75t_L g11255 ( 
.A(n_11090),
.B(n_10460),
.Y(n_11255)
);

OR2x2_ASAP7_75t_L g11256 ( 
.A(n_10653),
.B(n_10418),
.Y(n_11256)
);

BUFx2_ASAP7_75t_L g11257 ( 
.A(n_10676),
.Y(n_11257)
);

AND2x2_ASAP7_75t_L g11258 ( 
.A(n_11032),
.B(n_10204),
.Y(n_11258)
);

INVxp67_ASAP7_75t_L g11259 ( 
.A(n_11128),
.Y(n_11259)
);

INVx1_ASAP7_75t_L g11260 ( 
.A(n_10788),
.Y(n_11260)
);

AOI21xp5_ASAP7_75t_L g11261 ( 
.A1(n_10718),
.A2(n_10610),
.B(n_10576),
.Y(n_11261)
);

BUFx3_ASAP7_75t_L g11262 ( 
.A(n_10850),
.Y(n_11262)
);

NOR2xp33_ASAP7_75t_L g11263 ( 
.A(n_10647),
.B(n_10240),
.Y(n_11263)
);

AND2x2_ASAP7_75t_L g11264 ( 
.A(n_10791),
.B(n_10240),
.Y(n_11264)
);

CKINVDCx16_ASAP7_75t_R g11265 ( 
.A(n_10686),
.Y(n_11265)
);

AND2x4_ASAP7_75t_L g11266 ( 
.A(n_10990),
.B(n_10253),
.Y(n_11266)
);

O2A1O1Ixp33_ASAP7_75t_L g11267 ( 
.A1(n_10814),
.A2(n_10805),
.B(n_10730),
.C(n_10765),
.Y(n_11267)
);

INVx2_ASAP7_75t_SL g11268 ( 
.A(n_11016),
.Y(n_11268)
);

INVx1_ASAP7_75t_L g11269 ( 
.A(n_10819),
.Y(n_11269)
);

OAI21x1_ASAP7_75t_L g11270 ( 
.A1(n_10638),
.A2(n_10436),
.B(n_10317),
.Y(n_11270)
);

AND2x4_ASAP7_75t_L g11271 ( 
.A(n_10827),
.B(n_10253),
.Y(n_11271)
);

INVx1_ASAP7_75t_L g11272 ( 
.A(n_10874),
.Y(n_11272)
);

NAND2xp5_ASAP7_75t_L g11273 ( 
.A(n_11062),
.B(n_10436),
.Y(n_11273)
);

INVx1_ASAP7_75t_L g11274 ( 
.A(n_10708),
.Y(n_11274)
);

BUFx2_ASAP7_75t_L g11275 ( 
.A(n_11024),
.Y(n_11275)
);

CKINVDCx20_ASAP7_75t_R g11276 ( 
.A(n_10839),
.Y(n_11276)
);

NAND2xp33_ASAP7_75t_L g11277 ( 
.A(n_10688),
.B(n_10267),
.Y(n_11277)
);

BUFx6f_ASAP7_75t_L g11278 ( 
.A(n_10677),
.Y(n_11278)
);

INVx1_ASAP7_75t_L g11279 ( 
.A(n_10961),
.Y(n_11279)
);

INVx2_ASAP7_75t_SL g11280 ( 
.A(n_11016),
.Y(n_11280)
);

BUFx3_ASAP7_75t_L g11281 ( 
.A(n_10724),
.Y(n_11281)
);

INVx2_ASAP7_75t_L g11282 ( 
.A(n_11013),
.Y(n_11282)
);

NOR2xp33_ASAP7_75t_SL g11283 ( 
.A(n_10868),
.B(n_10420),
.Y(n_11283)
);

INVx1_ASAP7_75t_L g11284 ( 
.A(n_10711),
.Y(n_11284)
);

INVx2_ASAP7_75t_L g11285 ( 
.A(n_11130),
.Y(n_11285)
);

INVx1_ASAP7_75t_L g11286 ( 
.A(n_10717),
.Y(n_11286)
);

AOI21xp5_ASAP7_75t_L g11287 ( 
.A1(n_10795),
.A2(n_10413),
.B(n_10268),
.Y(n_11287)
);

AOI21xp5_ASAP7_75t_L g11288 ( 
.A1(n_10881),
.A2(n_10778),
.B(n_10733),
.Y(n_11288)
);

NAND2xp5_ASAP7_75t_SL g11289 ( 
.A(n_10662),
.B(n_10267),
.Y(n_11289)
);

AND2x2_ASAP7_75t_L g11290 ( 
.A(n_10981),
.B(n_10268),
.Y(n_11290)
);

A2O1A1Ixp33_ASAP7_75t_L g11291 ( 
.A1(n_10771),
.A2(n_10406),
.B(n_10431),
.C(n_10353),
.Y(n_11291)
);

AOI21xp5_ASAP7_75t_SL g11292 ( 
.A1(n_10825),
.A2(n_10406),
.B(n_10353),
.Y(n_11292)
);

NAND2xp5_ASAP7_75t_SL g11293 ( 
.A(n_10648),
.B(n_10431),
.Y(n_11293)
);

AOI21xp5_ASAP7_75t_L g11294 ( 
.A1(n_10731),
.A2(n_1165),
.B(n_1166),
.Y(n_11294)
);

NAND2xp5_ASAP7_75t_L g11295 ( 
.A(n_10674),
.B(n_1165),
.Y(n_11295)
);

AND2x4_ASAP7_75t_L g11296 ( 
.A(n_10672),
.B(n_1166),
.Y(n_11296)
);

INVx2_ASAP7_75t_L g11297 ( 
.A(n_10658),
.Y(n_11297)
);

INVx4_ASAP7_75t_L g11298 ( 
.A(n_10732),
.Y(n_11298)
);

INVx3_ASAP7_75t_L g11299 ( 
.A(n_10763),
.Y(n_11299)
);

OAI22xp5_ASAP7_75t_SL g11300 ( 
.A1(n_10776),
.A2(n_1169),
.B1(n_1167),
.B2(n_1168),
.Y(n_11300)
);

INVx1_ASAP7_75t_L g11301 ( 
.A(n_10704),
.Y(n_11301)
);

NAND2xp5_ASAP7_75t_SL g11302 ( 
.A(n_10656),
.B(n_10665),
.Y(n_11302)
);

OAI21xp33_ASAP7_75t_L g11303 ( 
.A1(n_10974),
.A2(n_1168),
.B(n_1169),
.Y(n_11303)
);

NAND2xp5_ASAP7_75t_L g11304 ( 
.A(n_10667),
.B(n_1170),
.Y(n_11304)
);

A2O1A1Ixp33_ASAP7_75t_L g11305 ( 
.A1(n_10982),
.A2(n_1172),
.B(n_1170),
.C(n_1171),
.Y(n_11305)
);

OR2x6_ASAP7_75t_L g11306 ( 
.A(n_11105),
.B(n_1171),
.Y(n_11306)
);

BUFx2_ASAP7_75t_L g11307 ( 
.A(n_10670),
.Y(n_11307)
);

NOR2xp33_ASAP7_75t_L g11308 ( 
.A(n_10831),
.B(n_1172),
.Y(n_11308)
);

OR2x2_ASAP7_75t_L g11309 ( 
.A(n_10675),
.B(n_1173),
.Y(n_11309)
);

AOI22xp33_ASAP7_75t_L g11310 ( 
.A1(n_11051),
.A2(n_1175),
.B1(n_1173),
.B2(n_1174),
.Y(n_11310)
);

NAND2xp5_ASAP7_75t_L g11311 ( 
.A(n_10645),
.B(n_1175),
.Y(n_11311)
);

INVx2_ASAP7_75t_L g11312 ( 
.A(n_10747),
.Y(n_11312)
);

OAI21xp5_ASAP7_75t_L g11313 ( 
.A1(n_10958),
.A2(n_1176),
.B(n_1177),
.Y(n_11313)
);

AOI22xp5_ASAP7_75t_L g11314 ( 
.A1(n_10750),
.A2(n_1178),
.B1(n_1176),
.B2(n_1177),
.Y(n_11314)
);

INVx1_ASAP7_75t_L g11315 ( 
.A(n_10828),
.Y(n_11315)
);

NOR3xp33_ASAP7_75t_L g11316 ( 
.A(n_10934),
.B(n_1178),
.C(n_1179),
.Y(n_11316)
);

BUFx6f_ASAP7_75t_L g11317 ( 
.A(n_10763),
.Y(n_11317)
);

INVx3_ASAP7_75t_SL g11318 ( 
.A(n_11127),
.Y(n_11318)
);

BUFx3_ASAP7_75t_L g11319 ( 
.A(n_11120),
.Y(n_11319)
);

AO21x1_ASAP7_75t_L g11320 ( 
.A1(n_10900),
.A2(n_1180),
.B(n_1181),
.Y(n_11320)
);

CKINVDCx5p33_ASAP7_75t_R g11321 ( 
.A(n_11092),
.Y(n_11321)
);

INVx2_ASAP7_75t_L g11322 ( 
.A(n_10965),
.Y(n_11322)
);

BUFx3_ASAP7_75t_L g11323 ( 
.A(n_10732),
.Y(n_11323)
);

INVx2_ASAP7_75t_L g11324 ( 
.A(n_10998),
.Y(n_11324)
);

OAI21xp5_ASAP7_75t_L g11325 ( 
.A1(n_10699),
.A2(n_1180),
.B(n_1182),
.Y(n_11325)
);

AOI21xp5_ASAP7_75t_L g11326 ( 
.A1(n_11022),
.A2(n_1182),
.B(n_1183),
.Y(n_11326)
);

BUFx6f_ASAP7_75t_L g11327 ( 
.A(n_10808),
.Y(n_11327)
);

A2O1A1Ixp33_ASAP7_75t_SL g11328 ( 
.A1(n_10734),
.A2(n_10772),
.B(n_10803),
.C(n_10796),
.Y(n_11328)
);

NAND2xp5_ASAP7_75t_L g11329 ( 
.A(n_10645),
.B(n_1183),
.Y(n_11329)
);

AOI21xp5_ASAP7_75t_L g11330 ( 
.A1(n_11033),
.A2(n_1185),
.B(n_1186),
.Y(n_11330)
);

OAI21xp5_ASAP7_75t_L g11331 ( 
.A1(n_10818),
.A2(n_1185),
.B(n_1187),
.Y(n_11331)
);

INVx1_ASAP7_75t_L g11332 ( 
.A(n_10851),
.Y(n_11332)
);

INVx1_ASAP7_75t_L g11333 ( 
.A(n_10854),
.Y(n_11333)
);

AOI21xp33_ASAP7_75t_L g11334 ( 
.A1(n_10914),
.A2(n_1188),
.B(n_1189),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_SL g11335 ( 
.A(n_10673),
.B(n_1188),
.Y(n_11335)
);

OR2x2_ASAP7_75t_SL g11336 ( 
.A(n_10997),
.B(n_1189),
.Y(n_11336)
);

INVx2_ASAP7_75t_SL g11337 ( 
.A(n_10691),
.Y(n_11337)
);

INVxp67_ASAP7_75t_L g11338 ( 
.A(n_11005),
.Y(n_11338)
);

NAND2xp5_ASAP7_75t_L g11339 ( 
.A(n_10738),
.B(n_1190),
.Y(n_11339)
);

AND2x4_ASAP7_75t_L g11340 ( 
.A(n_10876),
.B(n_1190),
.Y(n_11340)
);

A2O1A1Ixp33_ASAP7_75t_L g11341 ( 
.A1(n_11029),
.A2(n_1193),
.B(n_1191),
.C(n_1192),
.Y(n_11341)
);

INVx2_ASAP7_75t_L g11342 ( 
.A(n_10862),
.Y(n_11342)
);

INVx1_ASAP7_75t_SL g11343 ( 
.A(n_10885),
.Y(n_11343)
);

INVx1_ASAP7_75t_L g11344 ( 
.A(n_10860),
.Y(n_11344)
);

AND2x2_ASAP7_75t_L g11345 ( 
.A(n_10911),
.B(n_1191),
.Y(n_11345)
);

NAND2xp5_ASAP7_75t_L g11346 ( 
.A(n_10705),
.B(n_10979),
.Y(n_11346)
);

BUFx6f_ASAP7_75t_L g11347 ( 
.A(n_10808),
.Y(n_11347)
);

INVx3_ASAP7_75t_L g11348 ( 
.A(n_10892),
.Y(n_11348)
);

NAND2xp5_ASAP7_75t_L g11349 ( 
.A(n_10970),
.B(n_1192),
.Y(n_11349)
);

AOI22xp5_ASAP7_75t_L g11350 ( 
.A1(n_10897),
.A2(n_1195),
.B1(n_1193),
.B2(n_1194),
.Y(n_11350)
);

NAND2xp5_ASAP7_75t_L g11351 ( 
.A(n_10817),
.B(n_1194),
.Y(n_11351)
);

OAI22xp5_ASAP7_75t_L g11352 ( 
.A1(n_10762),
.A2(n_1197),
.B1(n_1195),
.B2(n_1196),
.Y(n_11352)
);

AOI21xp5_ASAP7_75t_L g11353 ( 
.A1(n_11040),
.A2(n_1196),
.B(n_1198),
.Y(n_11353)
);

AO21x2_ASAP7_75t_L g11354 ( 
.A1(n_10727),
.A2(n_1198),
.B(n_1199),
.Y(n_11354)
);

INVx1_ASAP7_75t_L g11355 ( 
.A(n_10746),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_10767),
.Y(n_11356)
);

INVx2_ASAP7_75t_L g11357 ( 
.A(n_10865),
.Y(n_11357)
);

HB1xp67_ASAP7_75t_L g11358 ( 
.A(n_10872),
.Y(n_11358)
);

NAND2xp5_ASAP7_75t_SL g11359 ( 
.A(n_11045),
.B(n_1199),
.Y(n_11359)
);

AND2x2_ASAP7_75t_L g11360 ( 
.A(n_10960),
.B(n_1200),
.Y(n_11360)
);

AND2x4_ASAP7_75t_L g11361 ( 
.A(n_10917),
.B(n_1201),
.Y(n_11361)
);

AOI21xp5_ASAP7_75t_L g11362 ( 
.A1(n_11071),
.A2(n_1201),
.B(n_1202),
.Y(n_11362)
);

INVx5_ASAP7_75t_L g11363 ( 
.A(n_11115),
.Y(n_11363)
);

HB1xp67_ASAP7_75t_L g11364 ( 
.A(n_10878),
.Y(n_11364)
);

OR2x2_ASAP7_75t_L g11365 ( 
.A(n_10790),
.B(n_1202),
.Y(n_11365)
);

INVx1_ASAP7_75t_L g11366 ( 
.A(n_10792),
.Y(n_11366)
);

A2O1A1Ixp33_ASAP7_75t_L g11367 ( 
.A1(n_10826),
.A2(n_1205),
.B(n_1203),
.C(n_1204),
.Y(n_11367)
);

BUFx6f_ASAP7_75t_L g11368 ( 
.A(n_10892),
.Y(n_11368)
);

OAI221xp5_ASAP7_75t_L g11369 ( 
.A1(n_10840),
.A2(n_1206),
.B1(n_1204),
.B2(n_1205),
.C(n_1207),
.Y(n_11369)
);

INVxp67_ASAP7_75t_L g11370 ( 
.A(n_11095),
.Y(n_11370)
);

INVx1_ASAP7_75t_L g11371 ( 
.A(n_10800),
.Y(n_11371)
);

AND2x2_ASAP7_75t_L g11372 ( 
.A(n_11002),
.B(n_1206),
.Y(n_11372)
);

NAND2x1p5_ASAP7_75t_L g11373 ( 
.A(n_10680),
.B(n_1207),
.Y(n_11373)
);

INVx4_ASAP7_75t_L g11374 ( 
.A(n_10973),
.Y(n_11374)
);

O2A1O1Ixp33_ASAP7_75t_L g11375 ( 
.A1(n_10690),
.A2(n_1210),
.B(n_1208),
.C(n_1209),
.Y(n_11375)
);

OAI21xp5_ASAP7_75t_L g11376 ( 
.A1(n_10844),
.A2(n_1208),
.B(n_1209),
.Y(n_11376)
);

O2A1O1Ixp33_ASAP7_75t_L g11377 ( 
.A1(n_11068),
.A2(n_11080),
.B(n_10685),
.C(n_10899),
.Y(n_11377)
);

NAND2xp5_ASAP7_75t_L g11378 ( 
.A(n_10812),
.B(n_1211),
.Y(n_11378)
);

OAI22xp5_ASAP7_75t_L g11379 ( 
.A1(n_10938),
.A2(n_1214),
.B1(n_1212),
.B2(n_1213),
.Y(n_11379)
);

INVx2_ASAP7_75t_L g11380 ( 
.A(n_10870),
.Y(n_11380)
);

INVx1_ASAP7_75t_L g11381 ( 
.A(n_10821),
.Y(n_11381)
);

INVx1_ASAP7_75t_L g11382 ( 
.A(n_10890),
.Y(n_11382)
);

AO21x2_ASAP7_75t_L g11383 ( 
.A1(n_10895),
.A2(n_1212),
.B(n_1213),
.Y(n_11383)
);

INVx1_ASAP7_75t_L g11384 ( 
.A(n_10893),
.Y(n_11384)
);

BUFx2_ASAP7_75t_L g11385 ( 
.A(n_10944),
.Y(n_11385)
);

AOI22xp33_ASAP7_75t_L g11386 ( 
.A1(n_10820),
.A2(n_1216),
.B1(n_1214),
.B2(n_1215),
.Y(n_11386)
);

NAND2xp5_ASAP7_75t_L g11387 ( 
.A(n_10901),
.B(n_1215),
.Y(n_11387)
);

OR2x6_ASAP7_75t_L g11388 ( 
.A(n_11115),
.B(n_11123),
.Y(n_11388)
);

AO32x2_ASAP7_75t_L g11389 ( 
.A1(n_10709),
.A2(n_1218),
.A3(n_1216),
.B1(n_1217),
.B2(n_1219),
.Y(n_11389)
);

INVx1_ASAP7_75t_L g11390 ( 
.A(n_10906),
.Y(n_11390)
);

OR2x2_ASAP7_75t_L g11391 ( 
.A(n_11038),
.B(n_1217),
.Y(n_11391)
);

INVx3_ASAP7_75t_SL g11392 ( 
.A(n_10640),
.Y(n_11392)
);

OAI21x1_ASAP7_75t_L g11393 ( 
.A1(n_10694),
.A2(n_10683),
.B(n_10823),
.Y(n_11393)
);

AND2x4_ASAP7_75t_L g11394 ( 
.A(n_11107),
.B(n_1218),
.Y(n_11394)
);

NAND2x1p5_ASAP7_75t_L g11395 ( 
.A(n_10774),
.B(n_1219),
.Y(n_11395)
);

A2O1A1Ixp33_ASAP7_75t_SL g11396 ( 
.A1(n_10846),
.A2(n_1222),
.B(n_1220),
.C(n_1221),
.Y(n_11396)
);

INVx3_ASAP7_75t_L g11397 ( 
.A(n_10973),
.Y(n_11397)
);

AND2x4_ASAP7_75t_L g11398 ( 
.A(n_10682),
.B(n_1220),
.Y(n_11398)
);

AOI21xp5_ASAP7_75t_L g11399 ( 
.A1(n_10707),
.A2(n_11010),
.B(n_10830),
.Y(n_11399)
);

AOI22xp5_ASAP7_75t_L g11400 ( 
.A1(n_11041),
.A2(n_1224),
.B1(n_1222),
.B2(n_1223),
.Y(n_11400)
);

OAI22xp5_ASAP7_75t_L g11401 ( 
.A1(n_10941),
.A2(n_1227),
.B1(n_1224),
.B2(n_1226),
.Y(n_11401)
);

NAND2xp5_ASAP7_75t_L g11402 ( 
.A(n_10689),
.B(n_1226),
.Y(n_11402)
);

INVx2_ASAP7_75t_L g11403 ( 
.A(n_10924),
.Y(n_11403)
);

NOR2xp33_ASAP7_75t_R g11404 ( 
.A(n_10936),
.B(n_1227),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_10943),
.Y(n_11405)
);

INVx1_ASAP7_75t_L g11406 ( 
.A(n_10801),
.Y(n_11406)
);

NAND2xp5_ASAP7_75t_L g11407 ( 
.A(n_10684),
.B(n_1228),
.Y(n_11407)
);

AND2x4_ASAP7_75t_L g11408 ( 
.A(n_11056),
.B(n_1228),
.Y(n_11408)
);

BUFx6f_ASAP7_75t_L g11409 ( 
.A(n_11020),
.Y(n_11409)
);

AOI21xp5_ASAP7_75t_L g11410 ( 
.A1(n_11042),
.A2(n_1229),
.B(n_1230),
.Y(n_11410)
);

AOI21xp5_ASAP7_75t_L g11411 ( 
.A1(n_11049),
.A2(n_1229),
.B(n_1231),
.Y(n_11411)
);

BUFx6f_ASAP7_75t_L g11412 ( 
.A(n_11020),
.Y(n_11412)
);

NAND2xp5_ASAP7_75t_L g11413 ( 
.A(n_11086),
.B(n_1232),
.Y(n_11413)
);

AOI21xp5_ASAP7_75t_L g11414 ( 
.A1(n_10856),
.A2(n_1232),
.B(n_1233),
.Y(n_11414)
);

BUFx12f_ASAP7_75t_L g11415 ( 
.A(n_10794),
.Y(n_11415)
);

INVx1_ASAP7_75t_L g11416 ( 
.A(n_10813),
.Y(n_11416)
);

INVx1_ASAP7_75t_L g11417 ( 
.A(n_10824),
.Y(n_11417)
);

AND2x2_ASAP7_75t_L g11418 ( 
.A(n_10931),
.B(n_1233),
.Y(n_11418)
);

INVx2_ASAP7_75t_SL g11419 ( 
.A(n_10880),
.Y(n_11419)
);

BUFx3_ASAP7_75t_L g11420 ( 
.A(n_10836),
.Y(n_11420)
);

BUFx3_ASAP7_75t_L g11421 ( 
.A(n_10848),
.Y(n_11421)
);

INVx3_ASAP7_75t_L g11422 ( 
.A(n_10909),
.Y(n_11422)
);

INVx3_ASAP7_75t_L g11423 ( 
.A(n_10933),
.Y(n_11423)
);

A2O1A1Ixp33_ASAP7_75t_L g11424 ( 
.A1(n_10992),
.A2(n_10715),
.B(n_10955),
.C(n_10952),
.Y(n_11424)
);

AND2x4_ASAP7_75t_L g11425 ( 
.A(n_10896),
.B(n_1234),
.Y(n_11425)
);

NOR2x1_ASAP7_75t_L g11426 ( 
.A(n_10835),
.B(n_1234),
.Y(n_11426)
);

INVx2_ASAP7_75t_L g11427 ( 
.A(n_10948),
.Y(n_11427)
);

INVx3_ASAP7_75t_L g11428 ( 
.A(n_10822),
.Y(n_11428)
);

INVx1_ASAP7_75t_L g11429 ( 
.A(n_10855),
.Y(n_11429)
);

AOI22xp33_ASAP7_75t_SL g11430 ( 
.A1(n_11081),
.A2(n_1237),
.B1(n_1235),
.B2(n_1236),
.Y(n_11430)
);

AO21x2_ASAP7_75t_L g11431 ( 
.A1(n_10898),
.A2(n_1236),
.B(n_1238),
.Y(n_11431)
);

INVx1_ASAP7_75t_L g11432 ( 
.A(n_10951),
.Y(n_11432)
);

BUFx3_ASAP7_75t_L g11433 ( 
.A(n_10712),
.Y(n_11433)
);

BUFx3_ASAP7_75t_L g11434 ( 
.A(n_11057),
.Y(n_11434)
);

HB1xp67_ASAP7_75t_L g11435 ( 
.A(n_10954),
.Y(n_11435)
);

OAI22xp5_ASAP7_75t_L g11436 ( 
.A1(n_10749),
.A2(n_1240),
.B1(n_1238),
.B2(n_1239),
.Y(n_11436)
);

NAND2x1_ASAP7_75t_L g11437 ( 
.A(n_10692),
.B(n_1239),
.Y(n_11437)
);

INVx3_ASAP7_75t_L g11438 ( 
.A(n_10949),
.Y(n_11438)
);

NAND2xp5_ASAP7_75t_L g11439 ( 
.A(n_10929),
.B(n_1241),
.Y(n_11439)
);

AND2x2_ASAP7_75t_L g11440 ( 
.A(n_10940),
.B(n_1241),
.Y(n_11440)
);

HB1xp67_ASAP7_75t_L g11441 ( 
.A(n_10742),
.Y(n_11441)
);

BUFx6f_ASAP7_75t_L g11442 ( 
.A(n_10748),
.Y(n_11442)
);

OAI22xp5_ASAP7_75t_L g11443 ( 
.A1(n_10946),
.A2(n_1244),
.B1(n_1242),
.B2(n_1243),
.Y(n_11443)
);

INVx4_ASAP7_75t_L g11444 ( 
.A(n_11097),
.Y(n_11444)
);

OAI22xp5_ASAP7_75t_L g11445 ( 
.A1(n_10867),
.A2(n_1246),
.B1(n_1242),
.B2(n_1245),
.Y(n_11445)
);

INVx1_ASAP7_75t_L g11446 ( 
.A(n_10913),
.Y(n_11446)
);

BUFx2_ASAP7_75t_L g11447 ( 
.A(n_10679),
.Y(n_11447)
);

NOR2xp67_ASAP7_75t_SL g11448 ( 
.A(n_11074),
.B(n_1247),
.Y(n_11448)
);

AOI21xp33_ASAP7_75t_SL g11449 ( 
.A1(n_10695),
.A2(n_1248),
.B(n_1249),
.Y(n_11449)
);

NAND2x1_ASAP7_75t_SL g11450 ( 
.A(n_10968),
.B(n_1249),
.Y(n_11450)
);

INVx3_ASAP7_75t_L g11451 ( 
.A(n_10681),
.Y(n_11451)
);

AND2x4_ASAP7_75t_L g11452 ( 
.A(n_10756),
.B(n_1250),
.Y(n_11452)
);

OAI22xp5_ASAP7_75t_L g11453 ( 
.A1(n_10978),
.A2(n_1252),
.B1(n_1250),
.B2(n_1251),
.Y(n_11453)
);

A2O1A1Ixp33_ASAP7_75t_SL g11454 ( 
.A1(n_10875),
.A2(n_1255),
.B(n_1253),
.C(n_1254),
.Y(n_11454)
);

OR2x2_ASAP7_75t_L g11455 ( 
.A(n_11052),
.B(n_11046),
.Y(n_11455)
);

INVx2_ASAP7_75t_SL g11456 ( 
.A(n_10915),
.Y(n_11456)
);

BUFx2_ASAP7_75t_SL g11457 ( 
.A(n_11126),
.Y(n_11457)
);

BUFx2_ASAP7_75t_L g11458 ( 
.A(n_10720),
.Y(n_11458)
);

HB1xp67_ASAP7_75t_L g11459 ( 
.A(n_10869),
.Y(n_11459)
);

INVx1_ASAP7_75t_L g11460 ( 
.A(n_10837),
.Y(n_11460)
);

NAND2xp5_ASAP7_75t_SL g11461 ( 
.A(n_10650),
.B(n_1254),
.Y(n_11461)
);

AND2x4_ASAP7_75t_L g11462 ( 
.A(n_10995),
.B(n_1255),
.Y(n_11462)
);

AND2x4_ASAP7_75t_L g11463 ( 
.A(n_10999),
.B(n_1256),
.Y(n_11463)
);

INVx2_ASAP7_75t_SL g11464 ( 
.A(n_11012),
.Y(n_11464)
);

INVx1_ASAP7_75t_L g11465 ( 
.A(n_10837),
.Y(n_11465)
);

NOR2x1_ASAP7_75t_SL g11466 ( 
.A(n_11018),
.B(n_1256),
.Y(n_11466)
);

INVx1_ASAP7_75t_L g11467 ( 
.A(n_10894),
.Y(n_11467)
);

INVx2_ASAP7_75t_SL g11468 ( 
.A(n_11011),
.Y(n_11468)
);

INVx1_ASAP7_75t_L g11469 ( 
.A(n_10905),
.Y(n_11469)
);

AOI222xp33_ASAP7_75t_L g11470 ( 
.A1(n_11015),
.A2(n_1260),
.B1(n_1262),
.B2(n_1257),
.C1(n_1258),
.C2(n_1261),
.Y(n_11470)
);

NOR2xp33_ASAP7_75t_L g11471 ( 
.A(n_11043),
.B(n_1257),
.Y(n_11471)
);

OAI22xp5_ASAP7_75t_L g11472 ( 
.A1(n_10975),
.A2(n_1263),
.B1(n_1258),
.B2(n_1260),
.Y(n_11472)
);

NAND3xp33_ASAP7_75t_SL g11473 ( 
.A(n_11108),
.B(n_1264),
.C(n_1265),
.Y(n_11473)
);

AO21x1_ASAP7_75t_L g11474 ( 
.A1(n_10910),
.A2(n_1264),
.B(n_1266),
.Y(n_11474)
);

OR2x2_ASAP7_75t_L g11475 ( 
.A(n_11047),
.B(n_1267),
.Y(n_11475)
);

INVx1_ASAP7_75t_SL g11476 ( 
.A(n_10983),
.Y(n_11476)
);

BUFx6f_ASAP7_75t_L g11477 ( 
.A(n_10993),
.Y(n_11477)
);

AND2x2_ASAP7_75t_L g11478 ( 
.A(n_10879),
.B(n_1267),
.Y(n_11478)
);

NAND2xp5_ASAP7_75t_L g11479 ( 
.A(n_11007),
.B(n_1268),
.Y(n_11479)
);

NOR2xp33_ASAP7_75t_L g11480 ( 
.A(n_11014),
.B(n_11017),
.Y(n_11480)
);

INVx2_ASAP7_75t_SL g11481 ( 
.A(n_11048),
.Y(n_11481)
);

INVx1_ASAP7_75t_L g11482 ( 
.A(n_10912),
.Y(n_11482)
);

INVx2_ASAP7_75t_L g11483 ( 
.A(n_10802),
.Y(n_11483)
);

NOR2x1_ASAP7_75t_SL g11484 ( 
.A(n_10921),
.B(n_10758),
.Y(n_11484)
);

AOI22xp33_ASAP7_75t_SL g11485 ( 
.A1(n_11085),
.A2(n_1272),
.B1(n_1269),
.B2(n_1271),
.Y(n_11485)
);

INVx4_ASAP7_75t_L g11486 ( 
.A(n_11064),
.Y(n_11486)
);

NAND2xp5_ASAP7_75t_L g11487 ( 
.A(n_11008),
.B(n_1269),
.Y(n_11487)
);

HB1xp67_ASAP7_75t_L g11488 ( 
.A(n_10882),
.Y(n_11488)
);

NAND2xp33_ASAP7_75t_L g11489 ( 
.A(n_10726),
.B(n_1271),
.Y(n_11489)
);

AOI21xp5_ASAP7_75t_L g11490 ( 
.A1(n_10783),
.A2(n_1272),
.B(n_1273),
.Y(n_11490)
);

NOR2x1_ASAP7_75t_L g11491 ( 
.A(n_11113),
.B(n_1274),
.Y(n_11491)
);

AOI21xp5_ASAP7_75t_L g11492 ( 
.A1(n_11087),
.A2(n_1274),
.B(n_1275),
.Y(n_11492)
);

BUFx3_ASAP7_75t_L g11493 ( 
.A(n_11119),
.Y(n_11493)
);

INVx5_ASAP7_75t_L g11494 ( 
.A(n_11079),
.Y(n_11494)
);

AND2x2_ASAP7_75t_L g11495 ( 
.A(n_10887),
.B(n_1276),
.Y(n_11495)
);

INVx1_ASAP7_75t_L g11496 ( 
.A(n_10920),
.Y(n_11496)
);

AOI22xp33_ASAP7_75t_L g11497 ( 
.A1(n_10959),
.A2(n_1279),
.B1(n_1277),
.B2(n_1278),
.Y(n_11497)
);

NOR2xp33_ASAP7_75t_SL g11498 ( 
.A(n_10700),
.B(n_1279),
.Y(n_11498)
);

BUFx3_ASAP7_75t_L g11499 ( 
.A(n_11122),
.Y(n_11499)
);

OAI22xp5_ASAP7_75t_L g11500 ( 
.A1(n_10975),
.A2(n_1282),
.B1(n_1280),
.B2(n_1281),
.Y(n_11500)
);

NAND2xp5_ASAP7_75t_L g11501 ( 
.A(n_11083),
.B(n_1281),
.Y(n_11501)
);

OR2x6_ASAP7_75t_L g11502 ( 
.A(n_10757),
.B(n_1282),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_10891),
.B(n_1283),
.Y(n_11503)
);

OAI22xp5_ASAP7_75t_L g11504 ( 
.A1(n_11099),
.A2(n_1285),
.B1(n_1283),
.B2(n_1284),
.Y(n_11504)
);

INVx1_ASAP7_75t_L g11505 ( 
.A(n_10930),
.Y(n_11505)
);

OR2x2_ASAP7_75t_L g11506 ( 
.A(n_11050),
.B(n_1285),
.Y(n_11506)
);

NAND2xp5_ASAP7_75t_L g11507 ( 
.A(n_11094),
.B(n_11129),
.Y(n_11507)
);

INVx2_ASAP7_75t_L g11508 ( 
.A(n_11451),
.Y(n_11508)
);

BUFx8_ASAP7_75t_L g11509 ( 
.A(n_11177),
.Y(n_11509)
);

BUFx8_ASAP7_75t_L g11510 ( 
.A(n_11160),
.Y(n_11510)
);

OAI22xp5_ASAP7_75t_L g11511 ( 
.A1(n_11222),
.A2(n_10918),
.B1(n_11093),
.B2(n_10985),
.Y(n_11511)
);

INVx1_ASAP7_75t_SL g11512 ( 
.A(n_11196),
.Y(n_11512)
);

INVx1_ASAP7_75t_SL g11513 ( 
.A(n_11318),
.Y(n_11513)
);

INVx5_ASAP7_75t_L g11514 ( 
.A(n_11160),
.Y(n_11514)
);

CKINVDCx20_ASAP7_75t_R g11515 ( 
.A(n_11276),
.Y(n_11515)
);

INVx3_ASAP7_75t_L g11516 ( 
.A(n_11281),
.Y(n_11516)
);

OAI22xp5_ASAP7_75t_L g11517 ( 
.A1(n_11306),
.A2(n_11064),
.B1(n_11075),
.B2(n_11004),
.Y(n_11517)
);

INVx6_ASAP7_75t_L g11518 ( 
.A(n_11245),
.Y(n_11518)
);

NAND2xp5_ASAP7_75t_L g11519 ( 
.A(n_11237),
.B(n_11103),
.Y(n_11519)
);

BUFx2_ASAP7_75t_SL g11520 ( 
.A(n_11494),
.Y(n_11520)
);

INVx1_ASAP7_75t_L g11521 ( 
.A(n_11140),
.Y(n_11521)
);

INVx1_ASAP7_75t_L g11522 ( 
.A(n_11150),
.Y(n_11522)
);

CKINVDCx20_ASAP7_75t_R g11523 ( 
.A(n_11265),
.Y(n_11523)
);

BUFx12f_ASAP7_75t_L g11524 ( 
.A(n_11136),
.Y(n_11524)
);

BUFx8_ASAP7_75t_L g11525 ( 
.A(n_11345),
.Y(n_11525)
);

INVx1_ASAP7_75t_L g11526 ( 
.A(n_11155),
.Y(n_11526)
);

CKINVDCx11_ASAP7_75t_R g11527 ( 
.A(n_11392),
.Y(n_11527)
);

OAI22xp5_ASAP7_75t_L g11528 ( 
.A1(n_11306),
.A2(n_11075),
.B1(n_11106),
.B2(n_11088),
.Y(n_11528)
);

CKINVDCx5p33_ASAP7_75t_R g11529 ( 
.A(n_11210),
.Y(n_11529)
);

INVx1_ASAP7_75t_L g11530 ( 
.A(n_11166),
.Y(n_11530)
);

OAI22xp5_ASAP7_75t_L g11531 ( 
.A1(n_11502),
.A2(n_10698),
.B1(n_11035),
.B2(n_11003),
.Y(n_11531)
);

CKINVDCx5p33_ASAP7_75t_R g11532 ( 
.A(n_11262),
.Y(n_11532)
);

OAI22xp33_ASAP7_75t_L g11533 ( 
.A1(n_11502),
.A2(n_10753),
.B1(n_11000),
.B2(n_10939),
.Y(n_11533)
);

AOI22xp33_ASAP7_75t_SL g11534 ( 
.A1(n_11484),
.A2(n_10986),
.B1(n_11098),
.B2(n_11067),
.Y(n_11534)
);

AOI22xp33_ASAP7_75t_L g11535 ( 
.A1(n_11288),
.A2(n_11065),
.B1(n_10922),
.B2(n_10809),
.Y(n_11535)
);

BUFx3_ASAP7_75t_L g11536 ( 
.A(n_11226),
.Y(n_11536)
);

INVx2_ASAP7_75t_L g11537 ( 
.A(n_11483),
.Y(n_11537)
);

BUFx6f_ASAP7_75t_L g11538 ( 
.A(n_11191),
.Y(n_11538)
);

NAND2xp5_ASAP7_75t_L g11539 ( 
.A(n_11432),
.B(n_11110),
.Y(n_11539)
);

OAI22xp33_ASAP7_75t_L g11540 ( 
.A1(n_11486),
.A2(n_11388),
.B1(n_11146),
.B2(n_11363),
.Y(n_11540)
);

CKINVDCx11_ASAP7_75t_R g11541 ( 
.A(n_11216),
.Y(n_11541)
);

INVx1_ASAP7_75t_L g11542 ( 
.A(n_11173),
.Y(n_11542)
);

INVx2_ASAP7_75t_L g11543 ( 
.A(n_11194),
.Y(n_11543)
);

AOI22xp33_ASAP7_75t_SL g11544 ( 
.A1(n_11179),
.A2(n_10721),
.B1(n_11073),
.B2(n_11078),
.Y(n_11544)
);

AOI22xp33_ASAP7_75t_SL g11545 ( 
.A1(n_11178),
.A2(n_11331),
.B1(n_11376),
.B2(n_11457),
.Y(n_11545)
);

INVx1_ASAP7_75t_L g11546 ( 
.A(n_11174),
.Y(n_11546)
);

NAND2x1p5_ASAP7_75t_L g11547 ( 
.A(n_11176),
.B(n_11076),
.Y(n_11547)
);

AOI22xp33_ASAP7_75t_L g11548 ( 
.A1(n_11212),
.A2(n_10728),
.B1(n_11061),
.B2(n_11025),
.Y(n_11548)
);

OAI22xp5_ASAP7_75t_L g11549 ( 
.A1(n_11305),
.A2(n_10926),
.B1(n_10942),
.B2(n_10967),
.Y(n_11549)
);

AOI21xp5_ASAP7_75t_SL g11550 ( 
.A1(n_11161),
.A2(n_10737),
.B(n_10740),
.Y(n_11550)
);

OAI22xp33_ASAP7_75t_L g11551 ( 
.A1(n_11388),
.A2(n_10925),
.B1(n_10916),
.B2(n_10971),
.Y(n_11551)
);

OR2x2_ASAP7_75t_L g11552 ( 
.A(n_11247),
.B(n_11118),
.Y(n_11552)
);

HB1xp67_ASAP7_75t_L g11553 ( 
.A(n_11157),
.Y(n_11553)
);

BUFx3_ASAP7_75t_L g11554 ( 
.A(n_11415),
.Y(n_11554)
);

INVx1_ASAP7_75t_L g11555 ( 
.A(n_11185),
.Y(n_11555)
);

CKINVDCx5p33_ASAP7_75t_R g11556 ( 
.A(n_11211),
.Y(n_11556)
);

INVx6_ASAP7_75t_L g11557 ( 
.A(n_11148),
.Y(n_11557)
);

OAI22xp5_ASAP7_75t_L g11558 ( 
.A1(n_11314),
.A2(n_10977),
.B1(n_10987),
.B2(n_10903),
.Y(n_11558)
);

AOI22xp33_ASAP7_75t_L g11559 ( 
.A1(n_11316),
.A2(n_10994),
.B1(n_10988),
.B2(n_11104),
.Y(n_11559)
);

AOI22xp33_ASAP7_75t_L g11560 ( 
.A1(n_11158),
.A2(n_11111),
.B1(n_10871),
.B2(n_11070),
.Y(n_11560)
);

AOI22xp33_ASAP7_75t_SL g11561 ( 
.A1(n_11369),
.A2(n_10697),
.B1(n_10702),
.B2(n_10775),
.Y(n_11561)
);

INVx2_ASAP7_75t_L g11562 ( 
.A(n_11202),
.Y(n_11562)
);

CKINVDCx20_ASAP7_75t_R g11563 ( 
.A(n_11319),
.Y(n_11563)
);

INVx1_ASAP7_75t_L g11564 ( 
.A(n_11197),
.Y(n_11564)
);

BUFx2_ASAP7_75t_L g11565 ( 
.A(n_11135),
.Y(n_11565)
);

AOI22xp33_ASAP7_75t_L g11566 ( 
.A1(n_11399),
.A2(n_11091),
.B1(n_10845),
.B2(n_11112),
.Y(n_11566)
);

CKINVDCx11_ASAP7_75t_R g11567 ( 
.A(n_11148),
.Y(n_11567)
);

OAI21xp33_ASAP7_75t_L g11568 ( 
.A1(n_11341),
.A2(n_11303),
.B(n_11424),
.Y(n_11568)
);

INVx6_ASAP7_75t_L g11569 ( 
.A(n_11298),
.Y(n_11569)
);

INVx1_ASAP7_75t_L g11570 ( 
.A(n_11200),
.Y(n_11570)
);

AOI22xp5_ASAP7_75t_L g11571 ( 
.A1(n_11448),
.A2(n_11489),
.B1(n_11359),
.B2(n_11470),
.Y(n_11571)
);

AOI22xp33_ASAP7_75t_SL g11572 ( 
.A1(n_11363),
.A2(n_10804),
.B1(n_10953),
.B2(n_10866),
.Y(n_11572)
);

INVx1_ASAP7_75t_SL g11573 ( 
.A(n_11447),
.Y(n_11573)
);

CKINVDCx5p33_ASAP7_75t_R g11574 ( 
.A(n_11192),
.Y(n_11574)
);

AOI22xp33_ASAP7_75t_L g11575 ( 
.A1(n_11326),
.A2(n_11037),
.B1(n_10861),
.B2(n_10807),
.Y(n_11575)
);

INVx6_ASAP7_75t_L g11576 ( 
.A(n_11227),
.Y(n_11576)
);

INVx1_ASAP7_75t_L g11577 ( 
.A(n_11149),
.Y(n_11577)
);

INVx6_ASAP7_75t_L g11578 ( 
.A(n_11323),
.Y(n_11578)
);

AOI22xp33_ASAP7_75t_SL g11579 ( 
.A1(n_11204),
.A2(n_11498),
.B1(n_11248),
.B2(n_11353),
.Y(n_11579)
);

AOI22xp33_ASAP7_75t_L g11580 ( 
.A1(n_11330),
.A2(n_11362),
.B1(n_11430),
.B2(n_11243),
.Y(n_11580)
);

BUFx12f_ASAP7_75t_L g11581 ( 
.A(n_11321),
.Y(n_11581)
);

AOI22xp33_ASAP7_75t_L g11582 ( 
.A1(n_11492),
.A2(n_10843),
.B1(n_10859),
.B2(n_11102),
.Y(n_11582)
);

OAI22xp33_ASAP7_75t_L g11583 ( 
.A1(n_11273),
.A2(n_10884),
.B1(n_10764),
.B2(n_11114),
.Y(n_11583)
);

AOI22xp33_ASAP7_75t_L g11584 ( 
.A1(n_11294),
.A2(n_10723),
.B1(n_11069),
.B2(n_11125),
.Y(n_11584)
);

NAND2xp5_ASAP7_75t_L g11585 ( 
.A(n_11382),
.B(n_11384),
.Y(n_11585)
);

INVx1_ASAP7_75t_L g11586 ( 
.A(n_11154),
.Y(n_11586)
);

INVx5_ASAP7_75t_L g11587 ( 
.A(n_11494),
.Y(n_11587)
);

INVx1_ASAP7_75t_L g11588 ( 
.A(n_11165),
.Y(n_11588)
);

INVx1_ASAP7_75t_L g11589 ( 
.A(n_11172),
.Y(n_11589)
);

NAND2xp5_ASAP7_75t_L g11590 ( 
.A(n_11390),
.B(n_11124),
.Y(n_11590)
);

INVx1_ASAP7_75t_L g11591 ( 
.A(n_11181),
.Y(n_11591)
);

AOI22xp33_ASAP7_75t_L g11592 ( 
.A1(n_11414),
.A2(n_10713),
.B1(n_11021),
.B2(n_11019),
.Y(n_11592)
);

BUFx6f_ASAP7_75t_L g11593 ( 
.A(n_11215),
.Y(n_11593)
);

BUFx4f_ASAP7_75t_SL g11594 ( 
.A(n_11141),
.Y(n_11594)
);

OAI22xp5_ASAP7_75t_L g11595 ( 
.A1(n_11152),
.A2(n_10793),
.B1(n_10877),
.B2(n_10816),
.Y(n_11595)
);

INVx2_ASAP7_75t_L g11596 ( 
.A(n_11188),
.Y(n_11596)
);

AOI22xp33_ASAP7_75t_SL g11597 ( 
.A1(n_11313),
.A2(n_11030),
.B1(n_11054),
.B2(n_11072),
.Y(n_11597)
);

INVx2_ASAP7_75t_L g11598 ( 
.A(n_11193),
.Y(n_11598)
);

INVx2_ASAP7_75t_L g11599 ( 
.A(n_11198),
.Y(n_11599)
);

INVx2_ASAP7_75t_L g11600 ( 
.A(n_11206),
.Y(n_11600)
);

AOI22xp33_ASAP7_75t_SL g11601 ( 
.A1(n_11325),
.A2(n_11101),
.B1(n_10996),
.B2(n_10963),
.Y(n_11601)
);

INVx4_ASAP7_75t_L g11602 ( 
.A(n_11215),
.Y(n_11602)
);

INVx1_ASAP7_75t_L g11603 ( 
.A(n_11208),
.Y(n_11603)
);

NAND2xp5_ASAP7_75t_L g11604 ( 
.A(n_11435),
.B(n_10659),
.Y(n_11604)
);

BUFx4_ASAP7_75t_R g11605 ( 
.A(n_11466),
.Y(n_11605)
);

INVx2_ASAP7_75t_L g11606 ( 
.A(n_11131),
.Y(n_11606)
);

OAI22xp33_ASAP7_75t_SL g11607 ( 
.A1(n_11370),
.A2(n_10793),
.B1(n_10877),
.B2(n_10816),
.Y(n_11607)
);

HB1xp67_ASAP7_75t_L g11608 ( 
.A(n_11459),
.Y(n_11608)
);

CKINVDCx20_ASAP7_75t_R g11609 ( 
.A(n_11404),
.Y(n_11609)
);

INVx6_ASAP7_75t_L g11610 ( 
.A(n_11477),
.Y(n_11610)
);

OAI22xp33_ASAP7_75t_L g11611 ( 
.A1(n_11311),
.A2(n_10984),
.B1(n_10725),
.B2(n_10864),
.Y(n_11611)
);

INVx4_ASAP7_75t_L g11612 ( 
.A(n_11229),
.Y(n_11612)
);

AOI22xp33_ASAP7_75t_L g11613 ( 
.A1(n_11490),
.A2(n_10966),
.B1(n_10980),
.B2(n_10962),
.Y(n_11613)
);

OAI22xp5_ASAP7_75t_L g11614 ( 
.A1(n_11485),
.A2(n_10984),
.B1(n_10725),
.B2(n_10864),
.Y(n_11614)
);

NAND2xp5_ASAP7_75t_L g11615 ( 
.A(n_11332),
.B(n_10659),
.Y(n_11615)
);

BUFx5_ASAP7_75t_L g11616 ( 
.A(n_11406),
.Y(n_11616)
);

CKINVDCx20_ASAP7_75t_R g11617 ( 
.A(n_11275),
.Y(n_11617)
);

BUFx3_ASAP7_75t_L g11618 ( 
.A(n_11434),
.Y(n_11618)
);

AOI22xp33_ASAP7_75t_SL g11619 ( 
.A1(n_11308),
.A2(n_11117),
.B1(n_11084),
.B2(n_10991),
.Y(n_11619)
);

AOI22xp33_ASAP7_75t_L g11620 ( 
.A1(n_11320),
.A2(n_11084),
.B1(n_11028),
.B2(n_10991),
.Y(n_11620)
);

BUFx12f_ASAP7_75t_L g11621 ( 
.A(n_11475),
.Y(n_11621)
);

BUFx3_ASAP7_75t_L g11622 ( 
.A(n_11433),
.Y(n_11622)
);

OAI22xp33_ASAP7_75t_L g11623 ( 
.A1(n_11329),
.A2(n_10976),
.B1(n_11066),
.B2(n_11109),
.Y(n_11623)
);

OAI22xp5_ASAP7_75t_L g11624 ( 
.A1(n_11400),
.A2(n_10976),
.B1(n_11066),
.B2(n_11109),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_11218),
.Y(n_11625)
);

CKINVDCx20_ASAP7_75t_R g11626 ( 
.A(n_11189),
.Y(n_11626)
);

INVx1_ASAP7_75t_SL g11627 ( 
.A(n_11183),
.Y(n_11627)
);

AOI22xp33_ASAP7_75t_L g11628 ( 
.A1(n_11474),
.A2(n_10888),
.B1(n_10782),
.B2(n_1288),
.Y(n_11628)
);

AOI22xp33_ASAP7_75t_L g11629 ( 
.A1(n_11334),
.A2(n_1292),
.B1(n_1286),
.B2(n_1287),
.Y(n_11629)
);

INVx1_ASAP7_75t_L g11630 ( 
.A(n_11234),
.Y(n_11630)
);

INVx4_ASAP7_75t_L g11631 ( 
.A(n_11229),
.Y(n_11631)
);

BUFx12f_ASAP7_75t_L g11632 ( 
.A(n_11506),
.Y(n_11632)
);

OAI22xp33_ASAP7_75t_L g11633 ( 
.A1(n_11289),
.A2(n_1292),
.B1(n_1286),
.B2(n_1287),
.Y(n_11633)
);

BUFx2_ASAP7_75t_L g11634 ( 
.A(n_11159),
.Y(n_11634)
);

INVx1_ASAP7_75t_SL g11635 ( 
.A(n_11171),
.Y(n_11635)
);

AND2x2_ASAP7_75t_L g11636 ( 
.A(n_11257),
.B(n_1293),
.Y(n_11636)
);

INVx1_ASAP7_75t_SL g11637 ( 
.A(n_11385),
.Y(n_11637)
);

NAND2xp5_ASAP7_75t_L g11638 ( 
.A(n_11333),
.B(n_1293),
.Y(n_11638)
);

INVx2_ASAP7_75t_L g11639 ( 
.A(n_11137),
.Y(n_11639)
);

INVx8_ASAP7_75t_L g11640 ( 
.A(n_11361),
.Y(n_11640)
);

BUFx3_ASAP7_75t_L g11641 ( 
.A(n_11420),
.Y(n_11641)
);

INVx1_ASAP7_75t_L g11642 ( 
.A(n_11235),
.Y(n_11642)
);

CKINVDCx20_ASAP7_75t_R g11643 ( 
.A(n_11421),
.Y(n_11643)
);

BUFx2_ASAP7_75t_L g11644 ( 
.A(n_11252),
.Y(n_11644)
);

INVxp67_ASAP7_75t_SL g11645 ( 
.A(n_11488),
.Y(n_11645)
);

AOI22xp33_ASAP7_75t_L g11646 ( 
.A1(n_11473),
.A2(n_11471),
.B1(n_11461),
.B2(n_11410),
.Y(n_11646)
);

INVx1_ASAP7_75t_SL g11647 ( 
.A(n_11151),
.Y(n_11647)
);

INVx1_ASAP7_75t_L g11648 ( 
.A(n_11274),
.Y(n_11648)
);

AOI22xp33_ASAP7_75t_L g11649 ( 
.A1(n_11411),
.A2(n_1298),
.B1(n_1295),
.B2(n_1297),
.Y(n_11649)
);

NAND2xp5_ASAP7_75t_L g11650 ( 
.A(n_11344),
.B(n_1297),
.Y(n_11650)
);

INVx2_ASAP7_75t_L g11651 ( 
.A(n_11219),
.Y(n_11651)
);

BUFx3_ASAP7_75t_L g11652 ( 
.A(n_11209),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_11156),
.Y(n_11653)
);

AOI22xp33_ASAP7_75t_SL g11654 ( 
.A1(n_11270),
.A2(n_1300),
.B1(n_1298),
.B2(n_1299),
.Y(n_11654)
);

BUFx8_ASAP7_75t_L g11655 ( 
.A(n_11360),
.Y(n_11655)
);

BUFx10_ASAP7_75t_L g11656 ( 
.A(n_11408),
.Y(n_11656)
);

BUFx10_ASAP7_75t_L g11657 ( 
.A(n_11394),
.Y(n_11657)
);

BUFx3_ASAP7_75t_L g11658 ( 
.A(n_11221),
.Y(n_11658)
);

BUFx4f_ASAP7_75t_SL g11659 ( 
.A(n_11343),
.Y(n_11659)
);

INVx1_ASAP7_75t_SL g11660 ( 
.A(n_11302),
.Y(n_11660)
);

AOI22xp33_ASAP7_75t_L g11661 ( 
.A1(n_11383),
.A2(n_1302),
.B1(n_1299),
.B2(n_1301),
.Y(n_11661)
);

BUFx3_ASAP7_75t_L g11662 ( 
.A(n_11254),
.Y(n_11662)
);

BUFx10_ASAP7_75t_L g11663 ( 
.A(n_11340),
.Y(n_11663)
);

BUFx6f_ASAP7_75t_SL g11664 ( 
.A(n_11268),
.Y(n_11664)
);

INVx1_ASAP7_75t_SL g11665 ( 
.A(n_11187),
.Y(n_11665)
);

AOI22xp33_ASAP7_75t_SL g11666 ( 
.A1(n_11352),
.A2(n_1305),
.B1(n_1303),
.B2(n_1304),
.Y(n_11666)
);

BUFx3_ASAP7_75t_L g11667 ( 
.A(n_11264),
.Y(n_11667)
);

INVx4_ASAP7_75t_L g11668 ( 
.A(n_11253),
.Y(n_11668)
);

AOI22xp33_ASAP7_75t_SL g11669 ( 
.A1(n_11504),
.A2(n_1306),
.B1(n_1304),
.B2(n_1305),
.Y(n_11669)
);

BUFx3_ASAP7_75t_L g11670 ( 
.A(n_11182),
.Y(n_11670)
);

INVx4_ASAP7_75t_L g11671 ( 
.A(n_11253),
.Y(n_11671)
);

BUFx2_ASAP7_75t_L g11672 ( 
.A(n_11170),
.Y(n_11672)
);

BUFx6f_ASAP7_75t_L g11673 ( 
.A(n_11278),
.Y(n_11673)
);

INVx1_ASAP7_75t_L g11674 ( 
.A(n_11416),
.Y(n_11674)
);

OAI22xp5_ASAP7_75t_L g11675 ( 
.A1(n_11350),
.A2(n_1308),
.B1(n_1306),
.B2(n_1307),
.Y(n_11675)
);

AOI22xp33_ASAP7_75t_L g11676 ( 
.A1(n_11431),
.A2(n_1309),
.B1(n_1307),
.B2(n_1308),
.Y(n_11676)
);

INVxp67_ASAP7_75t_SL g11677 ( 
.A(n_11346),
.Y(n_11677)
);

INVx6_ASAP7_75t_L g11678 ( 
.A(n_11477),
.Y(n_11678)
);

INVx4_ASAP7_75t_L g11679 ( 
.A(n_11278),
.Y(n_11679)
);

AOI22xp5_ASAP7_75t_L g11680 ( 
.A1(n_11453),
.A2(n_1311),
.B1(n_1309),
.B2(n_1310),
.Y(n_11680)
);

INVx2_ASAP7_75t_L g11681 ( 
.A(n_11220),
.Y(n_11681)
);

AND2x2_ASAP7_75t_L g11682 ( 
.A(n_11307),
.B(n_1310),
.Y(n_11682)
);

OAI22xp5_ASAP7_75t_L g11683 ( 
.A1(n_11145),
.A2(n_1313),
.B1(n_1311),
.B2(n_1312),
.Y(n_11683)
);

INVx1_ASAP7_75t_L g11684 ( 
.A(n_11417),
.Y(n_11684)
);

INVx1_ASAP7_75t_L g11685 ( 
.A(n_11429),
.Y(n_11685)
);

INVx2_ASAP7_75t_L g11686 ( 
.A(n_11322),
.Y(n_11686)
);

AOI22xp33_ASAP7_75t_L g11687 ( 
.A1(n_11458),
.A2(n_11436),
.B1(n_11224),
.B2(n_11444),
.Y(n_11687)
);

AOI22xp33_ASAP7_75t_L g11688 ( 
.A1(n_11441),
.A2(n_1314),
.B1(n_1312),
.B2(n_1313),
.Y(n_11688)
);

AOI22xp33_ASAP7_75t_L g11689 ( 
.A1(n_11443),
.A2(n_11445),
.B1(n_11499),
.B2(n_11493),
.Y(n_11689)
);

AOI22xp33_ASAP7_75t_L g11690 ( 
.A1(n_11310),
.A2(n_11225),
.B1(n_11168),
.B2(n_11169),
.Y(n_11690)
);

AOI22xp33_ASAP7_75t_SL g11691 ( 
.A1(n_11300),
.A2(n_1316),
.B1(n_1314),
.B2(n_1315),
.Y(n_11691)
);

NAND2xp5_ASAP7_75t_L g11692 ( 
.A(n_11355),
.B(n_1316),
.Y(n_11692)
);

BUFx12f_ASAP7_75t_L g11693 ( 
.A(n_11391),
.Y(n_11693)
);

INVx1_ASAP7_75t_L g11694 ( 
.A(n_11240),
.Y(n_11694)
);

AOI22xp33_ASAP7_75t_SL g11695 ( 
.A1(n_11395),
.A2(n_1319),
.B1(n_1317),
.B2(n_1318),
.Y(n_11695)
);

CKINVDCx11_ASAP7_75t_R g11696 ( 
.A(n_11317),
.Y(n_11696)
);

INVx4_ASAP7_75t_L g11697 ( 
.A(n_11317),
.Y(n_11697)
);

INVx1_ASAP7_75t_SL g11698 ( 
.A(n_11144),
.Y(n_11698)
);

BUFx6f_ASAP7_75t_L g11699 ( 
.A(n_11327),
.Y(n_11699)
);

NAND2xp5_ASAP7_75t_L g11700 ( 
.A(n_11356),
.B(n_11366),
.Y(n_11700)
);

OR2x2_ASAP7_75t_L g11701 ( 
.A(n_11297),
.B(n_1317),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_11249),
.Y(n_11702)
);

OAI22xp5_ASAP7_75t_L g11703 ( 
.A1(n_11377),
.A2(n_1320),
.B1(n_1318),
.B2(n_1319),
.Y(n_11703)
);

INVx11_ASAP7_75t_L g11704 ( 
.A(n_11419),
.Y(n_11704)
);

BUFx6f_ASAP7_75t_L g11705 ( 
.A(n_11327),
.Y(n_11705)
);

AOI22xp33_ASAP7_75t_SL g11706 ( 
.A1(n_11472),
.A2(n_11500),
.B1(n_11203),
.B2(n_11349),
.Y(n_11706)
);

CKINVDCx5p33_ASAP7_75t_R g11707 ( 
.A(n_11347),
.Y(n_11707)
);

BUFx3_ASAP7_75t_L g11708 ( 
.A(n_11134),
.Y(n_11708)
);

INVx1_ASAP7_75t_L g11709 ( 
.A(n_11260),
.Y(n_11709)
);

OAI22xp5_ASAP7_75t_L g11710 ( 
.A1(n_11291),
.A2(n_11367),
.B1(n_11336),
.B2(n_11426),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_11269),
.Y(n_11711)
);

BUFx10_ASAP7_75t_L g11712 ( 
.A(n_11280),
.Y(n_11712)
);

INVx2_ASAP7_75t_L g11713 ( 
.A(n_11324),
.Y(n_11713)
);

INVx2_ASAP7_75t_L g11714 ( 
.A(n_11272),
.Y(n_11714)
);

INVx1_ASAP7_75t_L g11715 ( 
.A(n_11279),
.Y(n_11715)
);

INVx1_ASAP7_75t_L g11716 ( 
.A(n_11301),
.Y(n_11716)
);

INVx2_ASAP7_75t_L g11717 ( 
.A(n_11199),
.Y(n_11717)
);

OAI22xp33_ASAP7_75t_L g11718 ( 
.A1(n_11373),
.A2(n_1324),
.B1(n_1322),
.B2(n_1323),
.Y(n_11718)
);

BUFx12f_ASAP7_75t_L g11719 ( 
.A(n_11372),
.Y(n_11719)
);

INVx1_ASAP7_75t_L g11720 ( 
.A(n_11315),
.Y(n_11720)
);

OAI22xp5_ASAP7_75t_L g11721 ( 
.A1(n_11267),
.A2(n_1325),
.B1(n_1322),
.B2(n_1323),
.Y(n_11721)
);

OAI22xp5_ASAP7_75t_L g11722 ( 
.A1(n_11439),
.A2(n_1328),
.B1(n_1325),
.B2(n_1327),
.Y(n_11722)
);

CKINVDCx5p33_ASAP7_75t_R g11723 ( 
.A(n_11347),
.Y(n_11723)
);

BUFx2_ASAP7_75t_L g11724 ( 
.A(n_11223),
.Y(n_11724)
);

OAI22xp5_ASAP7_75t_L g11725 ( 
.A1(n_11413),
.A2(n_1329),
.B1(n_1327),
.B2(n_1328),
.Y(n_11725)
);

CKINVDCx5p33_ASAP7_75t_R g11726 ( 
.A(n_11368),
.Y(n_11726)
);

INVx3_ASAP7_75t_L g11727 ( 
.A(n_11374),
.Y(n_11727)
);

AOI22xp33_ASAP7_75t_L g11728 ( 
.A1(n_11379),
.A2(n_1332),
.B1(n_1330),
.B2(n_1331),
.Y(n_11728)
);

NAND2xp5_ASAP7_75t_L g11729 ( 
.A(n_11371),
.B(n_1330),
.Y(n_11729)
);

INVx2_ASAP7_75t_SL g11730 ( 
.A(n_11132),
.Y(n_11730)
);

BUFx4f_ASAP7_75t_SL g11731 ( 
.A(n_11368),
.Y(n_11731)
);

BUFx8_ASAP7_75t_L g11732 ( 
.A(n_11418),
.Y(n_11732)
);

AOI22xp5_ASAP7_75t_L g11733 ( 
.A1(n_11401),
.A2(n_1333),
.B1(n_1331),
.B2(n_1332),
.Y(n_11733)
);

HB1xp67_ASAP7_75t_L g11734 ( 
.A(n_11467),
.Y(n_11734)
);

CKINVDCx5p33_ASAP7_75t_R g11735 ( 
.A(n_11409),
.Y(n_11735)
);

INVx4_ASAP7_75t_L g11736 ( 
.A(n_11409),
.Y(n_11736)
);

AOI22xp33_ASAP7_75t_L g11737 ( 
.A1(n_11469),
.A2(n_1335),
.B1(n_1333),
.B2(n_1334),
.Y(n_11737)
);

AOI22xp33_ASAP7_75t_L g11738 ( 
.A1(n_11482),
.A2(n_1336),
.B1(n_1334),
.B2(n_1335),
.Y(n_11738)
);

CKINVDCx20_ASAP7_75t_R g11739 ( 
.A(n_11290),
.Y(n_11739)
);

AOI22xp33_ASAP7_75t_L g11740 ( 
.A1(n_11496),
.A2(n_1339),
.B1(n_1336),
.B2(n_1337),
.Y(n_11740)
);

INVx1_ASAP7_75t_L g11741 ( 
.A(n_11180),
.Y(n_11741)
);

INVx1_ASAP7_75t_L g11742 ( 
.A(n_11259),
.Y(n_11742)
);

BUFx2_ASAP7_75t_L g11743 ( 
.A(n_11133),
.Y(n_11743)
);

BUFx12f_ASAP7_75t_L g11744 ( 
.A(n_11365),
.Y(n_11744)
);

INVx6_ASAP7_75t_L g11745 ( 
.A(n_11412),
.Y(n_11745)
);

INVx5_ASAP7_75t_L g11746 ( 
.A(n_11478),
.Y(n_11746)
);

INVx2_ASAP7_75t_L g11747 ( 
.A(n_11285),
.Y(n_11747)
);

CKINVDCx20_ASAP7_75t_R g11748 ( 
.A(n_11258),
.Y(n_11748)
);

AOI22xp33_ASAP7_75t_L g11749 ( 
.A1(n_11505),
.A2(n_1341),
.B1(n_1339),
.B2(n_1340),
.Y(n_11749)
);

BUFx10_ASAP7_75t_L g11750 ( 
.A(n_11263),
.Y(n_11750)
);

INVx2_ASAP7_75t_L g11751 ( 
.A(n_11233),
.Y(n_11751)
);

AOI22xp33_ASAP7_75t_L g11752 ( 
.A1(n_11462),
.A2(n_1343),
.B1(n_1340),
.B2(n_1342),
.Y(n_11752)
);

AOI22xp33_ASAP7_75t_L g11753 ( 
.A1(n_11463),
.A2(n_1346),
.B1(n_1343),
.B2(n_1345),
.Y(n_11753)
);

BUFx2_ASAP7_75t_L g11754 ( 
.A(n_11147),
.Y(n_11754)
);

BUFx12f_ASAP7_75t_L g11755 ( 
.A(n_11442),
.Y(n_11755)
);

AOI22xp33_ASAP7_75t_L g11756 ( 
.A1(n_11386),
.A2(n_1347),
.B1(n_1345),
.B2(n_1346),
.Y(n_11756)
);

BUFx3_ASAP7_75t_L g11757 ( 
.A(n_11138),
.Y(n_11757)
);

CKINVDCx5p33_ASAP7_75t_R g11758 ( 
.A(n_11412),
.Y(n_11758)
);

INVx2_ASAP7_75t_L g11759 ( 
.A(n_11241),
.Y(n_11759)
);

BUFx3_ASAP7_75t_L g11760 ( 
.A(n_11337),
.Y(n_11760)
);

AOI22xp33_ASAP7_75t_L g11761 ( 
.A1(n_11497),
.A2(n_1349),
.B1(n_1347),
.B2(n_1348),
.Y(n_11761)
);

INVx1_ASAP7_75t_L g11762 ( 
.A(n_11282),
.Y(n_11762)
);

AOI22xp33_ASAP7_75t_L g11763 ( 
.A1(n_11452),
.A2(n_1350),
.B1(n_1348),
.B2(n_1349),
.Y(n_11763)
);

OAI22xp33_ASAP7_75t_L g11764 ( 
.A1(n_11217),
.A2(n_1353),
.B1(n_1351),
.B2(n_1352),
.Y(n_11764)
);

BUFx2_ASAP7_75t_L g11765 ( 
.A(n_11422),
.Y(n_11765)
);

AOI22xp33_ASAP7_75t_L g11766 ( 
.A1(n_11464),
.A2(n_11481),
.B1(n_11468),
.B2(n_11236),
.Y(n_11766)
);

OAI22xp5_ASAP7_75t_L g11767 ( 
.A1(n_11375),
.A2(n_1354),
.B1(n_1352),
.B2(n_1353),
.Y(n_11767)
);

AOI22xp33_ASAP7_75t_L g11768 ( 
.A1(n_11284),
.A2(n_1356),
.B1(n_1354),
.B2(n_1355),
.Y(n_11768)
);

AOI22xp33_ASAP7_75t_L g11769 ( 
.A1(n_11286),
.A2(n_1357),
.B1(n_1355),
.B2(n_1356),
.Y(n_11769)
);

INVx1_ASAP7_75t_L g11770 ( 
.A(n_11312),
.Y(n_11770)
);

INVx1_ASAP7_75t_L g11771 ( 
.A(n_11460),
.Y(n_11771)
);

BUFx8_ASAP7_75t_L g11772 ( 
.A(n_11440),
.Y(n_11772)
);

AOI22xp33_ASAP7_75t_L g11773 ( 
.A1(n_11230),
.A2(n_1359),
.B1(n_1357),
.B2(n_1358),
.Y(n_11773)
);

CKINVDCx20_ASAP7_75t_R g11774 ( 
.A(n_11175),
.Y(n_11774)
);

INVx2_ASAP7_75t_L g11775 ( 
.A(n_11207),
.Y(n_11775)
);

CKINVDCx11_ASAP7_75t_R g11776 ( 
.A(n_11296),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_11465),
.Y(n_11777)
);

BUFx6f_ASAP7_75t_L g11778 ( 
.A(n_11442),
.Y(n_11778)
);

OAI22xp5_ASAP7_75t_L g11779 ( 
.A1(n_11261),
.A2(n_1360),
.B1(n_1358),
.B2(n_1359),
.Y(n_11779)
);

AOI22xp33_ASAP7_75t_L g11780 ( 
.A1(n_11358),
.A2(n_1363),
.B1(n_1360),
.B2(n_1361),
.Y(n_11780)
);

INVx1_ASAP7_75t_L g11781 ( 
.A(n_11364),
.Y(n_11781)
);

OAI22xp5_ASAP7_75t_L g11782 ( 
.A1(n_11338),
.A2(n_1364),
.B1(n_1361),
.B2(n_1363),
.Y(n_11782)
);

OAI22xp33_ASAP7_75t_L g11783 ( 
.A1(n_11162),
.A2(n_1366),
.B1(n_1364),
.B2(n_1365),
.Y(n_11783)
);

OAI22xp33_ASAP7_75t_L g11784 ( 
.A1(n_11283),
.A2(n_1368),
.B1(n_1366),
.B2(n_1367),
.Y(n_11784)
);

INVx2_ASAP7_75t_L g11785 ( 
.A(n_11205),
.Y(n_11785)
);

OAI22xp33_ASAP7_75t_L g11786 ( 
.A1(n_11184),
.A2(n_1370),
.B1(n_1367),
.B2(n_1369),
.Y(n_11786)
);

NAND2xp5_ASAP7_75t_L g11787 ( 
.A(n_11381),
.B(n_1369),
.Y(n_11787)
);

AND2x2_ASAP7_75t_L g11788 ( 
.A(n_11190),
.B(n_11342),
.Y(n_11788)
);

CKINVDCx11_ASAP7_75t_R g11789 ( 
.A(n_11425),
.Y(n_11789)
);

OAI22xp33_ASAP7_75t_L g11790 ( 
.A1(n_11195),
.A2(n_1372),
.B1(n_1370),
.B2(n_1371),
.Y(n_11790)
);

INVx2_ASAP7_75t_L g11791 ( 
.A(n_11266),
.Y(n_11791)
);

CKINVDCx11_ASAP7_75t_R g11792 ( 
.A(n_11476),
.Y(n_11792)
);

OAI21xp33_ASAP7_75t_L g11793 ( 
.A1(n_11450),
.A2(n_1371),
.B(n_1372),
.Y(n_11793)
);

OAI22xp5_ASAP7_75t_SL g11794 ( 
.A1(n_11153),
.A2(n_1375),
.B1(n_1373),
.B2(n_1374),
.Y(n_11794)
);

CKINVDCx5p33_ASAP7_75t_R g11795 ( 
.A(n_11214),
.Y(n_11795)
);

CKINVDCx11_ASAP7_75t_R g11796 ( 
.A(n_11398),
.Y(n_11796)
);

INVx1_ASAP7_75t_L g11797 ( 
.A(n_11163),
.Y(n_11797)
);

INVx1_ASAP7_75t_L g11798 ( 
.A(n_11403),
.Y(n_11798)
);

INVx2_ASAP7_75t_L g11799 ( 
.A(n_11428),
.Y(n_11799)
);

BUFx2_ASAP7_75t_L g11800 ( 
.A(n_11423),
.Y(n_11800)
);

OAI22xp5_ASAP7_75t_L g11801 ( 
.A1(n_11242),
.A2(n_1376),
.B1(n_1373),
.B2(n_1375),
.Y(n_11801)
);

AOI22xp33_ASAP7_75t_L g11802 ( 
.A1(n_11339),
.A2(n_11480),
.B1(n_11446),
.B2(n_11405),
.Y(n_11802)
);

BUFx10_ASAP7_75t_L g11803 ( 
.A(n_11239),
.Y(n_11803)
);

INVx2_ASAP7_75t_L g11804 ( 
.A(n_11438),
.Y(n_11804)
);

BUFx8_ASAP7_75t_L g11805 ( 
.A(n_11495),
.Y(n_11805)
);

OAI22xp33_ASAP7_75t_L g11806 ( 
.A1(n_11309),
.A2(n_1378),
.B1(n_1376),
.B2(n_1377),
.Y(n_11806)
);

CKINVDCx20_ASAP7_75t_R g11807 ( 
.A(n_11256),
.Y(n_11807)
);

INVx2_ASAP7_75t_L g11808 ( 
.A(n_11271),
.Y(n_11808)
);

BUFx8_ASAP7_75t_L g11809 ( 
.A(n_11503),
.Y(n_11809)
);

CKINVDCx11_ASAP7_75t_R g11810 ( 
.A(n_11357),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_11427),
.Y(n_11811)
);

INVx2_ASAP7_75t_L g11812 ( 
.A(n_11201),
.Y(n_11812)
);

OAI22xp33_ASAP7_75t_L g11813 ( 
.A1(n_11238),
.A2(n_1381),
.B1(n_1378),
.B2(n_1379),
.Y(n_11813)
);

BUFx2_ASAP7_75t_SL g11814 ( 
.A(n_11293),
.Y(n_11814)
);

AOI22xp5_ASAP7_75t_L g11815 ( 
.A1(n_11277),
.A2(n_1383),
.B1(n_1381),
.B2(n_1382),
.Y(n_11815)
);

AOI22xp33_ASAP7_75t_L g11816 ( 
.A1(n_11456),
.A2(n_1386),
.B1(n_1384),
.B2(n_1385),
.Y(n_11816)
);

AOI22xp33_ASAP7_75t_L g11817 ( 
.A1(n_11491),
.A2(n_1386),
.B1(n_1384),
.B2(n_1385),
.Y(n_11817)
);

AOI22xp33_ASAP7_75t_L g11818 ( 
.A1(n_11228),
.A2(n_1389),
.B1(n_1387),
.B2(n_1388),
.Y(n_11818)
);

INVx2_ASAP7_75t_L g11819 ( 
.A(n_11380),
.Y(n_11819)
);

INVxp67_ASAP7_75t_SL g11820 ( 
.A(n_11142),
.Y(n_11820)
);

AOI22xp33_ASAP7_75t_L g11821 ( 
.A1(n_11139),
.A2(n_1391),
.B1(n_1388),
.B2(n_1390),
.Y(n_11821)
);

INVx3_ASAP7_75t_L g11822 ( 
.A(n_11299),
.Y(n_11822)
);

AOI22xp33_ASAP7_75t_L g11823 ( 
.A1(n_11354),
.A2(n_1392),
.B1(n_1390),
.B2(n_1391),
.Y(n_11823)
);

AOI22xp33_ASAP7_75t_L g11824 ( 
.A1(n_11507),
.A2(n_1394),
.B1(n_1392),
.B2(n_1393),
.Y(n_11824)
);

BUFx3_ASAP7_75t_L g11825 ( 
.A(n_11348),
.Y(n_11825)
);

AOI22xp33_ASAP7_75t_L g11826 ( 
.A1(n_11455),
.A2(n_1395),
.B1(n_1393),
.B2(n_1394),
.Y(n_11826)
);

OAI22xp5_ASAP7_75t_L g11827 ( 
.A1(n_11292),
.A2(n_1397),
.B1(n_1395),
.B2(n_1396),
.Y(n_11827)
);

CKINVDCx11_ASAP7_75t_R g11828 ( 
.A(n_11397),
.Y(n_11828)
);

AOI22xp33_ASAP7_75t_L g11829 ( 
.A1(n_11143),
.A2(n_1399),
.B1(n_1397),
.B2(n_1398),
.Y(n_11829)
);

NAND2x1p5_ASAP7_75t_L g11830 ( 
.A(n_11437),
.B(n_1399),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_11213),
.B(n_1400),
.Y(n_11831)
);

AND2x2_ASAP7_75t_L g11832 ( 
.A(n_11186),
.B(n_1400),
.Y(n_11832)
);

BUFx8_ASAP7_75t_L g11833 ( 
.A(n_11389),
.Y(n_11833)
);

INVx1_ASAP7_75t_L g11834 ( 
.A(n_11231),
.Y(n_11834)
);

AOI22xp33_ASAP7_75t_L g11835 ( 
.A1(n_11167),
.A2(n_1403),
.B1(n_1401),
.B2(n_1402),
.Y(n_11835)
);

INVx2_ASAP7_75t_L g11836 ( 
.A(n_11255),
.Y(n_11836)
);

OAI21xp5_ASAP7_75t_L g11837 ( 
.A1(n_11328),
.A2(n_1401),
.B(n_1403),
.Y(n_11837)
);

CKINVDCx20_ASAP7_75t_R g11838 ( 
.A(n_11164),
.Y(n_11838)
);

NAND2xp5_ASAP7_75t_L g11839 ( 
.A(n_11232),
.B(n_1404),
.Y(n_11839)
);

BUFx12f_ASAP7_75t_L g11840 ( 
.A(n_11402),
.Y(n_11840)
);

AOI22xp33_ASAP7_75t_L g11841 ( 
.A1(n_11287),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_11841)
);

AOI22xp33_ASAP7_75t_L g11842 ( 
.A1(n_11244),
.A2(n_1407),
.B1(n_1405),
.B2(n_1406),
.Y(n_11842)
);

INVx6_ASAP7_75t_L g11843 ( 
.A(n_11250),
.Y(n_11843)
);

INVx2_ASAP7_75t_L g11844 ( 
.A(n_11616),
.Y(n_11844)
);

NAND2xp5_ASAP7_75t_L g11845 ( 
.A(n_11820),
.B(n_11295),
.Y(n_11845)
);

INVx2_ASAP7_75t_SL g11846 ( 
.A(n_11514),
.Y(n_11846)
);

AOI22xp33_ASAP7_75t_L g11847 ( 
.A1(n_11833),
.A2(n_11393),
.B1(n_11335),
.B2(n_11479),
.Y(n_11847)
);

OAI21x1_ASAP7_75t_L g11848 ( 
.A1(n_11812),
.A2(n_11508),
.B(n_11771),
.Y(n_11848)
);

AOI22xp33_ASAP7_75t_L g11849 ( 
.A1(n_11579),
.A2(n_11568),
.B1(n_11545),
.B2(n_11690),
.Y(n_11849)
);

CKINVDCx9p33_ASAP7_75t_R g11850 ( 
.A(n_11565),
.Y(n_11850)
);

AND2x2_ASAP7_75t_L g11851 ( 
.A(n_11634),
.B(n_11814),
.Y(n_11851)
);

BUFx3_ASAP7_75t_L g11852 ( 
.A(n_11510),
.Y(n_11852)
);

OR2x6_ASAP7_75t_L g11853 ( 
.A(n_11520),
.B(n_11407),
.Y(n_11853)
);

BUFx3_ASAP7_75t_L g11854 ( 
.A(n_11509),
.Y(n_11854)
);

BUFx6f_ASAP7_75t_L g11855 ( 
.A(n_11567),
.Y(n_11855)
);

INVx1_ASAP7_75t_L g11856 ( 
.A(n_11674),
.Y(n_11856)
);

NAND2x1p5_ASAP7_75t_L g11857 ( 
.A(n_11627),
.B(n_11304),
.Y(n_11857)
);

OAI22xp5_ASAP7_75t_SL g11858 ( 
.A1(n_11511),
.A2(n_11378),
.B1(n_11351),
.B2(n_11501),
.Y(n_11858)
);

AND2x2_ASAP7_75t_L g11859 ( 
.A(n_11746),
.B(n_11251),
.Y(n_11859)
);

AOI21x1_ASAP7_75t_L g11860 ( 
.A1(n_11724),
.A2(n_11487),
.B(n_11387),
.Y(n_11860)
);

BUFx6f_ASAP7_75t_L g11861 ( 
.A(n_11514),
.Y(n_11861)
);

INVx2_ASAP7_75t_L g11862 ( 
.A(n_11616),
.Y(n_11862)
);

NAND2xp33_ASAP7_75t_R g11863 ( 
.A(n_11556),
.B(n_11449),
.Y(n_11863)
);

INVx1_ASAP7_75t_L g11864 ( 
.A(n_11684),
.Y(n_11864)
);

HB1xp67_ASAP7_75t_L g11865 ( 
.A(n_11553),
.Y(n_11865)
);

BUFx2_ASAP7_75t_L g11866 ( 
.A(n_11617),
.Y(n_11866)
);

OAI21xp5_ASAP7_75t_L g11867 ( 
.A1(n_11580),
.A2(n_11396),
.B(n_11454),
.Y(n_11867)
);

INVx1_ASAP7_75t_L g11868 ( 
.A(n_11685),
.Y(n_11868)
);

OAI21x1_ASAP7_75t_L g11869 ( 
.A1(n_11777),
.A2(n_11246),
.B(n_11251),
.Y(n_11869)
);

OAI22xp5_ASAP7_75t_L g11870 ( 
.A1(n_11687),
.A2(n_11246),
.B1(n_11389),
.B2(n_1409),
.Y(n_11870)
);

AOI221xp5_ASAP7_75t_L g11871 ( 
.A1(n_11595),
.A2(n_1410),
.B1(n_1407),
.B2(n_1408),
.C(n_1411),
.Y(n_11871)
);

AOI22xp33_ASAP7_75t_L g11872 ( 
.A1(n_11534),
.A2(n_1412),
.B1(n_1408),
.B2(n_1410),
.Y(n_11872)
);

NOR2xp33_ASAP7_75t_L g11873 ( 
.A(n_11527),
.B(n_1412),
.Y(n_11873)
);

AND2x4_ASAP7_75t_L g11874 ( 
.A(n_11516),
.B(n_1413),
.Y(n_11874)
);

BUFx8_ASAP7_75t_SL g11875 ( 
.A(n_11581),
.Y(n_11875)
);

AOI21xp5_ASAP7_75t_L g11876 ( 
.A1(n_11533),
.A2(n_1414),
.B(n_1415),
.Y(n_11876)
);

AOI22xp5_ASAP7_75t_L g11877 ( 
.A1(n_11528),
.A2(n_1416),
.B1(n_1414),
.B2(n_1415),
.Y(n_11877)
);

NAND2xp5_ASAP7_75t_L g11878 ( 
.A(n_11677),
.B(n_11797),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11521),
.Y(n_11879)
);

AOI221xp5_ASAP7_75t_L g11880 ( 
.A1(n_11683),
.A2(n_11703),
.B1(n_11721),
.B2(n_11607),
.C(n_11710),
.Y(n_11880)
);

HB1xp67_ASAP7_75t_L g11881 ( 
.A(n_11608),
.Y(n_11881)
);

INVx2_ASAP7_75t_L g11882 ( 
.A(n_11616),
.Y(n_11882)
);

INVx3_ASAP7_75t_L g11883 ( 
.A(n_11518),
.Y(n_11883)
);

INVx1_ASAP7_75t_L g11884 ( 
.A(n_11522),
.Y(n_11884)
);

OAI22xp5_ASAP7_75t_SL g11885 ( 
.A1(n_11523),
.A2(n_1418),
.B1(n_1416),
.B2(n_1417),
.Y(n_11885)
);

NAND2xp5_ASAP7_75t_L g11886 ( 
.A(n_11519),
.B(n_1419),
.Y(n_11886)
);

OAI21x1_ASAP7_75t_L g11887 ( 
.A1(n_11615),
.A2(n_1420),
.B(n_1421),
.Y(n_11887)
);

NOR2xp33_ASAP7_75t_R g11888 ( 
.A(n_11609),
.B(n_1420),
.Y(n_11888)
);

AND2x2_ASAP7_75t_L g11889 ( 
.A(n_11746),
.B(n_1421),
.Y(n_11889)
);

INVx2_ASAP7_75t_SL g11890 ( 
.A(n_11704),
.Y(n_11890)
);

BUFx4f_ASAP7_75t_L g11891 ( 
.A(n_11524),
.Y(n_11891)
);

OAI22xp33_ASAP7_75t_L g11892 ( 
.A1(n_11571),
.A2(n_1424),
.B1(n_1422),
.B2(n_1423),
.Y(n_11892)
);

BUFx6f_ASAP7_75t_L g11893 ( 
.A(n_11541),
.Y(n_11893)
);

OAI22xp5_ASAP7_75t_L g11894 ( 
.A1(n_11706),
.A2(n_1425),
.B1(n_1422),
.B2(n_1424),
.Y(n_11894)
);

INVx3_ASAP7_75t_L g11895 ( 
.A(n_11712),
.Y(n_11895)
);

INVx3_ASAP7_75t_L g11896 ( 
.A(n_11538),
.Y(n_11896)
);

AOI22xp33_ASAP7_75t_L g11897 ( 
.A1(n_11535),
.A2(n_1427),
.B1(n_1425),
.B2(n_1426),
.Y(n_11897)
);

AND2x4_ASAP7_75t_L g11898 ( 
.A(n_11573),
.B(n_1426),
.Y(n_11898)
);

AND2x2_ASAP7_75t_L g11899 ( 
.A(n_11765),
.B(n_1427),
.Y(n_11899)
);

INVx3_ASAP7_75t_L g11900 ( 
.A(n_11538),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_11526),
.Y(n_11901)
);

AND2x4_ASAP7_75t_L g11902 ( 
.A(n_11727),
.B(n_1428),
.Y(n_11902)
);

OAI22xp33_ASAP7_75t_L g11903 ( 
.A1(n_11614),
.A2(n_1430),
.B1(n_1428),
.B2(n_1429),
.Y(n_11903)
);

OAI22xp5_ASAP7_75t_L g11904 ( 
.A1(n_11766),
.A2(n_1432),
.B1(n_1430),
.B2(n_1431),
.Y(n_11904)
);

INVx6_ASAP7_75t_L g11905 ( 
.A(n_11587),
.Y(n_11905)
);

OAI21xp5_ASAP7_75t_L g11906 ( 
.A1(n_11550),
.A2(n_1431),
.B(n_1433),
.Y(n_11906)
);

INVx1_ASAP7_75t_L g11907 ( 
.A(n_11530),
.Y(n_11907)
);

AOI22xp33_ASAP7_75t_L g11908 ( 
.A1(n_11531),
.A2(n_1435),
.B1(n_1433),
.B2(n_1434),
.Y(n_11908)
);

BUFx4f_ASAP7_75t_L g11909 ( 
.A(n_11576),
.Y(n_11909)
);

INVx1_ASAP7_75t_L g11910 ( 
.A(n_11542),
.Y(n_11910)
);

OAI22xp5_ASAP7_75t_L g11911 ( 
.A1(n_11620),
.A2(n_1437),
.B1(n_1435),
.B2(n_1436),
.Y(n_11911)
);

CKINVDCx5p33_ASAP7_75t_R g11912 ( 
.A(n_11515),
.Y(n_11912)
);

AOI22xp33_ASAP7_75t_SL g11913 ( 
.A1(n_11549),
.A2(n_1438),
.B1(n_1436),
.B2(n_1437),
.Y(n_11913)
);

OR2x2_ASAP7_75t_L g11914 ( 
.A(n_11604),
.B(n_1438),
.Y(n_11914)
);

AOI22xp33_ASAP7_75t_L g11915 ( 
.A1(n_11794),
.A2(n_11558),
.B1(n_11548),
.B2(n_11767),
.Y(n_11915)
);

AO21x2_ASAP7_75t_L g11916 ( 
.A1(n_11540),
.A2(n_1439),
.B(n_1440),
.Y(n_11916)
);

INVx1_ASAP7_75t_L g11917 ( 
.A(n_11546),
.Y(n_11917)
);

AND2x2_ASAP7_75t_L g11918 ( 
.A(n_11800),
.B(n_1439),
.Y(n_11918)
);

CKINVDCx20_ASAP7_75t_R g11919 ( 
.A(n_11626),
.Y(n_11919)
);

AOI22xp33_ASAP7_75t_L g11920 ( 
.A1(n_11544),
.A2(n_1442),
.B1(n_1440),
.B2(n_1441),
.Y(n_11920)
);

AOI22xp33_ASAP7_75t_L g11921 ( 
.A1(n_11827),
.A2(n_1445),
.B1(n_1442),
.B2(n_1444),
.Y(n_11921)
);

NAND2xp5_ASAP7_75t_L g11922 ( 
.A(n_11781),
.B(n_1445),
.Y(n_11922)
);

INVx1_ASAP7_75t_L g11923 ( 
.A(n_11555),
.Y(n_11923)
);

NAND2xp5_ASAP7_75t_L g11924 ( 
.A(n_11834),
.B(n_11741),
.Y(n_11924)
);

OAI221xp5_ASAP7_75t_L g11925 ( 
.A1(n_11646),
.A2(n_1449),
.B1(n_1446),
.B2(n_1448),
.C(n_1450),
.Y(n_11925)
);

NAND3xp33_ASAP7_75t_SL g11926 ( 
.A(n_11619),
.B(n_11837),
.C(n_11547),
.Y(n_11926)
);

INVx2_ASAP7_75t_L g11927 ( 
.A(n_11616),
.Y(n_11927)
);

BUFx4_ASAP7_75t_SL g11928 ( 
.A(n_11574),
.Y(n_11928)
);

AND2x2_ASAP7_75t_L g11929 ( 
.A(n_11660),
.B(n_1446),
.Y(n_11929)
);

AOI22xp33_ASAP7_75t_L g11930 ( 
.A1(n_11560),
.A2(n_1451),
.B1(n_1449),
.B2(n_1450),
.Y(n_11930)
);

INVx1_ASAP7_75t_L g11931 ( 
.A(n_11564),
.Y(n_11931)
);

AND2x4_ASAP7_75t_L g11932 ( 
.A(n_11672),
.B(n_1451),
.Y(n_11932)
);

INVx4_ASAP7_75t_L g11933 ( 
.A(n_11587),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11570),
.Y(n_11934)
);

INVx2_ASAP7_75t_L g11935 ( 
.A(n_11537),
.Y(n_11935)
);

OR2x6_ASAP7_75t_L g11936 ( 
.A(n_11755),
.B(n_1452),
.Y(n_11936)
);

AOI22xp5_ASAP7_75t_L g11937 ( 
.A1(n_11624),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_11937)
);

OA21x2_ASAP7_75t_L g11938 ( 
.A1(n_11644),
.A2(n_1453),
.B(n_1454),
.Y(n_11938)
);

OAI22xp5_ASAP7_75t_L g11939 ( 
.A1(n_11601),
.A2(n_1457),
.B1(n_1455),
.B2(n_1456),
.Y(n_11939)
);

AND2x4_ASAP7_75t_L g11940 ( 
.A(n_11667),
.B(n_1455),
.Y(n_11940)
);

INVx2_ASAP7_75t_L g11941 ( 
.A(n_11747),
.Y(n_11941)
);

BUFx12f_ASAP7_75t_L g11942 ( 
.A(n_11696),
.Y(n_11942)
);

OAI22xp33_ASAP7_75t_L g11943 ( 
.A1(n_11659),
.A2(n_1462),
.B1(n_1459),
.B2(n_1461),
.Y(n_11943)
);

NAND2xp5_ASAP7_75t_L g11944 ( 
.A(n_11742),
.B(n_11653),
.Y(n_11944)
);

NOR2xp33_ASAP7_75t_L g11945 ( 
.A(n_11512),
.B(n_1459),
.Y(n_11945)
);

INVx1_ASAP7_75t_L g11946 ( 
.A(n_11603),
.Y(n_11946)
);

NAND2xp5_ASAP7_75t_SL g11947 ( 
.A(n_11647),
.B(n_1461),
.Y(n_11947)
);

AOI21xp5_ASAP7_75t_L g11948 ( 
.A1(n_11623),
.A2(n_1462),
.B(n_1463),
.Y(n_11948)
);

BUFx10_ASAP7_75t_L g11949 ( 
.A(n_11664),
.Y(n_11949)
);

OR2x2_ASAP7_75t_L g11950 ( 
.A(n_11552),
.B(n_11754),
.Y(n_11950)
);

OA21x2_ASAP7_75t_L g11951 ( 
.A1(n_11645),
.A2(n_1463),
.B(n_1464),
.Y(n_11951)
);

OAI22xp5_ASAP7_75t_L g11952 ( 
.A1(n_11689),
.A2(n_1466),
.B1(n_1464),
.B2(n_1465),
.Y(n_11952)
);

INVx2_ASAP7_75t_L g11953 ( 
.A(n_11686),
.Y(n_11953)
);

AOI21xp33_ASAP7_75t_SL g11954 ( 
.A1(n_11784),
.A2(n_11830),
.B(n_11764),
.Y(n_11954)
);

NAND2xp5_ASAP7_75t_L g11955 ( 
.A(n_11802),
.B(n_1465),
.Y(n_11955)
);

INVx1_ASAP7_75t_L g11956 ( 
.A(n_11625),
.Y(n_11956)
);

INVx1_ASAP7_75t_L g11957 ( 
.A(n_11630),
.Y(n_11957)
);

OAI21x1_ASAP7_75t_L g11958 ( 
.A1(n_11539),
.A2(n_1467),
.B(n_1468),
.Y(n_11958)
);

AND2x4_ASAP7_75t_SL g11959 ( 
.A(n_11750),
.B(n_1467),
.Y(n_11959)
);

AOI22xp5_ASAP7_75t_L g11960 ( 
.A1(n_11779),
.A2(n_1470),
.B1(n_1468),
.B2(n_1469),
.Y(n_11960)
);

OAI21x1_ASAP7_75t_L g11961 ( 
.A1(n_11590),
.A2(n_1470),
.B(n_1471),
.Y(n_11961)
);

AND2x2_ASAP7_75t_L g11962 ( 
.A(n_11743),
.B(n_11751),
.Y(n_11962)
);

AOI22xp33_ASAP7_75t_L g11963 ( 
.A1(n_11566),
.A2(n_1473),
.B1(n_1471),
.B2(n_1472),
.Y(n_11963)
);

OR2x6_ASAP7_75t_L g11964 ( 
.A(n_11640),
.B(n_1473),
.Y(n_11964)
);

AOI22xp33_ASAP7_75t_L g11965 ( 
.A1(n_11559),
.A2(n_1476),
.B1(n_1474),
.B2(n_1475),
.Y(n_11965)
);

OR2x6_ASAP7_75t_L g11966 ( 
.A(n_11640),
.B(n_1474),
.Y(n_11966)
);

AND2x4_ASAP7_75t_L g11967 ( 
.A(n_11708),
.B(n_1475),
.Y(n_11967)
);

NAND2xp33_ASAP7_75t_R g11968 ( 
.A(n_11529),
.B(n_1476),
.Y(n_11968)
);

AND2x4_ASAP7_75t_L g11969 ( 
.A(n_11757),
.B(n_11652),
.Y(n_11969)
);

AOI22xp33_ASAP7_75t_L g11970 ( 
.A1(n_11561),
.A2(n_1479),
.B1(n_1477),
.B2(n_1478),
.Y(n_11970)
);

AOI22xp33_ASAP7_75t_SL g11971 ( 
.A1(n_11517),
.A2(n_1479),
.B1(n_1477),
.B2(n_1478),
.Y(n_11971)
);

INVx1_ASAP7_75t_L g11972 ( 
.A(n_11642),
.Y(n_11972)
);

INVx6_ASAP7_75t_L g11973 ( 
.A(n_11525),
.Y(n_11973)
);

INVx1_ASAP7_75t_L g11974 ( 
.A(n_11648),
.Y(n_11974)
);

BUFx4f_ASAP7_75t_SL g11975 ( 
.A(n_11563),
.Y(n_11975)
);

BUFx8_ASAP7_75t_L g11976 ( 
.A(n_11554),
.Y(n_11976)
);

INVx1_ASAP7_75t_L g11977 ( 
.A(n_11694),
.Y(n_11977)
);

OR2x2_ASAP7_75t_L g11978 ( 
.A(n_11698),
.B(n_1480),
.Y(n_11978)
);

BUFx3_ASAP7_75t_L g11979 ( 
.A(n_11643),
.Y(n_11979)
);

OAI22xp5_ASAP7_75t_L g11980 ( 
.A1(n_11597),
.A2(n_1482),
.B1(n_1480),
.B2(n_1481),
.Y(n_11980)
);

AOI22xp33_ASAP7_75t_L g11981 ( 
.A1(n_11669),
.A2(n_1483),
.B1(n_1481),
.B2(n_1482),
.Y(n_11981)
);

INVx1_ASAP7_75t_L g11982 ( 
.A(n_11702),
.Y(n_11982)
);

OAI22xp33_ASAP7_75t_L g11983 ( 
.A1(n_11635),
.A2(n_1485),
.B1(n_1483),
.B2(n_1484),
.Y(n_11983)
);

A2O1A1Ixp33_ASAP7_75t_L g11984 ( 
.A1(n_11793),
.A2(n_1486),
.B(n_1484),
.C(n_1485),
.Y(n_11984)
);

BUFx2_ASAP7_75t_SL g11985 ( 
.A(n_11774),
.Y(n_11985)
);

OAI22xp5_ASAP7_75t_L g11986 ( 
.A1(n_11575),
.A2(n_1488),
.B1(n_1486),
.B2(n_1487),
.Y(n_11986)
);

AOI21xp5_ASAP7_75t_L g11987 ( 
.A1(n_11611),
.A2(n_1487),
.B(n_1488),
.Y(n_11987)
);

INVx1_ASAP7_75t_L g11988 ( 
.A(n_11709),
.Y(n_11988)
);

CKINVDCx5p33_ASAP7_75t_R g11989 ( 
.A(n_11532),
.Y(n_11989)
);

AOI221xp5_ASAP7_75t_L g11990 ( 
.A1(n_11786),
.A2(n_1491),
.B1(n_1489),
.B2(n_1490),
.C(n_1492),
.Y(n_11990)
);

INVx3_ASAP7_75t_L g11991 ( 
.A(n_11569),
.Y(n_11991)
);

AOI22xp33_ASAP7_75t_L g11992 ( 
.A1(n_11805),
.A2(n_1492),
.B1(n_1489),
.B2(n_1491),
.Y(n_11992)
);

OAI22xp5_ASAP7_75t_L g11993 ( 
.A1(n_11592),
.A2(n_1495),
.B1(n_1493),
.B2(n_1494),
.Y(n_11993)
);

AOI22xp5_ASAP7_75t_L g11994 ( 
.A1(n_11790),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_11994)
);

INVx1_ASAP7_75t_L g11995 ( 
.A(n_11711),
.Y(n_11995)
);

AND2x2_ASAP7_75t_L g11996 ( 
.A(n_11759),
.B(n_11637),
.Y(n_11996)
);

AOI22xp33_ASAP7_75t_L g11997 ( 
.A1(n_11809),
.A2(n_1498),
.B1(n_1496),
.B2(n_1497),
.Y(n_11997)
);

OAI22xp5_ASAP7_75t_L g11998 ( 
.A1(n_11584),
.A2(n_1501),
.B1(n_1497),
.B2(n_1499),
.Y(n_11998)
);

AOI322xp5_ASAP7_75t_L g11999 ( 
.A1(n_11691),
.A2(n_1505),
.A3(n_1504),
.B1(n_1502),
.B2(n_1499),
.C1(n_1501),
.C2(n_1503),
.Y(n_11999)
);

AND2x2_ASAP7_75t_L g12000 ( 
.A(n_11543),
.B(n_1502),
.Y(n_12000)
);

INVx1_ASAP7_75t_L g12001 ( 
.A(n_11715),
.Y(n_12001)
);

INVx2_ASAP7_75t_L g12002 ( 
.A(n_11713),
.Y(n_12002)
);

AOI22xp33_ASAP7_75t_SL g12003 ( 
.A1(n_11838),
.A2(n_1505),
.B1(n_1503),
.B2(n_1504),
.Y(n_12003)
);

OAI22xp5_ASAP7_75t_L g12004 ( 
.A1(n_11582),
.A2(n_1508),
.B1(n_1506),
.B2(n_1507),
.Y(n_12004)
);

AOI22xp33_ASAP7_75t_L g12005 ( 
.A1(n_11773),
.A2(n_1510),
.B1(n_1507),
.B2(n_1509),
.Y(n_12005)
);

INVx3_ASAP7_75t_L g12006 ( 
.A(n_11778),
.Y(n_12006)
);

NAND2xp33_ASAP7_75t_R g12007 ( 
.A(n_11795),
.B(n_1509),
.Y(n_12007)
);

AOI22xp33_ASAP7_75t_L g12008 ( 
.A1(n_11666),
.A2(n_1513),
.B1(n_1511),
.B2(n_1512),
.Y(n_12008)
);

NAND2xp5_ASAP7_75t_L g12009 ( 
.A(n_11798),
.B(n_1511),
.Y(n_12009)
);

AND2x2_ASAP7_75t_L g12010 ( 
.A(n_11562),
.B(n_11799),
.Y(n_12010)
);

HB1xp67_ASAP7_75t_L g12011 ( 
.A(n_11734),
.Y(n_12011)
);

CKINVDCx5p33_ASAP7_75t_R g12012 ( 
.A(n_11594),
.Y(n_12012)
);

INVx2_ASAP7_75t_L g12013 ( 
.A(n_11651),
.Y(n_12013)
);

INVx1_ASAP7_75t_L g12014 ( 
.A(n_11716),
.Y(n_12014)
);

NAND3xp33_ASAP7_75t_SL g12015 ( 
.A(n_11815),
.B(n_1512),
.C(n_1513),
.Y(n_12015)
);

OAI22xp5_ASAP7_75t_L g12016 ( 
.A1(n_11661),
.A2(n_1516),
.B1(n_1514),
.B2(n_1515),
.Y(n_12016)
);

AOI22xp33_ASAP7_75t_L g12017 ( 
.A1(n_11675),
.A2(n_1517),
.B1(n_1514),
.B2(n_1516),
.Y(n_12017)
);

CKINVDCx20_ASAP7_75t_R g12018 ( 
.A(n_11828),
.Y(n_12018)
);

BUFx3_ASAP7_75t_L g12019 ( 
.A(n_11731),
.Y(n_12019)
);

NAND2xp5_ASAP7_75t_L g12020 ( 
.A(n_11811),
.B(n_1518),
.Y(n_12020)
);

NAND2xp5_ASAP7_75t_L g12021 ( 
.A(n_11585),
.B(n_1518),
.Y(n_12021)
);

BUFx6f_ASAP7_75t_L g12022 ( 
.A(n_11593),
.Y(n_12022)
);

INVx2_ASAP7_75t_L g12023 ( 
.A(n_11681),
.Y(n_12023)
);

INVx2_ASAP7_75t_L g12024 ( 
.A(n_11596),
.Y(n_12024)
);

OA21x2_ASAP7_75t_L g12025 ( 
.A1(n_11700),
.A2(n_1519),
.B(n_1520),
.Y(n_12025)
);

NOR2xp33_ASAP7_75t_R g12026 ( 
.A(n_11789),
.B(n_1519),
.Y(n_12026)
);

INVx2_ASAP7_75t_L g12027 ( 
.A(n_11598),
.Y(n_12027)
);

AOI22xp5_ASAP7_75t_L g12028 ( 
.A1(n_11680),
.A2(n_11813),
.B1(n_11733),
.B2(n_11654),
.Y(n_12028)
);

AOI22xp33_ASAP7_75t_L g12029 ( 
.A1(n_11744),
.A2(n_1523),
.B1(n_1520),
.B2(n_1521),
.Y(n_12029)
);

NAND2xp5_ASAP7_75t_L g12030 ( 
.A(n_11720),
.B(n_1521),
.Y(n_12030)
);

OAI22xp5_ASAP7_75t_L g12031 ( 
.A1(n_11676),
.A2(n_1525),
.B1(n_1523),
.B2(n_1524),
.Y(n_12031)
);

BUFx3_ASAP7_75t_L g12032 ( 
.A(n_11536),
.Y(n_12032)
);

NOR2xp33_ASAP7_75t_L g12033 ( 
.A(n_11513),
.B(n_1524),
.Y(n_12033)
);

AND2x2_ASAP7_75t_L g12034 ( 
.A(n_11804),
.B(n_11785),
.Y(n_12034)
);

CKINVDCx5p33_ASAP7_75t_R g12035 ( 
.A(n_11707),
.Y(n_12035)
);

O2A1O1Ixp33_ASAP7_75t_L g12036 ( 
.A1(n_11722),
.A2(n_1527),
.B(n_1525),
.C(n_1526),
.Y(n_12036)
);

INVx1_ASAP7_75t_L g12037 ( 
.A(n_11639),
.Y(n_12037)
);

AOI21xp5_ASAP7_75t_L g12038 ( 
.A1(n_11551),
.A2(n_1526),
.B(n_1527),
.Y(n_12038)
);

AO21x2_ASAP7_75t_L g12039 ( 
.A1(n_11636),
.A2(n_1528),
.B(n_1530),
.Y(n_12039)
);

OAI22xp5_ASAP7_75t_L g12040 ( 
.A1(n_11572),
.A2(n_1532),
.B1(n_1530),
.B2(n_1531),
.Y(n_12040)
);

INVx2_ASAP7_75t_L g12041 ( 
.A(n_11599),
.Y(n_12041)
);

AND2x2_ASAP7_75t_L g12042 ( 
.A(n_11717),
.B(n_1533),
.Y(n_12042)
);

AOI22xp33_ASAP7_75t_L g12043 ( 
.A1(n_11621),
.A2(n_1535),
.B1(n_1533),
.B2(n_1534),
.Y(n_12043)
);

AOI22xp5_ASAP7_75t_L g12044 ( 
.A1(n_11725),
.A2(n_1536),
.B1(n_1534),
.B2(n_1535),
.Y(n_12044)
);

AND2x2_ASAP7_75t_L g12045 ( 
.A(n_11808),
.B(n_1536),
.Y(n_12045)
);

BUFx10_ASAP7_75t_L g12046 ( 
.A(n_11578),
.Y(n_12046)
);

AOI222xp33_ASAP7_75t_L g12047 ( 
.A1(n_11817),
.A2(n_1540),
.B1(n_1542),
.B2(n_1538),
.C1(n_1539),
.C2(n_1541),
.Y(n_12047)
);

AND2x2_ASAP7_75t_L g12048 ( 
.A(n_11788),
.B(n_1540),
.Y(n_12048)
);

OAI22xp5_ASAP7_75t_L g12049 ( 
.A1(n_11613),
.A2(n_1544),
.B1(n_1541),
.B2(n_1543),
.Y(n_12049)
);

AOI22xp5_ASAP7_75t_L g12050 ( 
.A1(n_11583),
.A2(n_1546),
.B1(n_1544),
.B2(n_1545),
.Y(n_12050)
);

OAI22xp33_ASAP7_75t_L g12051 ( 
.A1(n_11665),
.A2(n_1547),
.B1(n_1545),
.B2(n_1546),
.Y(n_12051)
);

AND2x2_ASAP7_75t_L g12052 ( 
.A(n_11791),
.B(n_1547),
.Y(n_12052)
);

OAI21x1_ASAP7_75t_L g12053 ( 
.A1(n_11714),
.A2(n_1548),
.B(n_1549),
.Y(n_12053)
);

AOI22xp5_ASAP7_75t_L g12054 ( 
.A1(n_11633),
.A2(n_1550),
.B1(n_1548),
.B2(n_1549),
.Y(n_12054)
);

OA21x2_ASAP7_75t_L g12055 ( 
.A1(n_11577),
.A2(n_1550),
.B(n_1551),
.Y(n_12055)
);

OAI21x1_ASAP7_75t_L g12056 ( 
.A1(n_11600),
.A2(n_11606),
.B(n_11588),
.Y(n_12056)
);

AND2x4_ASAP7_75t_L g12057 ( 
.A(n_11658),
.B(n_1551),
.Y(n_12057)
);

BUFx2_ASAP7_75t_L g12058 ( 
.A(n_11719),
.Y(n_12058)
);

CKINVDCx6p67_ASAP7_75t_R g12059 ( 
.A(n_11792),
.Y(n_12059)
);

NOR2xp33_ASAP7_75t_L g12060 ( 
.A(n_11632),
.B(n_11557),
.Y(n_12060)
);

NAND2x1_ASAP7_75t_L g12061 ( 
.A(n_11843),
.B(n_1552),
.Y(n_12061)
);

AO31x2_ASAP7_75t_L g12062 ( 
.A1(n_11602),
.A2(n_1554),
.A3(n_1552),
.B(n_1553),
.Y(n_12062)
);

OAI22xp5_ASAP7_75t_L g12063 ( 
.A1(n_11818),
.A2(n_1556),
.B1(n_1554),
.B2(n_1555),
.Y(n_12063)
);

NAND2x1_ASAP7_75t_L g12064 ( 
.A(n_11610),
.B(n_1556),
.Y(n_12064)
);

NAND2xp5_ASAP7_75t_L g12065 ( 
.A(n_11832),
.B(n_1557),
.Y(n_12065)
);

OAI22xp5_ASAP7_75t_L g12066 ( 
.A1(n_11823),
.A2(n_1559),
.B1(n_1557),
.B2(n_1558),
.Y(n_12066)
);

INVx2_ASAP7_75t_L g12067 ( 
.A(n_11836),
.Y(n_12067)
);

AO31x2_ASAP7_75t_L g12068 ( 
.A1(n_11612),
.A2(n_1560),
.A3(n_1558),
.B(n_1559),
.Y(n_12068)
);

INVx2_ASAP7_75t_SL g12069 ( 
.A(n_11657),
.Y(n_12069)
);

OAI222xp33_ASAP7_75t_L g12070 ( 
.A1(n_11695),
.A2(n_1562),
.B1(n_1564),
.B2(n_1560),
.C1(n_1561),
.C2(n_1563),
.Y(n_12070)
);

INVx1_ASAP7_75t_L g12071 ( 
.A(n_11586),
.Y(n_12071)
);

NAND2xp5_ASAP7_75t_L g12072 ( 
.A(n_11682),
.B(n_1561),
.Y(n_12072)
);

AND2x4_ASAP7_75t_L g12073 ( 
.A(n_11662),
.B(n_1562),
.Y(n_12073)
);

INVx1_ASAP7_75t_L g12074 ( 
.A(n_11589),
.Y(n_12074)
);

AND2x4_ASAP7_75t_L g12075 ( 
.A(n_11825),
.B(n_1563),
.Y(n_12075)
);

CKINVDCx16_ASAP7_75t_R g12076 ( 
.A(n_11760),
.Y(n_12076)
);

HB1xp67_ASAP7_75t_L g12077 ( 
.A(n_11591),
.Y(n_12077)
);

NOR3xp33_ASAP7_75t_SL g12078 ( 
.A(n_11783),
.B(n_1564),
.C(n_1565),
.Y(n_12078)
);

INVx1_ASAP7_75t_L g12079 ( 
.A(n_11770),
.Y(n_12079)
);

INVx2_ASAP7_75t_L g12080 ( 
.A(n_11762),
.Y(n_12080)
);

BUFx3_ASAP7_75t_L g12081 ( 
.A(n_11776),
.Y(n_12081)
);

OR2x6_ASAP7_75t_L g12082 ( 
.A(n_11778),
.B(n_1565),
.Y(n_12082)
);

BUFx3_ASAP7_75t_L g12083 ( 
.A(n_11655),
.Y(n_12083)
);

INVx6_ASAP7_75t_L g12084 ( 
.A(n_11656),
.Y(n_12084)
);

NAND2xp5_ASAP7_75t_L g12085 ( 
.A(n_11638),
.B(n_1566),
.Y(n_12085)
);

OAI22xp33_ASAP7_75t_L g12086 ( 
.A1(n_11678),
.A2(n_1568),
.B1(n_1566),
.B2(n_1567),
.Y(n_12086)
);

NAND2xp33_ASAP7_75t_SL g12087 ( 
.A(n_11748),
.B(n_11807),
.Y(n_12087)
);

AOI22xp33_ASAP7_75t_L g12088 ( 
.A1(n_11841),
.A2(n_1570),
.B1(n_1567),
.B2(n_1569),
.Y(n_12088)
);

A2O1A1Ixp33_ASAP7_75t_L g12089 ( 
.A1(n_11728),
.A2(n_1572),
.B(n_1570),
.C(n_1571),
.Y(n_12089)
);

AND2x4_ASAP7_75t_L g12090 ( 
.A(n_11622),
.B(n_1572),
.Y(n_12090)
);

AND2x6_ASAP7_75t_L g12091 ( 
.A(n_11593),
.B(n_1573),
.Y(n_12091)
);

HB1xp67_ASAP7_75t_L g12092 ( 
.A(n_11819),
.Y(n_12092)
);

INVx2_ASAP7_75t_SL g12093 ( 
.A(n_11663),
.Y(n_12093)
);

INVx1_ASAP7_75t_L g12094 ( 
.A(n_11701),
.Y(n_12094)
);

INVxp67_ASAP7_75t_L g12095 ( 
.A(n_11650),
.Y(n_12095)
);

BUFx6f_ASAP7_75t_L g12096 ( 
.A(n_11673),
.Y(n_12096)
);

INVx1_ASAP7_75t_L g12097 ( 
.A(n_11692),
.Y(n_12097)
);

INVx1_ASAP7_75t_L g12098 ( 
.A(n_11729),
.Y(n_12098)
);

OR2x6_ASAP7_75t_SL g12099 ( 
.A(n_11723),
.B(n_1573),
.Y(n_12099)
);

OR2x2_ASAP7_75t_L g12100 ( 
.A(n_11775),
.B(n_11730),
.Y(n_12100)
);

OA21x2_ASAP7_75t_L g12101 ( 
.A1(n_11787),
.A2(n_1574),
.B(n_1576),
.Y(n_12101)
);

OAI22xp33_ASAP7_75t_L g12102 ( 
.A1(n_11670),
.A2(n_1578),
.B1(n_1574),
.B2(n_1576),
.Y(n_12102)
);

AOI22xp33_ASAP7_75t_SL g12103 ( 
.A1(n_11693),
.A2(n_1581),
.B1(n_1578),
.B2(n_1579),
.Y(n_12103)
);

AOI22xp33_ASAP7_75t_L g12104 ( 
.A1(n_11840),
.A2(n_1582),
.B1(n_1579),
.B2(n_1581),
.Y(n_12104)
);

INVx2_ASAP7_75t_L g12105 ( 
.A(n_11822),
.Y(n_12105)
);

NAND2x1_ASAP7_75t_L g12106 ( 
.A(n_11631),
.B(n_11668),
.Y(n_12106)
);

AOI21xp5_ASAP7_75t_L g12107 ( 
.A1(n_11718),
.A2(n_1582),
.B(n_1583),
.Y(n_12107)
);

AOI22xp5_ASAP7_75t_L g12108 ( 
.A1(n_11801),
.A2(n_11649),
.B1(n_11629),
.B2(n_11688),
.Y(n_12108)
);

INVx3_ASAP7_75t_L g12109 ( 
.A(n_11671),
.Y(n_12109)
);

INVx3_ASAP7_75t_L g12110 ( 
.A(n_11679),
.Y(n_12110)
);

INVx2_ASAP7_75t_SL g12111 ( 
.A(n_11745),
.Y(n_12111)
);

NAND2xp5_ASAP7_75t_L g12112 ( 
.A(n_11839),
.B(n_1583),
.Y(n_12112)
);

INVx4_ASAP7_75t_L g12113 ( 
.A(n_11726),
.Y(n_12113)
);

INVx1_ASAP7_75t_L g12114 ( 
.A(n_11831),
.Y(n_12114)
);

OAI22xp33_ASAP7_75t_L g12115 ( 
.A1(n_11641),
.A2(n_11618),
.B1(n_11739),
.B2(n_11736),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_11803),
.Y(n_12116)
);

OAI22xp5_ASAP7_75t_L g12117 ( 
.A1(n_11737),
.A2(n_1586),
.B1(n_1584),
.B2(n_1585),
.Y(n_12117)
);

OAI21xp5_ASAP7_75t_L g12118 ( 
.A1(n_11806),
.A2(n_1584),
.B(n_1585),
.Y(n_12118)
);

NOR2xp33_ASAP7_75t_L g12119 ( 
.A(n_11605),
.B(n_1586),
.Y(n_12119)
);

AOI22xp33_ASAP7_75t_L g12120 ( 
.A1(n_11756),
.A2(n_1589),
.B1(n_1587),
.B2(n_1588),
.Y(n_12120)
);

AOI22xp33_ASAP7_75t_L g12121 ( 
.A1(n_11761),
.A2(n_1590),
.B1(n_1587),
.B2(n_1588),
.Y(n_12121)
);

INVx3_ASAP7_75t_L g12122 ( 
.A(n_11697),
.Y(n_12122)
);

OAI211xp5_ASAP7_75t_SL g12123 ( 
.A1(n_11821),
.A2(n_1592),
.B(n_1590),
.C(n_1591),
.Y(n_12123)
);

NAND2xp5_ASAP7_75t_L g12124 ( 
.A(n_11673),
.B(n_1591),
.Y(n_12124)
);

AOI22xp33_ASAP7_75t_SL g12125 ( 
.A1(n_11732),
.A2(n_1594),
.B1(n_1592),
.B2(n_1593),
.Y(n_12125)
);

AND2x4_ASAP7_75t_L g12126 ( 
.A(n_11699),
.B(n_1594),
.Y(n_12126)
);

AOI22xp33_ASAP7_75t_L g12127 ( 
.A1(n_11796),
.A2(n_1597),
.B1(n_1595),
.B2(n_1596),
.Y(n_12127)
);

NAND2xp5_ASAP7_75t_L g12128 ( 
.A(n_11699),
.B(n_1595),
.Y(n_12128)
);

OAI21x1_ASAP7_75t_L g12129 ( 
.A1(n_11782),
.A2(n_1596),
.B(n_1597),
.Y(n_12129)
);

CKINVDCx6p67_ASAP7_75t_R g12130 ( 
.A(n_11810),
.Y(n_12130)
);

OR2x6_ASAP7_75t_L g12131 ( 
.A(n_11705),
.B(n_1598),
.Y(n_12131)
);

AOI22xp33_ASAP7_75t_SL g12132 ( 
.A1(n_11772),
.A2(n_1600),
.B1(n_1598),
.B2(n_1599),
.Y(n_12132)
);

NAND2x1p5_ASAP7_75t_L g12133 ( 
.A(n_11705),
.B(n_1600),
.Y(n_12133)
);

CKINVDCx6p67_ASAP7_75t_R g12134 ( 
.A(n_11735),
.Y(n_12134)
);

NAND3xp33_ASAP7_75t_L g12135 ( 
.A(n_11829),
.B(n_1601),
.C(n_1602),
.Y(n_12135)
);

INVx1_ASAP7_75t_L g12136 ( 
.A(n_11758),
.Y(n_12136)
);

AOI22xp33_ASAP7_75t_L g12137 ( 
.A1(n_11835),
.A2(n_1603),
.B1(n_1601),
.B2(n_1602),
.Y(n_12137)
);

INVx3_ASAP7_75t_L g12138 ( 
.A(n_11752),
.Y(n_12138)
);

INVxp33_ASAP7_75t_SL g12139 ( 
.A(n_11753),
.Y(n_12139)
);

INVx2_ASAP7_75t_L g12140 ( 
.A(n_11763),
.Y(n_12140)
);

AOI22xp33_ASAP7_75t_L g12141 ( 
.A1(n_11824),
.A2(n_11738),
.B1(n_11749),
.B2(n_11740),
.Y(n_12141)
);

INVx2_ASAP7_75t_L g12142 ( 
.A(n_11842),
.Y(n_12142)
);

INVxp67_ASAP7_75t_SL g12143 ( 
.A(n_11816),
.Y(n_12143)
);

BUFx4f_ASAP7_75t_L g12144 ( 
.A(n_11780),
.Y(n_12144)
);

OR2x2_ASAP7_75t_L g12145 ( 
.A(n_11826),
.B(n_1603),
.Y(n_12145)
);

NAND2x1_ASAP7_75t_L g12146 ( 
.A(n_11769),
.B(n_1604),
.Y(n_12146)
);

NAND2xp33_ASAP7_75t_R g12147 ( 
.A(n_11768),
.B(n_1605),
.Y(n_12147)
);

BUFx3_ASAP7_75t_L g12148 ( 
.A(n_11628),
.Y(n_12148)
);

INVx6_ASAP7_75t_L g12149 ( 
.A(n_11510),
.Y(n_12149)
);

INVx1_ASAP7_75t_L g12150 ( 
.A(n_11674),
.Y(n_12150)
);

NAND2xp5_ASAP7_75t_L g12151 ( 
.A(n_11820),
.B(n_1605),
.Y(n_12151)
);

INVx1_ASAP7_75t_L g12152 ( 
.A(n_11674),
.Y(n_12152)
);

AOI221xp5_ASAP7_75t_L g12153 ( 
.A1(n_11568),
.A2(n_1608),
.B1(n_1606),
.B2(n_1607),
.C(n_1609),
.Y(n_12153)
);

OAI22xp5_ASAP7_75t_L g12154 ( 
.A1(n_11579),
.A2(n_1610),
.B1(n_1606),
.B2(n_1609),
.Y(n_12154)
);

NOR2x1_ASAP7_75t_SL g12155 ( 
.A(n_11814),
.B(n_1610),
.Y(n_12155)
);

BUFx2_ASAP7_75t_SL g12156 ( 
.A(n_11523),
.Y(n_12156)
);

BUFx3_ASAP7_75t_L g12157 ( 
.A(n_11510),
.Y(n_12157)
);

NAND2xp5_ASAP7_75t_L g12158 ( 
.A(n_11820),
.B(n_1611),
.Y(n_12158)
);

OAI21x1_ASAP7_75t_L g12159 ( 
.A1(n_11812),
.A2(n_1611),
.B(n_1612),
.Y(n_12159)
);

A2O1A1Ixp33_ASAP7_75t_L g12160 ( 
.A1(n_11568),
.A2(n_1614),
.B(n_1612),
.C(n_1613),
.Y(n_12160)
);

INVx2_ASAP7_75t_SL g12161 ( 
.A(n_11514),
.Y(n_12161)
);

AOI22xp33_ASAP7_75t_L g12162 ( 
.A1(n_11833),
.A2(n_1616),
.B1(n_1614),
.B2(n_1615),
.Y(n_12162)
);

INVx6_ASAP7_75t_L g12163 ( 
.A(n_11510),
.Y(n_12163)
);

OAI22xp33_ASAP7_75t_L g12164 ( 
.A1(n_11595),
.A2(n_1617),
.B1(n_1615),
.B2(n_1616),
.Y(n_12164)
);

NAND2xp5_ASAP7_75t_L g12165 ( 
.A(n_11820),
.B(n_1619),
.Y(n_12165)
);

NAND2x1p5_ASAP7_75t_L g12166 ( 
.A(n_11634),
.B(n_1619),
.Y(n_12166)
);

INVx6_ASAP7_75t_L g12167 ( 
.A(n_11510),
.Y(n_12167)
);

AOI22xp33_ASAP7_75t_L g12168 ( 
.A1(n_11833),
.A2(n_1622),
.B1(n_1620),
.B2(n_1621),
.Y(n_12168)
);

AO21x2_ASAP7_75t_L g12169 ( 
.A1(n_11540),
.A2(n_1620),
.B(n_1621),
.Y(n_12169)
);

INVx1_ASAP7_75t_L g12170 ( 
.A(n_11674),
.Y(n_12170)
);

AOI222xp33_ASAP7_75t_L g12171 ( 
.A1(n_11568),
.A2(n_1625),
.B1(n_1627),
.B2(n_1623),
.C1(n_1624),
.C2(n_1626),
.Y(n_12171)
);

NAND2xp5_ASAP7_75t_SL g12172 ( 
.A(n_11540),
.B(n_1623),
.Y(n_12172)
);

INVx2_ASAP7_75t_L g12173 ( 
.A(n_11616),
.Y(n_12173)
);

OR2x6_ASAP7_75t_L g12174 ( 
.A(n_11520),
.B(n_1624),
.Y(n_12174)
);

CKINVDCx11_ASAP7_75t_R g12175 ( 
.A(n_11541),
.Y(n_12175)
);

AND2x2_ASAP7_75t_L g12176 ( 
.A(n_11565),
.B(n_1625),
.Y(n_12176)
);

OAI21xp33_ASAP7_75t_L g12177 ( 
.A1(n_11849),
.A2(n_1626),
.B(n_1627),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_11856),
.Y(n_12178)
);

BUFx8_ASAP7_75t_SL g12179 ( 
.A(n_11893),
.Y(n_12179)
);

OAI22xp33_ASAP7_75t_L g12180 ( 
.A1(n_11926),
.A2(n_1630),
.B1(n_1628),
.B2(n_1629),
.Y(n_12180)
);

INVx3_ASAP7_75t_L g12181 ( 
.A(n_11942),
.Y(n_12181)
);

BUFx12f_ASAP7_75t_L g12182 ( 
.A(n_12175),
.Y(n_12182)
);

AOI22xp33_ASAP7_75t_L g12183 ( 
.A1(n_12148),
.A2(n_1631),
.B1(n_1629),
.B2(n_1630),
.Y(n_12183)
);

OAI21xp5_ASAP7_75t_SL g12184 ( 
.A1(n_11915),
.A2(n_1631),
.B(n_1632),
.Y(n_12184)
);

AOI22xp5_ASAP7_75t_L g12185 ( 
.A1(n_12154),
.A2(n_1634),
.B1(n_1632),
.B2(n_1633),
.Y(n_12185)
);

NOR2xp33_ASAP7_75t_L g12186 ( 
.A(n_12149),
.B(n_1635),
.Y(n_12186)
);

NAND2xp5_ASAP7_75t_L g12187 ( 
.A(n_11987),
.B(n_1635),
.Y(n_12187)
);

AOI22xp33_ASAP7_75t_L g12188 ( 
.A1(n_11880),
.A2(n_12144),
.B1(n_12139),
.B2(n_11870),
.Y(n_12188)
);

INVx3_ASAP7_75t_L g12189 ( 
.A(n_11861),
.Y(n_12189)
);

AOI22xp5_ASAP7_75t_L g12190 ( 
.A1(n_12172),
.A2(n_1638),
.B1(n_1636),
.B2(n_1637),
.Y(n_12190)
);

AOI22xp33_ASAP7_75t_L g12191 ( 
.A1(n_11906),
.A2(n_1638),
.B1(n_1636),
.B2(n_1637),
.Y(n_12191)
);

BUFx12f_ASAP7_75t_L g12192 ( 
.A(n_12149),
.Y(n_12192)
);

AOI22xp33_ASAP7_75t_SL g12193 ( 
.A1(n_12155),
.A2(n_1641),
.B1(n_1639),
.B2(n_1640),
.Y(n_12193)
);

INVx2_ASAP7_75t_L g12194 ( 
.A(n_11846),
.Y(n_12194)
);

AOI22xp33_ASAP7_75t_SL g12195 ( 
.A1(n_12143),
.A2(n_1641),
.B1(n_1639),
.B2(n_1640),
.Y(n_12195)
);

AOI22xp33_ASAP7_75t_L g12196 ( 
.A1(n_12138),
.A2(n_1644),
.B1(n_1642),
.B2(n_1643),
.Y(n_12196)
);

INVx1_ASAP7_75t_L g12197 ( 
.A(n_11864),
.Y(n_12197)
);

AOI22xp33_ASAP7_75t_L g12198 ( 
.A1(n_11939),
.A2(n_1646),
.B1(n_1642),
.B2(n_1645),
.Y(n_12198)
);

INVx1_ASAP7_75t_L g12199 ( 
.A(n_11868),
.Y(n_12199)
);

INVx1_ASAP7_75t_L g12200 ( 
.A(n_12150),
.Y(n_12200)
);

OAI21xp33_ASAP7_75t_L g12201 ( 
.A1(n_12162),
.A2(n_1645),
.B(n_1646),
.Y(n_12201)
);

OAI22xp5_ASAP7_75t_SL g12202 ( 
.A1(n_11858),
.A2(n_1649),
.B1(n_1647),
.B2(n_1648),
.Y(n_12202)
);

AOI22xp33_ASAP7_75t_L g12203 ( 
.A1(n_11876),
.A2(n_1649),
.B1(n_1647),
.B2(n_1648),
.Y(n_12203)
);

BUFx12f_ASAP7_75t_L g12204 ( 
.A(n_12163),
.Y(n_12204)
);

OAI22xp5_ASAP7_75t_L g12205 ( 
.A1(n_11847),
.A2(n_12168),
.B1(n_11971),
.B2(n_12076),
.Y(n_12205)
);

INVx1_ASAP7_75t_L g12206 ( 
.A(n_12152),
.Y(n_12206)
);

AOI22xp33_ASAP7_75t_L g12207 ( 
.A1(n_11894),
.A2(n_1652),
.B1(n_1650),
.B2(n_1651),
.Y(n_12207)
);

INVx2_ASAP7_75t_L g12208 ( 
.A(n_12161),
.Y(n_12208)
);

AND2x2_ASAP7_75t_L g12209 ( 
.A(n_11851),
.B(n_11895),
.Y(n_12209)
);

AOI22xp33_ASAP7_75t_L g12210 ( 
.A1(n_11867),
.A2(n_1652),
.B1(n_1650),
.B2(n_1651),
.Y(n_12210)
);

OAI21xp5_ASAP7_75t_SL g12211 ( 
.A1(n_11877),
.A2(n_1653),
.B(n_1654),
.Y(n_12211)
);

BUFx2_ASAP7_75t_L g12212 ( 
.A(n_11933),
.Y(n_12212)
);

AOI22xp33_ASAP7_75t_SL g12213 ( 
.A1(n_11985),
.A2(n_1655),
.B1(n_1653),
.B2(n_1654),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_12170),
.Y(n_12214)
);

AOI22xp33_ASAP7_75t_L g12215 ( 
.A1(n_11980),
.A2(n_12040),
.B1(n_11871),
.B2(n_11913),
.Y(n_12215)
);

OAI21xp5_ASAP7_75t_SL g12216 ( 
.A1(n_11872),
.A2(n_1656),
.B(n_1657),
.Y(n_12216)
);

AOI22xp33_ASAP7_75t_L g12217 ( 
.A1(n_11916),
.A2(n_12169),
.B1(n_12015),
.B2(n_12038),
.Y(n_12217)
);

AOI22xp33_ASAP7_75t_L g12218 ( 
.A1(n_12142),
.A2(n_1658),
.B1(n_1656),
.B2(n_1657),
.Y(n_12218)
);

AOI22xp5_ASAP7_75t_L g12219 ( 
.A1(n_12007),
.A2(n_1660),
.B1(n_1658),
.B2(n_1659),
.Y(n_12219)
);

INVx1_ASAP7_75t_L g12220 ( 
.A(n_11879),
.Y(n_12220)
);

INVx2_ASAP7_75t_L g12221 ( 
.A(n_11905),
.Y(n_12221)
);

AND2x2_ASAP7_75t_L g12222 ( 
.A(n_11962),
.B(n_1659),
.Y(n_12222)
);

OAI21xp5_ASAP7_75t_SL g12223 ( 
.A1(n_12028),
.A2(n_1661),
.B(n_1663),
.Y(n_12223)
);

AOI22xp33_ASAP7_75t_L g12224 ( 
.A1(n_12140),
.A2(n_1665),
.B1(n_1661),
.B2(n_1664),
.Y(n_12224)
);

OAI22xp33_ASAP7_75t_SL g12225 ( 
.A1(n_12084),
.A2(n_1669),
.B1(n_1666),
.B2(n_1668),
.Y(n_12225)
);

INVx1_ASAP7_75t_L g12226 ( 
.A(n_11884),
.Y(n_12226)
);

BUFx4f_ASAP7_75t_SL g12227 ( 
.A(n_12018),
.Y(n_12227)
);

AOI22xp33_ASAP7_75t_L g12228 ( 
.A1(n_11970),
.A2(n_1672),
.B1(n_1670),
.B2(n_1671),
.Y(n_12228)
);

AOI22xp33_ASAP7_75t_L g12229 ( 
.A1(n_11892),
.A2(n_1672),
.B1(n_1670),
.B2(n_1671),
.Y(n_12229)
);

BUFx2_ASAP7_75t_L g12230 ( 
.A(n_11850),
.Y(n_12230)
);

AOI22xp33_ASAP7_75t_SL g12231 ( 
.A1(n_11859),
.A2(n_1675),
.B1(n_1673),
.B2(n_1674),
.Y(n_12231)
);

BUFx3_ASAP7_75t_L g12232 ( 
.A(n_11855),
.Y(n_12232)
);

AOI22xp33_ASAP7_75t_L g12233 ( 
.A1(n_12153),
.A2(n_1676),
.B1(n_1673),
.B2(n_1674),
.Y(n_12233)
);

INVx2_ASAP7_75t_L g12234 ( 
.A(n_11905),
.Y(n_12234)
);

INVx2_ASAP7_75t_L g12235 ( 
.A(n_12084),
.Y(n_12235)
);

NAND2xp5_ASAP7_75t_SL g12236 ( 
.A(n_12115),
.B(n_1676),
.Y(n_12236)
);

AOI22xp33_ASAP7_75t_L g12237 ( 
.A1(n_11925),
.A2(n_1680),
.B1(n_1677),
.B2(n_1679),
.Y(n_12237)
);

AND2x4_ASAP7_75t_L g12238 ( 
.A(n_12069),
.B(n_1677),
.Y(n_12238)
);

AND2x2_ASAP7_75t_L g12239 ( 
.A(n_11996),
.B(n_1679),
.Y(n_12239)
);

AOI222xp33_ASAP7_75t_L g12240 ( 
.A1(n_11885),
.A2(n_1682),
.B1(n_1684),
.B2(n_1680),
.C1(n_1681),
.C2(n_1683),
.Y(n_12240)
);

OAI22xp5_ASAP7_75t_L g12241 ( 
.A1(n_12050),
.A2(n_11937),
.B1(n_12141),
.B2(n_12099),
.Y(n_12241)
);

AOI22xp33_ASAP7_75t_L g12242 ( 
.A1(n_12171),
.A2(n_1685),
.B1(n_1681),
.B2(n_1682),
.Y(n_12242)
);

INVx1_ASAP7_75t_L g12243 ( 
.A(n_11901),
.Y(n_12243)
);

AOI22xp33_ASAP7_75t_SL g12244 ( 
.A1(n_11952),
.A2(n_1687),
.B1(n_1685),
.B2(n_1686),
.Y(n_12244)
);

OAI22xp5_ASAP7_75t_L g12245 ( 
.A1(n_11920),
.A2(n_1688),
.B1(n_1686),
.B2(n_1687),
.Y(n_12245)
);

OAI22xp5_ASAP7_75t_L g12246 ( 
.A1(n_11908),
.A2(n_1690),
.B1(n_1688),
.B2(n_1689),
.Y(n_12246)
);

AOI22xp33_ASAP7_75t_L g12247 ( 
.A1(n_12135),
.A2(n_1691),
.B1(n_1689),
.B2(n_1690),
.Y(n_12247)
);

INVx5_ASAP7_75t_L g12248 ( 
.A(n_12163),
.Y(n_12248)
);

AOI22xp33_ASAP7_75t_L g12249 ( 
.A1(n_12118),
.A2(n_1693),
.B1(n_1691),
.B2(n_1692),
.Y(n_12249)
);

OAI22xp5_ASAP7_75t_L g12250 ( 
.A1(n_12164),
.A2(n_1694),
.B1(n_1692),
.B2(n_1693),
.Y(n_12250)
);

AOI22xp33_ASAP7_75t_L g12251 ( 
.A1(n_11948),
.A2(n_1696),
.B1(n_1694),
.B2(n_1695),
.Y(n_12251)
);

OAI21xp5_ASAP7_75t_SL g12252 ( 
.A1(n_12108),
.A2(n_1697),
.B(n_1698),
.Y(n_12252)
);

AOI22xp33_ASAP7_75t_L g12253 ( 
.A1(n_12123),
.A2(n_1699),
.B1(n_1697),
.B2(n_1698),
.Y(n_12253)
);

OR2x2_ASAP7_75t_L g12254 ( 
.A(n_11950),
.B(n_1699),
.Y(n_12254)
);

AOI222xp33_ASAP7_75t_L g12255 ( 
.A1(n_11903),
.A2(n_1702),
.B1(n_1704),
.B2(n_1700),
.C1(n_1701),
.C2(n_1703),
.Y(n_12255)
);

NAND2xp5_ASAP7_75t_L g12256 ( 
.A(n_12094),
.B(n_1700),
.Y(n_12256)
);

OAI21xp5_ASAP7_75t_SL g12257 ( 
.A1(n_11954),
.A2(n_1701),
.B(n_1702),
.Y(n_12257)
);

BUFx4f_ASAP7_75t_L g12258 ( 
.A(n_12167),
.Y(n_12258)
);

OAI22xp5_ASAP7_75t_SL g12259 ( 
.A1(n_11853),
.A2(n_1706),
.B1(n_1704),
.B2(n_1705),
.Y(n_12259)
);

INVx3_ASAP7_75t_L g12260 ( 
.A(n_11861),
.Y(n_12260)
);

CKINVDCx20_ASAP7_75t_R g12261 ( 
.A(n_11919),
.Y(n_12261)
);

INVx1_ASAP7_75t_L g12262 ( 
.A(n_11907),
.Y(n_12262)
);

AOI22xp33_ASAP7_75t_L g12263 ( 
.A1(n_12049),
.A2(n_1707),
.B1(n_1705),
.B2(n_1706),
.Y(n_12263)
);

OAI22xp33_ASAP7_75t_L g12264 ( 
.A1(n_11968),
.A2(n_1710),
.B1(n_1708),
.B2(n_1709),
.Y(n_12264)
);

NOR2xp33_ASAP7_75t_SL g12265 ( 
.A(n_12059),
.B(n_1708),
.Y(n_12265)
);

BUFx2_ASAP7_75t_L g12266 ( 
.A(n_12130),
.Y(n_12266)
);

BUFx4f_ASAP7_75t_SL g12267 ( 
.A(n_11893),
.Y(n_12267)
);

INVx1_ASAP7_75t_L g12268 ( 
.A(n_11910),
.Y(n_12268)
);

OAI21xp5_ASAP7_75t_L g12269 ( 
.A1(n_11869),
.A2(n_1710),
.B(n_1711),
.Y(n_12269)
);

AOI22xp33_ASAP7_75t_L g12270 ( 
.A1(n_11993),
.A2(n_1713),
.B1(n_1711),
.B2(n_1712),
.Y(n_12270)
);

AOI22xp33_ASAP7_75t_L g12271 ( 
.A1(n_12004),
.A2(n_1714),
.B1(n_1712),
.B2(n_1713),
.Y(n_12271)
);

INVx5_ASAP7_75t_SL g12272 ( 
.A(n_12174),
.Y(n_12272)
);

HB1xp67_ASAP7_75t_L g12273 ( 
.A(n_11865),
.Y(n_12273)
);

AOI22xp33_ASAP7_75t_L g12274 ( 
.A1(n_11986),
.A2(n_1717),
.B1(n_1714),
.B2(n_1716),
.Y(n_12274)
);

INVx2_ASAP7_75t_L g12275 ( 
.A(n_12058),
.Y(n_12275)
);

NAND2xp5_ASAP7_75t_L g12276 ( 
.A(n_12095),
.B(n_1716),
.Y(n_12276)
);

OAI22xp5_ASAP7_75t_L g12277 ( 
.A1(n_11853),
.A2(n_1719),
.B1(n_1717),
.B2(n_1718),
.Y(n_12277)
);

INVx1_ASAP7_75t_L g12278 ( 
.A(n_11917),
.Y(n_12278)
);

INVx2_ASAP7_75t_L g12279 ( 
.A(n_12093),
.Y(n_12279)
);

BUFx2_ASAP7_75t_L g12280 ( 
.A(n_12081),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_11923),
.Y(n_12281)
);

AOI22xp33_ASAP7_75t_SL g12282 ( 
.A1(n_12026),
.A2(n_1720),
.B1(n_1718),
.B2(n_1719),
.Y(n_12282)
);

AOI22xp33_ASAP7_75t_SL g12283 ( 
.A1(n_11998),
.A2(n_1722),
.B1(n_1720),
.B2(n_1721),
.Y(n_12283)
);

AOI22xp33_ASAP7_75t_L g12284 ( 
.A1(n_11990),
.A2(n_1724),
.B1(n_1722),
.B2(n_1723),
.Y(n_12284)
);

NAND2xp5_ASAP7_75t_L g12285 ( 
.A(n_12025),
.B(n_1723),
.Y(n_12285)
);

NAND2xp5_ASAP7_75t_L g12286 ( 
.A(n_12097),
.B(n_1725),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_11931),
.Y(n_12287)
);

HB1xp67_ASAP7_75t_L g12288 ( 
.A(n_11881),
.Y(n_12288)
);

INVx1_ASAP7_75t_L g12289 ( 
.A(n_11934),
.Y(n_12289)
);

AND2x2_ASAP7_75t_L g12290 ( 
.A(n_12105),
.B(n_1725),
.Y(n_12290)
);

BUFx3_ASAP7_75t_L g12291 ( 
.A(n_11855),
.Y(n_12291)
);

BUFx3_ASAP7_75t_L g12292 ( 
.A(n_12167),
.Y(n_12292)
);

AND2x2_ASAP7_75t_L g12293 ( 
.A(n_12010),
.B(n_1726),
.Y(n_12293)
);

CKINVDCx20_ASAP7_75t_R g12294 ( 
.A(n_11975),
.Y(n_12294)
);

OAI21xp33_ASAP7_75t_L g12295 ( 
.A1(n_12078),
.A2(n_1727),
.B(n_1728),
.Y(n_12295)
);

OAI21xp5_ASAP7_75t_L g12296 ( 
.A1(n_12160),
.A2(n_1727),
.B(n_1728),
.Y(n_12296)
);

OAI22xp5_ASAP7_75t_L g12297 ( 
.A1(n_11938),
.A2(n_1731),
.B1(n_1729),
.B2(n_1730),
.Y(n_12297)
);

AOI22xp33_ASAP7_75t_L g12298 ( 
.A1(n_11911),
.A2(n_11930),
.B1(n_12119),
.B2(n_12087),
.Y(n_12298)
);

AOI22xp33_ASAP7_75t_L g12299 ( 
.A1(n_12047),
.A2(n_12114),
.B1(n_11897),
.B2(n_11878),
.Y(n_12299)
);

OAI22xp5_ASAP7_75t_L g12300 ( 
.A1(n_12116),
.A2(n_1732),
.B1(n_1729),
.B2(n_1731),
.Y(n_12300)
);

HB1xp67_ASAP7_75t_L g12301 ( 
.A(n_12011),
.Y(n_12301)
);

NOR2xp33_ASAP7_75t_R g12302 ( 
.A(n_11973),
.B(n_1732),
.Y(n_12302)
);

NAND2xp5_ASAP7_75t_L g12303 ( 
.A(n_12098),
.B(n_1733),
.Y(n_12303)
);

AOI22xp33_ASAP7_75t_SL g12304 ( 
.A1(n_11866),
.A2(n_1735),
.B1(n_1733),
.B2(n_1734),
.Y(n_12304)
);

AOI22xp33_ASAP7_75t_L g12305 ( 
.A1(n_12063),
.A2(n_1736),
.B1(n_1734),
.B2(n_1735),
.Y(n_12305)
);

AOI22xp33_ASAP7_75t_SL g12306 ( 
.A1(n_12166),
.A2(n_1738),
.B1(n_1736),
.B2(n_1737),
.Y(n_12306)
);

OAI22xp5_ASAP7_75t_L g12307 ( 
.A1(n_11857),
.A2(n_1740),
.B1(n_1737),
.B2(n_1739),
.Y(n_12307)
);

NOR2xp33_ASAP7_75t_L g12308 ( 
.A(n_11854),
.B(n_1740),
.Y(n_12308)
);

INVx1_ASAP7_75t_L g12309 ( 
.A(n_11946),
.Y(n_12309)
);

NAND3xp33_ASAP7_75t_L g12310 ( 
.A(n_11999),
.B(n_1741),
.C(n_1742),
.Y(n_12310)
);

OAI21xp5_ASAP7_75t_SL g12311 ( 
.A1(n_12036),
.A2(n_1741),
.B(n_1743),
.Y(n_12311)
);

AOI22xp33_ASAP7_75t_L g12312 ( 
.A1(n_11955),
.A2(n_1745),
.B1(n_1743),
.B2(n_1744),
.Y(n_12312)
);

HB1xp67_ASAP7_75t_L g12313 ( 
.A(n_11951),
.Y(n_12313)
);

AND2x2_ASAP7_75t_L g12314 ( 
.A(n_12034),
.B(n_1744),
.Y(n_12314)
);

INVx6_ASAP7_75t_L g12315 ( 
.A(n_11976),
.Y(n_12315)
);

AOI22xp33_ASAP7_75t_L g12316 ( 
.A1(n_12146),
.A2(n_12156),
.B1(n_12117),
.B2(n_12016),
.Y(n_12316)
);

INVx4_ASAP7_75t_L g12317 ( 
.A(n_11973),
.Y(n_12317)
);

AOI22xp33_ASAP7_75t_L g12318 ( 
.A1(n_12031),
.A2(n_1747),
.B1(n_1745),
.B2(n_1746),
.Y(n_12318)
);

INVx2_ASAP7_75t_L g12319 ( 
.A(n_12109),
.Y(n_12319)
);

NAND2xp5_ASAP7_75t_L g12320 ( 
.A(n_12101),
.B(n_11914),
.Y(n_12320)
);

OAI22xp33_ASAP7_75t_L g12321 ( 
.A1(n_12147),
.A2(n_1748),
.B1(n_1746),
.B2(n_1747),
.Y(n_12321)
);

INVx1_ASAP7_75t_L g12322 ( 
.A(n_11956),
.Y(n_12322)
);

BUFx2_ASAP7_75t_L g12323 ( 
.A(n_11875),
.Y(n_12323)
);

OAI21xp5_ASAP7_75t_SL g12324 ( 
.A1(n_11965),
.A2(n_1748),
.B(n_1749),
.Y(n_12324)
);

AOI22xp33_ASAP7_75t_SL g12325 ( 
.A1(n_11904),
.A2(n_1751),
.B1(n_1749),
.B2(n_1750),
.Y(n_12325)
);

OAI222xp33_ASAP7_75t_L g12326 ( 
.A1(n_11860),
.A2(n_1753),
.B1(n_1755),
.B2(n_1751),
.C1(n_1752),
.C2(n_1754),
.Y(n_12326)
);

INVx1_ASAP7_75t_L g12327 ( 
.A(n_11957),
.Y(n_12327)
);

OAI22xp5_ASAP7_75t_L g12328 ( 
.A1(n_11994),
.A2(n_1754),
.B1(n_1752),
.B2(n_1753),
.Y(n_12328)
);

AOI22xp33_ASAP7_75t_SL g12329 ( 
.A1(n_12039),
.A2(n_1758),
.B1(n_1756),
.B2(n_1757),
.Y(n_12329)
);

NOR2x1_ASAP7_75t_R g12330 ( 
.A(n_11852),
.B(n_1757),
.Y(n_12330)
);

OAI21xp33_ASAP7_75t_L g12331 ( 
.A1(n_11921),
.A2(n_1758),
.B(n_1759),
.Y(n_12331)
);

INVxp67_ASAP7_75t_L g12332 ( 
.A(n_11863),
.Y(n_12332)
);

CKINVDCx11_ASAP7_75t_R g12333 ( 
.A(n_11949),
.Y(n_12333)
);

BUFx3_ASAP7_75t_L g12334 ( 
.A(n_12157),
.Y(n_12334)
);

AOI22xp33_ASAP7_75t_L g12335 ( 
.A1(n_12066),
.A2(n_1763),
.B1(n_1760),
.B2(n_1761),
.Y(n_12335)
);

INVx1_ASAP7_75t_L g12336 ( 
.A(n_11972),
.Y(n_12336)
);

OAI22xp5_ASAP7_75t_L g12337 ( 
.A1(n_12110),
.A2(n_1765),
.B1(n_1763),
.B2(n_1764),
.Y(n_12337)
);

INVx5_ASAP7_75t_SL g12338 ( 
.A(n_12174),
.Y(n_12338)
);

INVx1_ASAP7_75t_L g12339 ( 
.A(n_11977),
.Y(n_12339)
);

INVx1_ASAP7_75t_L g12340 ( 
.A(n_11982),
.Y(n_12340)
);

OR2x2_ASAP7_75t_L g12341 ( 
.A(n_11924),
.B(n_1764),
.Y(n_12341)
);

AOI22xp33_ASAP7_75t_SL g12342 ( 
.A1(n_11889),
.A2(n_1767),
.B1(n_1765),
.B2(n_1766),
.Y(n_12342)
);

CKINVDCx5p33_ASAP7_75t_R g12343 ( 
.A(n_11928),
.Y(n_12343)
);

INVx1_ASAP7_75t_L g12344 ( 
.A(n_11988),
.Y(n_12344)
);

INVx1_ASAP7_75t_L g12345 ( 
.A(n_11995),
.Y(n_12345)
);

AOI22xp33_ASAP7_75t_L g12346 ( 
.A1(n_11845),
.A2(n_1768),
.B1(n_1766),
.B2(n_1767),
.Y(n_12346)
);

AND2x2_ASAP7_75t_L g12347 ( 
.A(n_12122),
.B(n_1768),
.Y(n_12347)
);

INVx2_ASAP7_75t_L g12348 ( 
.A(n_11896),
.Y(n_12348)
);

BUFx6f_ASAP7_75t_L g12349 ( 
.A(n_12083),
.Y(n_12349)
);

INVx1_ASAP7_75t_L g12350 ( 
.A(n_12001),
.Y(n_12350)
);

INVx1_ASAP7_75t_L g12351 ( 
.A(n_12014),
.Y(n_12351)
);

INVx2_ASAP7_75t_L g12352 ( 
.A(n_11900),
.Y(n_12352)
);

INVx2_ASAP7_75t_L g12353 ( 
.A(n_12006),
.Y(n_12353)
);

AOI22xp33_ASAP7_75t_L g12354 ( 
.A1(n_11963),
.A2(n_12107),
.B1(n_12017),
.B2(n_11981),
.Y(n_12354)
);

BUFx8_ASAP7_75t_SL g12355 ( 
.A(n_11891),
.Y(n_12355)
);

AOI22xp33_ASAP7_75t_L g12356 ( 
.A1(n_12008),
.A2(n_1771),
.B1(n_1769),
.B2(n_1770),
.Y(n_12356)
);

OAI22xp33_ASAP7_75t_SL g12357 ( 
.A1(n_12061),
.A2(n_1774),
.B1(n_1769),
.B2(n_1773),
.Y(n_12357)
);

AOI22xp33_ASAP7_75t_L g12358 ( 
.A1(n_12005),
.A2(n_1775),
.B1(n_1773),
.B2(n_1774),
.Y(n_12358)
);

OAI22x1_ASAP7_75t_L g12359 ( 
.A1(n_11969),
.A2(n_1777),
.B1(n_1775),
.B2(n_1776),
.Y(n_12359)
);

BUFx3_ASAP7_75t_L g12360 ( 
.A(n_11909),
.Y(n_12360)
);

INVx1_ASAP7_75t_L g12361 ( 
.A(n_11974),
.Y(n_12361)
);

AND2x2_ASAP7_75t_L g12362 ( 
.A(n_12111),
.B(n_1776),
.Y(n_12362)
);

INVx1_ASAP7_75t_L g12363 ( 
.A(n_12077),
.Y(n_12363)
);

BUFx3_ASAP7_75t_L g12364 ( 
.A(n_12019),
.Y(n_12364)
);

NAND2xp5_ASAP7_75t_L g12365 ( 
.A(n_11886),
.B(n_1777),
.Y(n_12365)
);

BUFx3_ASAP7_75t_L g12366 ( 
.A(n_11979),
.Y(n_12366)
);

AOI22xp33_ASAP7_75t_L g12367 ( 
.A1(n_12067),
.A2(n_1780),
.B1(n_1778),
.B2(n_1779),
.Y(n_12367)
);

AOI22xp33_ASAP7_75t_L g12368 ( 
.A1(n_12145),
.A2(n_12088),
.B1(n_12003),
.B2(n_12137),
.Y(n_12368)
);

INVx1_ASAP7_75t_L g12369 ( 
.A(n_12071),
.Y(n_12369)
);

BUFx3_ASAP7_75t_L g12370 ( 
.A(n_12134),
.Y(n_12370)
);

AOI222xp33_ASAP7_75t_L g12371 ( 
.A1(n_12070),
.A2(n_1782),
.B1(n_1784),
.B2(n_1778),
.C1(n_1781),
.C2(n_1783),
.Y(n_12371)
);

BUFx2_ASAP7_75t_L g12372 ( 
.A(n_11991),
.Y(n_12372)
);

INVx1_ASAP7_75t_L g12373 ( 
.A(n_12074),
.Y(n_12373)
);

AOI22xp33_ASAP7_75t_L g12374 ( 
.A1(n_12044),
.A2(n_1783),
.B1(n_1781),
.B2(n_1782),
.Y(n_12374)
);

CKINVDCx20_ASAP7_75t_R g12375 ( 
.A(n_12012),
.Y(n_12375)
);

INVx1_ASAP7_75t_L g12376 ( 
.A(n_12079),
.Y(n_12376)
);

INVx2_ASAP7_75t_L g12377 ( 
.A(n_12022),
.Y(n_12377)
);

BUFx12f_ASAP7_75t_L g12378 ( 
.A(n_11936),
.Y(n_12378)
);

AOI22xp5_ASAP7_75t_L g12379 ( 
.A1(n_12054),
.A2(n_1786),
.B1(n_1784),
.B2(n_1785),
.Y(n_12379)
);

AOI22xp33_ASAP7_75t_L g12380 ( 
.A1(n_11883),
.A2(n_1789),
.B1(n_1785),
.B2(n_1787),
.Y(n_12380)
);

OAI21xp5_ASAP7_75t_SL g12381 ( 
.A1(n_12125),
.A2(n_1787),
.B(n_1789),
.Y(n_12381)
);

AOI22xp33_ASAP7_75t_L g12382 ( 
.A1(n_12120),
.A2(n_1792),
.B1(n_1790),
.B2(n_1791),
.Y(n_12382)
);

BUFx3_ASAP7_75t_L g12383 ( 
.A(n_12046),
.Y(n_12383)
);

NOR2xp33_ASAP7_75t_L g12384 ( 
.A(n_12113),
.B(n_1790),
.Y(n_12384)
);

INVx1_ASAP7_75t_L g12385 ( 
.A(n_11944),
.Y(n_12385)
);

AOI22xp33_ASAP7_75t_L g12386 ( 
.A1(n_12121),
.A2(n_1793),
.B1(n_1791),
.B2(n_1792),
.Y(n_12386)
);

OAI22xp5_ASAP7_75t_L g12387 ( 
.A1(n_11960),
.A2(n_1796),
.B1(n_1793),
.B2(n_1794),
.Y(n_12387)
);

OAI21xp5_ASAP7_75t_SL g12388 ( 
.A1(n_12132),
.A2(n_1794),
.B(n_1796),
.Y(n_12388)
);

BUFx6f_ASAP7_75t_L g12389 ( 
.A(n_12075),
.Y(n_12389)
);

BUFx6f_ASAP7_75t_L g12390 ( 
.A(n_12057),
.Y(n_12390)
);

AOI22xp33_ASAP7_75t_L g12391 ( 
.A1(n_12103),
.A2(n_1799),
.B1(n_1797),
.B2(n_1798),
.Y(n_12391)
);

INVx1_ASAP7_75t_L g12392 ( 
.A(n_12080),
.Y(n_12392)
);

AOI22xp33_ASAP7_75t_SL g12393 ( 
.A1(n_11888),
.A2(n_1800),
.B1(n_1797),
.B2(n_1799),
.Y(n_12393)
);

CKINVDCx5p33_ASAP7_75t_R g12394 ( 
.A(n_11912),
.Y(n_12394)
);

INVx4_ASAP7_75t_L g12395 ( 
.A(n_12035),
.Y(n_12395)
);

OAI22xp5_ASAP7_75t_L g12396 ( 
.A1(n_12100),
.A2(n_1803),
.B1(n_1801),
.B2(n_1802),
.Y(n_12396)
);

AOI22xp33_ASAP7_75t_L g12397 ( 
.A1(n_11992),
.A2(n_1805),
.B1(n_1801),
.B2(n_1804),
.Y(n_12397)
);

AOI22xp33_ASAP7_75t_L g12398 ( 
.A1(n_11997),
.A2(n_1806),
.B1(n_1804),
.B2(n_1805),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_12127),
.A2(n_1808),
.B1(n_1806),
.B2(n_1807),
.Y(n_12399)
);

OAI22xp5_ASAP7_75t_L g12400 ( 
.A1(n_11984),
.A2(n_1810),
.B1(n_1807),
.B2(n_1809),
.Y(n_12400)
);

INVx6_ASAP7_75t_L g12401 ( 
.A(n_11964),
.Y(n_12401)
);

AOI22xp33_ASAP7_75t_SL g12402 ( 
.A1(n_12055),
.A2(n_1811),
.B1(n_1809),
.B2(n_1810),
.Y(n_12402)
);

INVx1_ASAP7_75t_L g12403 ( 
.A(n_12037),
.Y(n_12403)
);

OAI22xp5_ASAP7_75t_L g12404 ( 
.A1(n_12106),
.A2(n_1813),
.B1(n_1811),
.B2(n_1812),
.Y(n_12404)
);

AOI22xp33_ASAP7_75t_L g12405 ( 
.A1(n_11953),
.A2(n_1815),
.B1(n_1812),
.B2(n_1814),
.Y(n_12405)
);

AOI22xp33_ASAP7_75t_L g12406 ( 
.A1(n_12002),
.A2(n_1817),
.B1(n_1815),
.B2(n_1816),
.Y(n_12406)
);

AOI22xp33_ASAP7_75t_L g12407 ( 
.A1(n_11873),
.A2(n_1820),
.B1(n_1818),
.B2(n_1819),
.Y(n_12407)
);

OAI22xp33_ASAP7_75t_L g12408 ( 
.A1(n_12151),
.A2(n_1820),
.B1(n_1818),
.B2(n_1819),
.Y(n_12408)
);

NAND2xp5_ASAP7_75t_L g12409 ( 
.A(n_11887),
.B(n_1821),
.Y(n_12409)
);

NAND2xp5_ASAP7_75t_L g12410 ( 
.A(n_11929),
.B(n_1821),
.Y(n_12410)
);

AOI22xp33_ASAP7_75t_L g12411 ( 
.A1(n_12032),
.A2(n_1824),
.B1(n_1822),
.B2(n_1823),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_12024),
.Y(n_12412)
);

AND2x2_ASAP7_75t_L g12413 ( 
.A(n_12176),
.B(n_1822),
.Y(n_12413)
);

AOI22xp33_ASAP7_75t_L g12414 ( 
.A1(n_11941),
.A2(n_1825),
.B1(n_1823),
.B2(n_1824),
.Y(n_12414)
);

OAI22xp5_ASAP7_75t_L g12415 ( 
.A1(n_12158),
.A2(n_1827),
.B1(n_1825),
.B2(n_1826),
.Y(n_12415)
);

AOI222xp33_ASAP7_75t_L g12416 ( 
.A1(n_12029),
.A2(n_1829),
.B1(n_1831),
.B2(n_1827),
.C1(n_1828),
.C2(n_1830),
.Y(n_12416)
);

INVx3_ASAP7_75t_L g12417 ( 
.A(n_12022),
.Y(n_12417)
);

NAND2xp5_ASAP7_75t_L g12418 ( 
.A(n_12165),
.B(n_1828),
.Y(n_12418)
);

AND2x2_ASAP7_75t_L g12419 ( 
.A(n_12092),
.B(n_1829),
.Y(n_12419)
);

HB1xp67_ASAP7_75t_L g12420 ( 
.A(n_12027),
.Y(n_12420)
);

OAI21xp5_ASAP7_75t_L g12421 ( 
.A1(n_11958),
.A2(n_1832),
.B(n_1833),
.Y(n_12421)
);

INVx1_ASAP7_75t_L g12422 ( 
.A(n_12041),
.Y(n_12422)
);

OAI22xp33_ASAP7_75t_L g12423 ( 
.A1(n_11964),
.A2(n_1835),
.B1(n_1832),
.B2(n_1834),
.Y(n_12423)
);

NAND2xp5_ASAP7_75t_L g12424 ( 
.A(n_11899),
.B(n_1834),
.Y(n_12424)
);

NAND2xp5_ASAP7_75t_SL g12425 ( 
.A(n_11890),
.B(n_12096),
.Y(n_12425)
);

BUFx3_ASAP7_75t_L g12426 ( 
.A(n_11959),
.Y(n_12426)
);

AOI22xp33_ASAP7_75t_SL g12427 ( 
.A1(n_12091),
.A2(n_1837),
.B1(n_1835),
.B2(n_1836),
.Y(n_12427)
);

INVx2_ASAP7_75t_L g12428 ( 
.A(n_12096),
.Y(n_12428)
);

OAI22xp5_ASAP7_75t_L g12429 ( 
.A1(n_12089),
.A2(n_1838),
.B1(n_1836),
.B2(n_1837),
.Y(n_12429)
);

CKINVDCx5p33_ASAP7_75t_R g12430 ( 
.A(n_11989),
.Y(n_12430)
);

NAND2xp5_ASAP7_75t_L g12431 ( 
.A(n_11918),
.B(n_1838),
.Y(n_12431)
);

INVx1_ASAP7_75t_L g12432 ( 
.A(n_12013),
.Y(n_12432)
);

INVx1_ASAP7_75t_L g12433 ( 
.A(n_12023),
.Y(n_12433)
);

CKINVDCx5p33_ASAP7_75t_R g12434 ( 
.A(n_11936),
.Y(n_12434)
);

BUFx4f_ASAP7_75t_SL g12435 ( 
.A(n_12091),
.Y(n_12435)
);

INVx1_ASAP7_75t_L g12436 ( 
.A(n_12030),
.Y(n_12436)
);

AOI22xp33_ASAP7_75t_L g12437 ( 
.A1(n_12043),
.A2(n_1841),
.B1(n_1839),
.B2(n_1840),
.Y(n_12437)
);

AOI22xp33_ASAP7_75t_SL g12438 ( 
.A1(n_12091),
.A2(n_1842),
.B1(n_1839),
.B2(n_1841),
.Y(n_12438)
);

NOR2xp33_ASAP7_75t_L g12439 ( 
.A(n_12060),
.B(n_1842),
.Y(n_12439)
);

HB1xp67_ASAP7_75t_L g12440 ( 
.A(n_11935),
.Y(n_12440)
);

AOI22xp33_ASAP7_75t_L g12441 ( 
.A1(n_11947),
.A2(n_1845),
.B1(n_1843),
.B2(n_1844),
.Y(n_12441)
);

AND2x2_ASAP7_75t_L g12442 ( 
.A(n_12048),
.B(n_1843),
.Y(n_12442)
);

AOI22xp33_ASAP7_75t_L g12443 ( 
.A1(n_12104),
.A2(n_1848),
.B1(n_1846),
.B2(n_1847),
.Y(n_12443)
);

AND2x2_ASAP7_75t_L g12444 ( 
.A(n_12042),
.B(n_1846),
.Y(n_12444)
);

BUFx2_ASAP7_75t_L g12445 ( 
.A(n_11966),
.Y(n_12445)
);

BUFx4f_ASAP7_75t_SL g12446 ( 
.A(n_11967),
.Y(n_12446)
);

INVx1_ASAP7_75t_L g12447 ( 
.A(n_12009),
.Y(n_12447)
);

AOI22xp33_ASAP7_75t_SL g12448 ( 
.A1(n_12133),
.A2(n_1849),
.B1(n_1847),
.B2(n_1848),
.Y(n_12448)
);

HB1xp67_ASAP7_75t_L g12449 ( 
.A(n_12056),
.Y(n_12449)
);

AOI22xp33_ASAP7_75t_L g12450 ( 
.A1(n_11945),
.A2(n_11943),
.B1(n_12033),
.B2(n_12136),
.Y(n_12450)
);

OAI21xp5_ASAP7_75t_SL g12451 ( 
.A1(n_11983),
.A2(n_1849),
.B(n_1850),
.Y(n_12451)
);

AOI22xp33_ASAP7_75t_L g12452 ( 
.A1(n_11966),
.A2(n_1853),
.B1(n_1850),
.B2(n_1851),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_12020),
.Y(n_12453)
);

INVx4_ASAP7_75t_L g12454 ( 
.A(n_12082),
.Y(n_12454)
);

NAND2xp5_ASAP7_75t_SL g12455 ( 
.A(n_11932),
.B(n_1853),
.Y(n_12455)
);

INVx1_ASAP7_75t_L g12456 ( 
.A(n_11922),
.Y(n_12456)
);

INVx1_ASAP7_75t_L g12457 ( 
.A(n_11978),
.Y(n_12457)
);

AOI22xp33_ASAP7_75t_L g12458 ( 
.A1(n_12102),
.A2(n_12051),
.B1(n_12064),
.B2(n_12131),
.Y(n_12458)
);

BUFx6f_ASAP7_75t_L g12459 ( 
.A(n_12073),
.Y(n_12459)
);

NAND2xp5_ASAP7_75t_L g12460 ( 
.A(n_11961),
.B(n_1854),
.Y(n_12460)
);

INVx1_ASAP7_75t_L g12461 ( 
.A(n_12000),
.Y(n_12461)
);

AOI22xp33_ASAP7_75t_L g12462 ( 
.A1(n_12131),
.A2(n_12065),
.B1(n_12082),
.B2(n_12112),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_12053),
.Y(n_12463)
);

BUFx3_ASAP7_75t_L g12464 ( 
.A(n_12090),
.Y(n_12464)
);

AOI22xp33_ASAP7_75t_SL g12465 ( 
.A1(n_12129),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.Y(n_12465)
);

INVx3_ASAP7_75t_L g12466 ( 
.A(n_11874),
.Y(n_12466)
);

OAI22xp5_ASAP7_75t_L g12467 ( 
.A1(n_12021),
.A2(n_1857),
.B1(n_1855),
.B2(n_1856),
.Y(n_12467)
);

OR2x2_ASAP7_75t_L g12468 ( 
.A(n_12085),
.B(n_1857),
.Y(n_12468)
);

AO22x1_ASAP7_75t_L g12469 ( 
.A1(n_11898),
.A2(n_1861),
.B1(n_1859),
.B2(n_1860),
.Y(n_12469)
);

AOI22xp33_ASAP7_75t_SL g12470 ( 
.A1(n_11940),
.A2(n_1862),
.B1(n_1859),
.B2(n_1861),
.Y(n_12470)
);

OAI21xp33_ASAP7_75t_L g12471 ( 
.A1(n_12072),
.A2(n_1863),
.B(n_1864),
.Y(n_12471)
);

AOI22xp33_ASAP7_75t_L g12472 ( 
.A1(n_12086),
.A2(n_1865),
.B1(n_1863),
.B2(n_1864),
.Y(n_12472)
);

CKINVDCx6p67_ASAP7_75t_R g12473 ( 
.A(n_12126),
.Y(n_12473)
);

OAI21xp5_ASAP7_75t_L g12474 ( 
.A1(n_12159),
.A2(n_1865),
.B(n_1866),
.Y(n_12474)
);

INVx1_ASAP7_75t_L g12475 ( 
.A(n_12045),
.Y(n_12475)
);

OAI22xp33_ASAP7_75t_L g12476 ( 
.A1(n_11844),
.A2(n_1868),
.B1(n_1866),
.B2(n_1867),
.Y(n_12476)
);

HB1xp67_ASAP7_75t_L g12477 ( 
.A(n_12062),
.Y(n_12477)
);

NAND2xp5_ASAP7_75t_L g12478 ( 
.A(n_12052),
.B(n_1868),
.Y(n_12478)
);

AND2x2_ASAP7_75t_L g12479 ( 
.A(n_11902),
.B(n_1870),
.Y(n_12479)
);

OAI21xp5_ASAP7_75t_SL g12480 ( 
.A1(n_12124),
.A2(n_1871),
.B(n_1872),
.Y(n_12480)
);

INVx5_ASAP7_75t_L g12481 ( 
.A(n_11862),
.Y(n_12481)
);

NAND2xp5_ASAP7_75t_L g12482 ( 
.A(n_12062),
.B(n_1872),
.Y(n_12482)
);

INVx1_ASAP7_75t_L g12483 ( 
.A(n_12068),
.Y(n_12483)
);

BUFx3_ASAP7_75t_L g12484 ( 
.A(n_12128),
.Y(n_12484)
);

CKINVDCx20_ASAP7_75t_R g12485 ( 
.A(n_11882),
.Y(n_12485)
);

OAI22xp5_ASAP7_75t_L g12486 ( 
.A1(n_11927),
.A2(n_1875),
.B1(n_1873),
.B2(n_1874),
.Y(n_12486)
);

HB1xp67_ASAP7_75t_L g12487 ( 
.A(n_12068),
.Y(n_12487)
);

HB1xp67_ASAP7_75t_L g12488 ( 
.A(n_11848),
.Y(n_12488)
);

AND2x2_ASAP7_75t_L g12489 ( 
.A(n_12173),
.B(n_1873),
.Y(n_12489)
);

CKINVDCx20_ASAP7_75t_R g12490 ( 
.A(n_12175),
.Y(n_12490)
);

OAI21xp5_ASAP7_75t_L g12491 ( 
.A1(n_11849),
.A2(n_1874),
.B(n_1876),
.Y(n_12491)
);

OAI211xp5_ASAP7_75t_L g12492 ( 
.A1(n_11849),
.A2(n_1878),
.B(n_1876),
.C(n_1877),
.Y(n_12492)
);

CKINVDCx5p33_ASAP7_75t_R g12493 ( 
.A(n_12175),
.Y(n_12493)
);

AND2x2_ASAP7_75t_L g12494 ( 
.A(n_11851),
.B(n_1878),
.Y(n_12494)
);

AOI22xp33_ASAP7_75t_L g12495 ( 
.A1(n_11926),
.A2(n_1881),
.B1(n_1879),
.B2(n_1880),
.Y(n_12495)
);

INVx2_ASAP7_75t_L g12496 ( 
.A(n_11846),
.Y(n_12496)
);

AOI22xp33_ASAP7_75t_L g12497 ( 
.A1(n_11926),
.A2(n_1881),
.B1(n_1879),
.B2(n_1880),
.Y(n_12497)
);

INVx2_ASAP7_75t_L g12498 ( 
.A(n_11846),
.Y(n_12498)
);

AND2x2_ASAP7_75t_L g12499 ( 
.A(n_11851),
.B(n_1882),
.Y(n_12499)
);

NOR2x1_ASAP7_75t_L g12500 ( 
.A(n_11933),
.B(n_1882),
.Y(n_12500)
);

BUFx2_ASAP7_75t_L g12501 ( 
.A(n_11933),
.Y(n_12501)
);

AOI22xp33_ASAP7_75t_SL g12502 ( 
.A1(n_11870),
.A2(n_1885),
.B1(n_1883),
.B2(n_1884),
.Y(n_12502)
);

OAI22xp5_ASAP7_75t_L g12503 ( 
.A1(n_11847),
.A2(n_1888),
.B1(n_1886),
.B2(n_1887),
.Y(n_12503)
);

AOI22xp33_ASAP7_75t_L g12504 ( 
.A1(n_11926),
.A2(n_1889),
.B1(n_1886),
.B2(n_1888),
.Y(n_12504)
);

INVx3_ASAP7_75t_L g12505 ( 
.A(n_11942),
.Y(n_12505)
);

INVx5_ASAP7_75t_SL g12506 ( 
.A(n_12174),
.Y(n_12506)
);

AOI22xp33_ASAP7_75t_L g12507 ( 
.A1(n_11926),
.A2(n_1891),
.B1(n_1889),
.B2(n_1890),
.Y(n_12507)
);

OAI222xp33_ASAP7_75t_L g12508 ( 
.A1(n_11870),
.A2(n_1892),
.B1(n_1894),
.B2(n_1890),
.C1(n_1891),
.C2(n_1893),
.Y(n_12508)
);

AOI22xp33_ASAP7_75t_SL g12509 ( 
.A1(n_11870),
.A2(n_1896),
.B1(n_1892),
.B2(n_1895),
.Y(n_12509)
);

INVx1_ASAP7_75t_L g12510 ( 
.A(n_11856),
.Y(n_12510)
);

AOI22xp33_ASAP7_75t_L g12511 ( 
.A1(n_11926),
.A2(n_1897),
.B1(n_1895),
.B2(n_1896),
.Y(n_12511)
);

BUFx4f_ASAP7_75t_SL g12512 ( 
.A(n_11942),
.Y(n_12512)
);

AOI22xp33_ASAP7_75t_SL g12513 ( 
.A1(n_11870),
.A2(n_1899),
.B1(n_1897),
.B2(n_1898),
.Y(n_12513)
);

AOI22xp33_ASAP7_75t_SL g12514 ( 
.A1(n_11870),
.A2(n_1900),
.B1(n_1898),
.B2(n_1899),
.Y(n_12514)
);

OAI21xp5_ASAP7_75t_SL g12515 ( 
.A1(n_11849),
.A2(n_1900),
.B(n_1902),
.Y(n_12515)
);

INVx3_ASAP7_75t_L g12516 ( 
.A(n_12179),
.Y(n_12516)
);

INVx2_ASAP7_75t_L g12517 ( 
.A(n_12334),
.Y(n_12517)
);

AND2x2_ASAP7_75t_L g12518 ( 
.A(n_12372),
.B(n_1902),
.Y(n_12518)
);

AND2x2_ASAP7_75t_L g12519 ( 
.A(n_12280),
.B(n_1903),
.Y(n_12519)
);

BUFx6f_ASAP7_75t_L g12520 ( 
.A(n_12258),
.Y(n_12520)
);

INVx1_ASAP7_75t_L g12521 ( 
.A(n_12273),
.Y(n_12521)
);

OAI21xp5_ASAP7_75t_SL g12522 ( 
.A1(n_12188),
.A2(n_1903),
.B(n_1904),
.Y(n_12522)
);

OR2x2_ASAP7_75t_SL g12523 ( 
.A(n_12313),
.B(n_1905),
.Y(n_12523)
);

INVx2_ASAP7_75t_L g12524 ( 
.A(n_12292),
.Y(n_12524)
);

AND2x2_ASAP7_75t_L g12525 ( 
.A(n_12230),
.B(n_1905),
.Y(n_12525)
);

OR2x2_ASAP7_75t_L g12526 ( 
.A(n_12320),
.B(n_1906),
.Y(n_12526)
);

INVx1_ASAP7_75t_L g12527 ( 
.A(n_12288),
.Y(n_12527)
);

AND2x2_ASAP7_75t_L g12528 ( 
.A(n_12266),
.B(n_1906),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_12301),
.Y(n_12529)
);

AND2x2_ASAP7_75t_L g12530 ( 
.A(n_12445),
.B(n_1907),
.Y(n_12530)
);

BUFx2_ASAP7_75t_L g12531 ( 
.A(n_12182),
.Y(n_12531)
);

AND2x2_ASAP7_75t_L g12532 ( 
.A(n_12209),
.B(n_1908),
.Y(n_12532)
);

NAND2xp5_ASAP7_75t_L g12533 ( 
.A(n_12217),
.B(n_1908),
.Y(n_12533)
);

AOI222xp33_ASAP7_75t_L g12534 ( 
.A1(n_12241),
.A2(n_12310),
.B1(n_12202),
.B2(n_12257),
.C1(n_12295),
.C2(n_12508),
.Y(n_12534)
);

INVx1_ASAP7_75t_L g12535 ( 
.A(n_12392),
.Y(n_12535)
);

BUFx4f_ASAP7_75t_SL g12536 ( 
.A(n_12192),
.Y(n_12536)
);

INVx3_ASAP7_75t_L g12537 ( 
.A(n_12204),
.Y(n_12537)
);

INVx1_ASAP7_75t_L g12538 ( 
.A(n_12178),
.Y(n_12538)
);

AND2x2_ASAP7_75t_L g12539 ( 
.A(n_12189),
.B(n_1909),
.Y(n_12539)
);

INVx4_ASAP7_75t_L g12540 ( 
.A(n_12248),
.Y(n_12540)
);

INVx1_ASAP7_75t_L g12541 ( 
.A(n_12197),
.Y(n_12541)
);

AND2x2_ASAP7_75t_L g12542 ( 
.A(n_12260),
.B(n_12212),
.Y(n_12542)
);

INVx1_ASAP7_75t_L g12543 ( 
.A(n_12199),
.Y(n_12543)
);

INVx3_ASAP7_75t_L g12544 ( 
.A(n_12267),
.Y(n_12544)
);

OAI22xp5_ASAP7_75t_L g12545 ( 
.A1(n_12502),
.A2(n_1911),
.B1(n_1909),
.B2(n_1910),
.Y(n_12545)
);

OR2x2_ASAP7_75t_L g12546 ( 
.A(n_12457),
.B(n_1911),
.Y(n_12546)
);

AND2x2_ASAP7_75t_L g12547 ( 
.A(n_12501),
.B(n_1912),
.Y(n_12547)
);

INVx1_ASAP7_75t_SL g12548 ( 
.A(n_12333),
.Y(n_12548)
);

AND2x2_ASAP7_75t_L g12549 ( 
.A(n_12235),
.B(n_1912),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_12383),
.B(n_1913),
.Y(n_12550)
);

INVx3_ASAP7_75t_L g12551 ( 
.A(n_12315),
.Y(n_12551)
);

INVx3_ASAP7_75t_L g12552 ( 
.A(n_12315),
.Y(n_12552)
);

HB1xp67_ASAP7_75t_L g12553 ( 
.A(n_12477),
.Y(n_12553)
);

INVx2_ASAP7_75t_L g12554 ( 
.A(n_12364),
.Y(n_12554)
);

OR2x2_ASAP7_75t_L g12555 ( 
.A(n_12194),
.B(n_1913),
.Y(n_12555)
);

INVx1_ASAP7_75t_L g12556 ( 
.A(n_12200),
.Y(n_12556)
);

INVx2_ASAP7_75t_L g12557 ( 
.A(n_12232),
.Y(n_12557)
);

INVx1_ASAP7_75t_L g12558 ( 
.A(n_12206),
.Y(n_12558)
);

INVx3_ASAP7_75t_L g12559 ( 
.A(n_12317),
.Y(n_12559)
);

INVx1_ASAP7_75t_L g12560 ( 
.A(n_12214),
.Y(n_12560)
);

BUFx3_ASAP7_75t_L g12561 ( 
.A(n_12490),
.Y(n_12561)
);

AND2x2_ASAP7_75t_L g12562 ( 
.A(n_12221),
.B(n_1914),
.Y(n_12562)
);

HB1xp67_ASAP7_75t_L g12563 ( 
.A(n_12487),
.Y(n_12563)
);

NAND2xp5_ASAP7_75t_L g12564 ( 
.A(n_12180),
.B(n_1914),
.Y(n_12564)
);

HB1xp67_ASAP7_75t_L g12565 ( 
.A(n_12208),
.Y(n_12565)
);

INVx3_ASAP7_75t_L g12566 ( 
.A(n_12291),
.Y(n_12566)
);

OR2x2_ASAP7_75t_L g12567 ( 
.A(n_12496),
.B(n_1915),
.Y(n_12567)
);

AND2x2_ASAP7_75t_L g12568 ( 
.A(n_12234),
.B(n_1915),
.Y(n_12568)
);

INVx2_ASAP7_75t_L g12569 ( 
.A(n_12349),
.Y(n_12569)
);

AOI22xp33_ASAP7_75t_L g12570 ( 
.A1(n_12509),
.A2(n_1918),
.B1(n_1916),
.B2(n_1917),
.Y(n_12570)
);

INVx1_ASAP7_75t_L g12571 ( 
.A(n_12220),
.Y(n_12571)
);

INVx1_ASAP7_75t_L g12572 ( 
.A(n_12226),
.Y(n_12572)
);

AOI22xp33_ASAP7_75t_L g12573 ( 
.A1(n_12513),
.A2(n_1919),
.B1(n_1916),
.B2(n_1917),
.Y(n_12573)
);

INVx2_ASAP7_75t_L g12574 ( 
.A(n_12349),
.Y(n_12574)
);

AND2x2_ASAP7_75t_L g12575 ( 
.A(n_12498),
.B(n_1919),
.Y(n_12575)
);

INVxp67_ASAP7_75t_L g12576 ( 
.A(n_12330),
.Y(n_12576)
);

OR2x6_ASAP7_75t_L g12577 ( 
.A(n_12378),
.B(n_1920),
.Y(n_12577)
);

HB1xp67_ASAP7_75t_L g12578 ( 
.A(n_12254),
.Y(n_12578)
);

NAND2x1_ASAP7_75t_L g12579 ( 
.A(n_12401),
.B(n_12454),
.Y(n_12579)
);

INVx3_ASAP7_75t_L g12580 ( 
.A(n_12360),
.Y(n_12580)
);

INVx2_ASAP7_75t_SL g12581 ( 
.A(n_12248),
.Y(n_12581)
);

INVx2_ASAP7_75t_L g12582 ( 
.A(n_12401),
.Y(n_12582)
);

AND2x2_ASAP7_75t_L g12583 ( 
.A(n_12275),
.B(n_1920),
.Y(n_12583)
);

INVx4_ASAP7_75t_L g12584 ( 
.A(n_12248),
.Y(n_12584)
);

AOI22xp33_ASAP7_75t_L g12585 ( 
.A1(n_12514),
.A2(n_1923),
.B1(n_1921),
.B2(n_1922),
.Y(n_12585)
);

AND2x4_ASAP7_75t_L g12586 ( 
.A(n_12181),
.B(n_1921),
.Y(n_12586)
);

OR2x2_ASAP7_75t_L g12587 ( 
.A(n_12456),
.B(n_1923),
.Y(n_12587)
);

AND2x2_ASAP7_75t_L g12588 ( 
.A(n_12323),
.B(n_1924),
.Y(n_12588)
);

HB1xp67_ASAP7_75t_L g12589 ( 
.A(n_12420),
.Y(n_12589)
);

INVx2_ASAP7_75t_L g12590 ( 
.A(n_12505),
.Y(n_12590)
);

AOI21xp33_ASAP7_75t_L g12591 ( 
.A1(n_12332),
.A2(n_1925),
.B(n_1926),
.Y(n_12591)
);

AND2x2_ASAP7_75t_L g12592 ( 
.A(n_12279),
.B(n_12319),
.Y(n_12592)
);

AND2x2_ASAP7_75t_L g12593 ( 
.A(n_12348),
.B(n_1925),
.Y(n_12593)
);

INVx2_ASAP7_75t_SL g12594 ( 
.A(n_12512),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_12389),
.Y(n_12595)
);

AND2x2_ASAP7_75t_L g12596 ( 
.A(n_12352),
.B(n_1927),
.Y(n_12596)
);

INVx2_ASAP7_75t_L g12597 ( 
.A(n_12389),
.Y(n_12597)
);

INVx2_ASAP7_75t_L g12598 ( 
.A(n_12390),
.Y(n_12598)
);

NAND2xp5_ASAP7_75t_L g12599 ( 
.A(n_12475),
.B(n_1927),
.Y(n_12599)
);

INVx2_ASAP7_75t_L g12600 ( 
.A(n_12390),
.Y(n_12600)
);

AND2x2_ASAP7_75t_L g12601 ( 
.A(n_12417),
.B(n_1928),
.Y(n_12601)
);

AND2x2_ASAP7_75t_L g12602 ( 
.A(n_12353),
.B(n_12377),
.Y(n_12602)
);

INVx2_ASAP7_75t_L g12603 ( 
.A(n_12459),
.Y(n_12603)
);

AND2x2_ASAP7_75t_L g12604 ( 
.A(n_12428),
.B(n_1928),
.Y(n_12604)
);

INVx1_ASAP7_75t_L g12605 ( 
.A(n_12243),
.Y(n_12605)
);

INVx1_ASAP7_75t_L g12606 ( 
.A(n_12262),
.Y(n_12606)
);

AND2x2_ASAP7_75t_L g12607 ( 
.A(n_12272),
.B(n_1929),
.Y(n_12607)
);

AND2x4_ASAP7_75t_SL g12608 ( 
.A(n_12294),
.B(n_12375),
.Y(n_12608)
);

AND2x2_ASAP7_75t_L g12609 ( 
.A(n_12272),
.B(n_1929),
.Y(n_12609)
);

AND2x2_ASAP7_75t_L g12610 ( 
.A(n_12338),
.B(n_1930),
.Y(n_12610)
);

OAI22xp33_ASAP7_75t_L g12611 ( 
.A1(n_12205),
.A2(n_12269),
.B1(n_12223),
.B2(n_12252),
.Y(n_12611)
);

AND2x2_ASAP7_75t_L g12612 ( 
.A(n_12338),
.B(n_1930),
.Y(n_12612)
);

INVx3_ASAP7_75t_L g12613 ( 
.A(n_12459),
.Y(n_12613)
);

AND2x2_ASAP7_75t_L g12614 ( 
.A(n_12506),
.B(n_1931),
.Y(n_12614)
);

INVx2_ASAP7_75t_L g12615 ( 
.A(n_12464),
.Y(n_12615)
);

AND2x2_ASAP7_75t_L g12616 ( 
.A(n_12506),
.B(n_1931),
.Y(n_12616)
);

INVx1_ASAP7_75t_L g12617 ( 
.A(n_12268),
.Y(n_12617)
);

INVx2_ASAP7_75t_L g12618 ( 
.A(n_12466),
.Y(n_12618)
);

NOR2xp33_ASAP7_75t_R g12619 ( 
.A(n_12493),
.B(n_1932),
.Y(n_12619)
);

AOI22xp33_ASAP7_75t_L g12620 ( 
.A1(n_12215),
.A2(n_1934),
.B1(n_1932),
.B2(n_1933),
.Y(n_12620)
);

INVx1_ASAP7_75t_L g12621 ( 
.A(n_12278),
.Y(n_12621)
);

INVx2_ASAP7_75t_SL g12622 ( 
.A(n_12343),
.Y(n_12622)
);

AND2x2_ASAP7_75t_L g12623 ( 
.A(n_12370),
.B(n_1933),
.Y(n_12623)
);

AND2x2_ASAP7_75t_L g12624 ( 
.A(n_12461),
.B(n_12484),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12281),
.Y(n_12625)
);

AND2x2_ASAP7_75t_L g12626 ( 
.A(n_12425),
.B(n_12494),
.Y(n_12626)
);

HB1xp67_ASAP7_75t_L g12627 ( 
.A(n_12440),
.Y(n_12627)
);

INVx2_ASAP7_75t_L g12628 ( 
.A(n_12366),
.Y(n_12628)
);

AND2x2_ASAP7_75t_L g12629 ( 
.A(n_12499),
.B(n_1934),
.Y(n_12629)
);

INVx2_ASAP7_75t_L g12630 ( 
.A(n_12426),
.Y(n_12630)
);

INVx2_ASAP7_75t_L g12631 ( 
.A(n_12435),
.Y(n_12631)
);

AOI22xp33_ASAP7_75t_L g12632 ( 
.A1(n_12491),
.A2(n_1937),
.B1(n_1935),
.B2(n_1936),
.Y(n_12632)
);

NOR2xp33_ASAP7_75t_L g12633 ( 
.A(n_12355),
.B(n_1935),
.Y(n_12633)
);

INVx3_ASAP7_75t_L g12634 ( 
.A(n_12227),
.Y(n_12634)
);

INVx1_ASAP7_75t_L g12635 ( 
.A(n_12287),
.Y(n_12635)
);

HB1xp67_ASAP7_75t_L g12636 ( 
.A(n_12483),
.Y(n_12636)
);

INVx1_ASAP7_75t_L g12637 ( 
.A(n_12289),
.Y(n_12637)
);

AND2x2_ASAP7_75t_L g12638 ( 
.A(n_12447),
.B(n_1936),
.Y(n_12638)
);

OAI22xp5_ASAP7_75t_L g12639 ( 
.A1(n_12495),
.A2(n_1939),
.B1(n_1937),
.B2(n_1938),
.Y(n_12639)
);

INVx1_ASAP7_75t_L g12640 ( 
.A(n_12309),
.Y(n_12640)
);

NAND2xp5_ASAP7_75t_L g12641 ( 
.A(n_12299),
.B(n_1938),
.Y(n_12641)
);

INVx1_ASAP7_75t_L g12642 ( 
.A(n_12322),
.Y(n_12642)
);

INVx1_ASAP7_75t_L g12643 ( 
.A(n_12327),
.Y(n_12643)
);

OAI22xp5_ASAP7_75t_L g12644 ( 
.A1(n_12497),
.A2(n_1941),
.B1(n_1939),
.B2(n_1940),
.Y(n_12644)
);

INVx2_ASAP7_75t_L g12645 ( 
.A(n_12446),
.Y(n_12645)
);

AND2x2_ASAP7_75t_L g12646 ( 
.A(n_12453),
.B(n_1940),
.Y(n_12646)
);

AND2x2_ASAP7_75t_L g12647 ( 
.A(n_12436),
.B(n_1941),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_12336),
.Y(n_12648)
);

BUFx3_ASAP7_75t_L g12649 ( 
.A(n_12261),
.Y(n_12649)
);

OAI22xp5_ASAP7_75t_L g12650 ( 
.A1(n_12504),
.A2(n_1944),
.B1(n_1942),
.B2(n_1943),
.Y(n_12650)
);

BUFx2_ASAP7_75t_L g12651 ( 
.A(n_12434),
.Y(n_12651)
);

AND2x2_ASAP7_75t_L g12652 ( 
.A(n_12222),
.B(n_1942),
.Y(n_12652)
);

AND2x2_ASAP7_75t_L g12653 ( 
.A(n_12239),
.B(n_1943),
.Y(n_12653)
);

AND2x2_ASAP7_75t_L g12654 ( 
.A(n_12463),
.B(n_1945),
.Y(n_12654)
);

INVx2_ASAP7_75t_L g12655 ( 
.A(n_12481),
.Y(n_12655)
);

INVx1_ASAP7_75t_L g12656 ( 
.A(n_12339),
.Y(n_12656)
);

INVx1_ASAP7_75t_L g12657 ( 
.A(n_12340),
.Y(n_12657)
);

AOI22xp33_ASAP7_75t_L g12658 ( 
.A1(n_12236),
.A2(n_1948),
.B1(n_1946),
.B2(n_1947),
.Y(n_12658)
);

INVx1_ASAP7_75t_L g12659 ( 
.A(n_12344),
.Y(n_12659)
);

INVx2_ASAP7_75t_L g12660 ( 
.A(n_12481),
.Y(n_12660)
);

AND2x2_ASAP7_75t_L g12661 ( 
.A(n_12473),
.B(n_1946),
.Y(n_12661)
);

AOI22xp33_ASAP7_75t_L g12662 ( 
.A1(n_12507),
.A2(n_1951),
.B1(n_1949),
.B2(n_1950),
.Y(n_12662)
);

INVx2_ASAP7_75t_L g12663 ( 
.A(n_12481),
.Y(n_12663)
);

INVx1_ASAP7_75t_L g12664 ( 
.A(n_12345),
.Y(n_12664)
);

INVx1_ASAP7_75t_SL g12665 ( 
.A(n_12302),
.Y(n_12665)
);

INVxp67_ASAP7_75t_SL g12666 ( 
.A(n_12500),
.Y(n_12666)
);

INVx2_ASAP7_75t_L g12667 ( 
.A(n_12485),
.Y(n_12667)
);

AND2x2_ASAP7_75t_L g12668 ( 
.A(n_12293),
.B(n_1950),
.Y(n_12668)
);

NAND2xp5_ASAP7_75t_L g12669 ( 
.A(n_12316),
.B(n_1951),
.Y(n_12669)
);

AND2x2_ASAP7_75t_L g12670 ( 
.A(n_12314),
.B(n_1952),
.Y(n_12670)
);

OAI22xp5_ASAP7_75t_L g12671 ( 
.A1(n_12511),
.A2(n_1954),
.B1(n_1952),
.B2(n_1953),
.Y(n_12671)
);

BUFx6f_ASAP7_75t_L g12672 ( 
.A(n_12238),
.Y(n_12672)
);

AND2x2_ASAP7_75t_L g12673 ( 
.A(n_12462),
.B(n_1953),
.Y(n_12673)
);

INVx1_ASAP7_75t_L g12674 ( 
.A(n_12350),
.Y(n_12674)
);

NAND2xp5_ASAP7_75t_L g12675 ( 
.A(n_12419),
.B(n_1954),
.Y(n_12675)
);

AND2x2_ASAP7_75t_L g12676 ( 
.A(n_12395),
.B(n_1955),
.Y(n_12676)
);

AND2x2_ASAP7_75t_L g12677 ( 
.A(n_12362),
.B(n_1955),
.Y(n_12677)
);

INVx1_ASAP7_75t_L g12678 ( 
.A(n_12351),
.Y(n_12678)
);

INVx2_ASAP7_75t_L g12679 ( 
.A(n_12489),
.Y(n_12679)
);

AND2x2_ASAP7_75t_L g12680 ( 
.A(n_12290),
.B(n_1956),
.Y(n_12680)
);

INVx2_ASAP7_75t_L g12681 ( 
.A(n_12412),
.Y(n_12681)
);

BUFx2_ASAP7_75t_L g12682 ( 
.A(n_12363),
.Y(n_12682)
);

OR2x2_ASAP7_75t_L g12683 ( 
.A(n_12341),
.B(n_12385),
.Y(n_12683)
);

INVx2_ASAP7_75t_L g12684 ( 
.A(n_12422),
.Y(n_12684)
);

AND2x2_ASAP7_75t_L g12685 ( 
.A(n_12413),
.B(n_1957),
.Y(n_12685)
);

INVx2_ASAP7_75t_L g12686 ( 
.A(n_12432),
.Y(n_12686)
);

INVx2_ASAP7_75t_L g12687 ( 
.A(n_12433),
.Y(n_12687)
);

INVx1_ASAP7_75t_L g12688 ( 
.A(n_12361),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_12510),
.Y(n_12689)
);

AND2x2_ASAP7_75t_L g12690 ( 
.A(n_12442),
.B(n_1957),
.Y(n_12690)
);

INVx2_ASAP7_75t_L g12691 ( 
.A(n_12347),
.Y(n_12691)
);

AND2x2_ASAP7_75t_L g12692 ( 
.A(n_12444),
.B(n_1958),
.Y(n_12692)
);

BUFx3_ASAP7_75t_L g12693 ( 
.A(n_12394),
.Y(n_12693)
);

AND2x2_ASAP7_75t_L g12694 ( 
.A(n_12458),
.B(n_12450),
.Y(n_12694)
);

AOI22xp33_ASAP7_75t_L g12695 ( 
.A1(n_12177),
.A2(n_1961),
.B1(n_1959),
.B2(n_1960),
.Y(n_12695)
);

AND2x4_ASAP7_75t_SL g12696 ( 
.A(n_12479),
.B(n_1959),
.Y(n_12696)
);

INVx1_ASAP7_75t_L g12697 ( 
.A(n_12369),
.Y(n_12697)
);

BUFx2_ASAP7_75t_L g12698 ( 
.A(n_12430),
.Y(n_12698)
);

AND2x2_ASAP7_75t_L g12699 ( 
.A(n_12256),
.B(n_1960),
.Y(n_12699)
);

AND2x2_ASAP7_75t_L g12700 ( 
.A(n_12298),
.B(n_1961),
.Y(n_12700)
);

AND2x4_ASAP7_75t_L g12701 ( 
.A(n_12421),
.B(n_1962),
.Y(n_12701)
);

NOR2x1_ASAP7_75t_L g12702 ( 
.A(n_12264),
.B(n_1962),
.Y(n_12702)
);

NOR2xp33_ASAP7_75t_L g12703 ( 
.A(n_12265),
.B(n_1963),
.Y(n_12703)
);

INVx1_ASAP7_75t_L g12704 ( 
.A(n_12373),
.Y(n_12704)
);

AND2x2_ASAP7_75t_L g12705 ( 
.A(n_12403),
.B(n_1963),
.Y(n_12705)
);

INVx1_ASAP7_75t_SL g12706 ( 
.A(n_12259),
.Y(n_12706)
);

AOI22xp33_ASAP7_75t_L g12707 ( 
.A1(n_12296),
.A2(n_1966),
.B1(n_1964),
.B2(n_1965),
.Y(n_12707)
);

AOI22xp33_ASAP7_75t_L g12708 ( 
.A1(n_12242),
.A2(n_1966),
.B1(n_1964),
.B2(n_1965),
.Y(n_12708)
);

NAND2xp5_ASAP7_75t_L g12709 ( 
.A(n_12184),
.B(n_1968),
.Y(n_12709)
);

INVx2_ASAP7_75t_L g12710 ( 
.A(n_12376),
.Y(n_12710)
);

AND2x4_ASAP7_75t_L g12711 ( 
.A(n_12455),
.B(n_1969),
.Y(n_12711)
);

INVx1_ASAP7_75t_L g12712 ( 
.A(n_12286),
.Y(n_12712)
);

INVx1_ASAP7_75t_L g12713 ( 
.A(n_12303),
.Y(n_12713)
);

INVx1_ASAP7_75t_L g12714 ( 
.A(n_12276),
.Y(n_12714)
);

INVx3_ASAP7_75t_L g12715 ( 
.A(n_12468),
.Y(n_12715)
);

INVx1_ASAP7_75t_L g12716 ( 
.A(n_12285),
.Y(n_12716)
);

INVxp67_ASAP7_75t_L g12717 ( 
.A(n_12186),
.Y(n_12717)
);

BUFx3_ASAP7_75t_L g12718 ( 
.A(n_12308),
.Y(n_12718)
);

INVx1_ASAP7_75t_L g12719 ( 
.A(n_12482),
.Y(n_12719)
);

INVx3_ASAP7_75t_L g12720 ( 
.A(n_12410),
.Y(n_12720)
);

INVx1_ASAP7_75t_L g12721 ( 
.A(n_12418),
.Y(n_12721)
);

BUFx2_ASAP7_75t_L g12722 ( 
.A(n_12449),
.Y(n_12722)
);

INVx2_ASAP7_75t_SL g12723 ( 
.A(n_12478),
.Y(n_12723)
);

BUFx3_ASAP7_75t_L g12724 ( 
.A(n_12424),
.Y(n_12724)
);

OR2x2_ASAP7_75t_L g12725 ( 
.A(n_12365),
.B(n_1969),
.Y(n_12725)
);

INVx2_ASAP7_75t_L g12726 ( 
.A(n_12488),
.Y(n_12726)
);

INVx1_ASAP7_75t_L g12727 ( 
.A(n_12409),
.Y(n_12727)
);

AND2x2_ASAP7_75t_L g12728 ( 
.A(n_12384),
.B(n_1970),
.Y(n_12728)
);

INVx2_ASAP7_75t_L g12729 ( 
.A(n_12460),
.Y(n_12729)
);

INVx2_ASAP7_75t_L g12730 ( 
.A(n_12359),
.Y(n_12730)
);

INVx2_ASAP7_75t_SL g12731 ( 
.A(n_12469),
.Y(n_12731)
);

INVx1_ASAP7_75t_L g12732 ( 
.A(n_12431),
.Y(n_12732)
);

AND2x2_ASAP7_75t_L g12733 ( 
.A(n_12439),
.B(n_1971),
.Y(n_12733)
);

INVx1_ASAP7_75t_L g12734 ( 
.A(n_12297),
.Y(n_12734)
);

AND2x2_ASAP7_75t_L g12735 ( 
.A(n_12474),
.B(n_1973),
.Y(n_12735)
);

INVx1_ASAP7_75t_L g12736 ( 
.A(n_12187),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_12480),
.B(n_1973),
.Y(n_12737)
);

INVx1_ASAP7_75t_SL g12738 ( 
.A(n_12193),
.Y(n_12738)
);

NAND2x1_ASAP7_75t_L g12739 ( 
.A(n_12219),
.B(n_1974),
.Y(n_12739)
);

INVx3_ASAP7_75t_L g12740 ( 
.A(n_12225),
.Y(n_12740)
);

AND2x2_ASAP7_75t_L g12741 ( 
.A(n_12307),
.B(n_12368),
.Y(n_12741)
);

INVx2_ASAP7_75t_L g12742 ( 
.A(n_12404),
.Y(n_12742)
);

AND2x2_ASAP7_75t_L g12743 ( 
.A(n_12402),
.B(n_1974),
.Y(n_12743)
);

AND2x2_ASAP7_75t_L g12744 ( 
.A(n_12503),
.B(n_1975),
.Y(n_12744)
);

NAND2xp5_ASAP7_75t_L g12745 ( 
.A(n_12515),
.B(n_1975),
.Y(n_12745)
);

INVx1_ASAP7_75t_L g12746 ( 
.A(n_12396),
.Y(n_12746)
);

AND2x2_ASAP7_75t_L g12747 ( 
.A(n_12471),
.B(n_1976),
.Y(n_12747)
);

AOI22xp33_ASAP7_75t_L g12748 ( 
.A1(n_12201),
.A2(n_1978),
.B1(n_1976),
.B2(n_1977),
.Y(n_12748)
);

OR2x2_ASAP7_75t_L g12749 ( 
.A(n_12415),
.B(n_1977),
.Y(n_12749)
);

NAND2xp5_ASAP7_75t_L g12750 ( 
.A(n_12408),
.B(n_1978),
.Y(n_12750)
);

INVx1_ASAP7_75t_L g12751 ( 
.A(n_12486),
.Y(n_12751)
);

AND2x2_ASAP7_75t_L g12752 ( 
.A(n_12277),
.B(n_1979),
.Y(n_12752)
);

INVx1_ASAP7_75t_L g12753 ( 
.A(n_12467),
.Y(n_12753)
);

NOR2xp33_ASAP7_75t_L g12754 ( 
.A(n_12451),
.B(n_1979),
.Y(n_12754)
);

OAI22xp5_ASAP7_75t_L g12755 ( 
.A1(n_12191),
.A2(n_1982),
.B1(n_1980),
.B2(n_1981),
.Y(n_12755)
);

NAND2xp5_ASAP7_75t_L g12756 ( 
.A(n_12329),
.B(n_1981),
.Y(n_12756)
);

AND2x2_ASAP7_75t_L g12757 ( 
.A(n_12354),
.B(n_1982),
.Y(n_12757)
);

INVx2_ASAP7_75t_L g12758 ( 
.A(n_12190),
.Y(n_12758)
);

HB1xp67_ASAP7_75t_L g12759 ( 
.A(n_12326),
.Y(n_12759)
);

HB1xp67_ASAP7_75t_L g12760 ( 
.A(n_12357),
.Y(n_12760)
);

INVx1_ASAP7_75t_L g12761 ( 
.A(n_12476),
.Y(n_12761)
);

AND2x2_ASAP7_75t_L g12762 ( 
.A(n_12465),
.B(n_1983),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_12282),
.B(n_1983),
.Y(n_12763)
);

INVxp67_ASAP7_75t_L g12764 ( 
.A(n_12492),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_12321),
.B(n_1984),
.Y(n_12765)
);

AOI22xp33_ASAP7_75t_L g12766 ( 
.A1(n_12371),
.A2(n_1987),
.B1(n_1985),
.B2(n_1986),
.Y(n_12766)
);

INVx1_ASAP7_75t_L g12767 ( 
.A(n_12250),
.Y(n_12767)
);

HB1xp67_ASAP7_75t_L g12768 ( 
.A(n_12337),
.Y(n_12768)
);

OR2x2_ASAP7_75t_L g12769 ( 
.A(n_12731),
.B(n_12311),
.Y(n_12769)
);

INVx2_ASAP7_75t_L g12770 ( 
.A(n_12561),
.Y(n_12770)
);

AND2x2_ASAP7_75t_L g12771 ( 
.A(n_12548),
.B(n_12393),
.Y(n_12771)
);

AND2x2_ASAP7_75t_L g12772 ( 
.A(n_12531),
.B(n_12342),
.Y(n_12772)
);

INVx1_ASAP7_75t_L g12773 ( 
.A(n_12589),
.Y(n_12773)
);

AOI22xp33_ASAP7_75t_L g12774 ( 
.A1(n_12759),
.A2(n_12233),
.B1(n_12210),
.B2(n_12429),
.Y(n_12774)
);

INVx5_ASAP7_75t_L g12775 ( 
.A(n_12520),
.Y(n_12775)
);

INVx2_ASAP7_75t_SL g12776 ( 
.A(n_12520),
.Y(n_12776)
);

INVx2_ASAP7_75t_L g12777 ( 
.A(n_12634),
.Y(n_12777)
);

INVx2_ASAP7_75t_SL g12778 ( 
.A(n_12516),
.Y(n_12778)
);

AND2x2_ASAP7_75t_L g12779 ( 
.A(n_12580),
.B(n_12427),
.Y(n_12779)
);

INVx2_ASAP7_75t_L g12780 ( 
.A(n_12540),
.Y(n_12780)
);

INVx1_ASAP7_75t_L g12781 ( 
.A(n_12627),
.Y(n_12781)
);

BUFx3_ASAP7_75t_L g12782 ( 
.A(n_12536),
.Y(n_12782)
);

HB1xp67_ASAP7_75t_L g12783 ( 
.A(n_12565),
.Y(n_12783)
);

AND2x4_ASAP7_75t_L g12784 ( 
.A(n_12551),
.B(n_12379),
.Y(n_12784)
);

INVx2_ASAP7_75t_L g12785 ( 
.A(n_12584),
.Y(n_12785)
);

INVx2_ASAP7_75t_L g12786 ( 
.A(n_12552),
.Y(n_12786)
);

AND2x2_ASAP7_75t_L g12787 ( 
.A(n_12542),
.B(n_12438),
.Y(n_12787)
);

AND2x2_ASAP7_75t_L g12788 ( 
.A(n_12559),
.B(n_12231),
.Y(n_12788)
);

INVx2_ASAP7_75t_L g12789 ( 
.A(n_12544),
.Y(n_12789)
);

AND2x2_ASAP7_75t_L g12790 ( 
.A(n_12537),
.B(n_12213),
.Y(n_12790)
);

INVx1_ASAP7_75t_L g12791 ( 
.A(n_12636),
.Y(n_12791)
);

AND2x4_ASAP7_75t_L g12792 ( 
.A(n_12608),
.B(n_12407),
.Y(n_12792)
);

INVx2_ASAP7_75t_L g12793 ( 
.A(n_12672),
.Y(n_12793)
);

AND2x2_ASAP7_75t_L g12794 ( 
.A(n_12651),
.B(n_12195),
.Y(n_12794)
);

AOI22xp33_ASAP7_75t_L g12795 ( 
.A1(n_12694),
.A2(n_12400),
.B1(n_12331),
.B2(n_12240),
.Y(n_12795)
);

AND2x2_ASAP7_75t_L g12796 ( 
.A(n_12645),
.B(n_12470),
.Y(n_12796)
);

INVx3_ASAP7_75t_L g12797 ( 
.A(n_12649),
.Y(n_12797)
);

AND2x4_ASAP7_75t_L g12798 ( 
.A(n_12581),
.B(n_12185),
.Y(n_12798)
);

AND2x4_ASAP7_75t_SL g12799 ( 
.A(n_12566),
.B(n_12452),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12553),
.Y(n_12800)
);

INVx1_ASAP7_75t_L g12801 ( 
.A(n_12563),
.Y(n_12801)
);

INVx1_ASAP7_75t_L g12802 ( 
.A(n_12521),
.Y(n_12802)
);

AND2x2_ASAP7_75t_L g12803 ( 
.A(n_12524),
.B(n_12306),
.Y(n_12803)
);

OR2x2_ASAP7_75t_L g12804 ( 
.A(n_12730),
.B(n_12211),
.Y(n_12804)
);

OR2x2_ASAP7_75t_L g12805 ( 
.A(n_12734),
.B(n_12300),
.Y(n_12805)
);

OAI22xp33_ASAP7_75t_L g12806 ( 
.A1(n_12740),
.A2(n_12388),
.B1(n_12381),
.B2(n_12216),
.Y(n_12806)
);

BUFx2_ASAP7_75t_L g12807 ( 
.A(n_12666),
.Y(n_12807)
);

INVx4_ASAP7_75t_L g12808 ( 
.A(n_12577),
.Y(n_12808)
);

INVx1_ASAP7_75t_L g12809 ( 
.A(n_12527),
.Y(n_12809)
);

NAND2xp5_ASAP7_75t_L g12810 ( 
.A(n_12706),
.B(n_12423),
.Y(n_12810)
);

HB1xp67_ASAP7_75t_L g12811 ( 
.A(n_12578),
.Y(n_12811)
);

INVx1_ASAP7_75t_L g12812 ( 
.A(n_12529),
.Y(n_12812)
);

AND2x2_ASAP7_75t_L g12813 ( 
.A(n_12590),
.B(n_12304),
.Y(n_12813)
);

OR2x2_ASAP7_75t_L g12814 ( 
.A(n_12760),
.B(n_12328),
.Y(n_12814)
);

INVx2_ASAP7_75t_L g12815 ( 
.A(n_12672),
.Y(n_12815)
);

INVx1_ASAP7_75t_L g12816 ( 
.A(n_12682),
.Y(n_12816)
);

INVx2_ASAP7_75t_L g12817 ( 
.A(n_12631),
.Y(n_12817)
);

INVx1_ASAP7_75t_L g12818 ( 
.A(n_12705),
.Y(n_12818)
);

AO21x2_ASAP7_75t_L g12819 ( 
.A1(n_12533),
.A2(n_12387),
.B(n_12324),
.Y(n_12819)
);

AND2x2_ASAP7_75t_L g12820 ( 
.A(n_12517),
.B(n_12448),
.Y(n_12820)
);

INVx1_ASAP7_75t_L g12821 ( 
.A(n_12546),
.Y(n_12821)
);

INVx1_ASAP7_75t_L g12822 ( 
.A(n_12710),
.Y(n_12822)
);

INVx1_ASAP7_75t_L g12823 ( 
.A(n_12538),
.Y(n_12823)
);

HB1xp67_ASAP7_75t_L g12824 ( 
.A(n_12525),
.Y(n_12824)
);

INVx1_ASAP7_75t_L g12825 ( 
.A(n_12541),
.Y(n_12825)
);

INVx1_ASAP7_75t_L g12826 ( 
.A(n_12543),
.Y(n_12826)
);

INVx2_ASAP7_75t_L g12827 ( 
.A(n_12630),
.Y(n_12827)
);

INVx2_ASAP7_75t_SL g12828 ( 
.A(n_12579),
.Y(n_12828)
);

AND2x2_ASAP7_75t_L g12829 ( 
.A(n_12626),
.B(n_12183),
.Y(n_12829)
);

HB1xp67_ASAP7_75t_L g12830 ( 
.A(n_12722),
.Y(n_12830)
);

INVx2_ASAP7_75t_L g12831 ( 
.A(n_12613),
.Y(n_12831)
);

NOR2x1_ASAP7_75t_L g12832 ( 
.A(n_12702),
.B(n_12245),
.Y(n_12832)
);

AND2x2_ASAP7_75t_L g12833 ( 
.A(n_12569),
.B(n_12312),
.Y(n_12833)
);

INVx1_ASAP7_75t_L g12834 ( 
.A(n_12556),
.Y(n_12834)
);

AND2x2_ASAP7_75t_L g12835 ( 
.A(n_12574),
.B(n_12203),
.Y(n_12835)
);

NAND2xp5_ASAP7_75t_L g12836 ( 
.A(n_12534),
.B(n_12218),
.Y(n_12836)
);

BUFx3_ASAP7_75t_L g12837 ( 
.A(n_12594),
.Y(n_12837)
);

INVx2_ASAP7_75t_SL g12838 ( 
.A(n_12655),
.Y(n_12838)
);

OR2x2_ASAP7_75t_SL g12839 ( 
.A(n_12582),
.B(n_12255),
.Y(n_12839)
);

AND2x2_ASAP7_75t_L g12840 ( 
.A(n_12667),
.B(n_12346),
.Y(n_12840)
);

INVx1_ASAP7_75t_L g12841 ( 
.A(n_12558),
.Y(n_12841)
);

INVxp67_ASAP7_75t_SL g12842 ( 
.A(n_12576),
.Y(n_12842)
);

BUFx3_ASAP7_75t_L g12843 ( 
.A(n_12693),
.Y(n_12843)
);

INVxp67_ASAP7_75t_SL g12844 ( 
.A(n_12718),
.Y(n_12844)
);

AND2x6_ASAP7_75t_L g12845 ( 
.A(n_12665),
.B(n_12244),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_12738),
.B(n_12224),
.Y(n_12846)
);

INVx1_ASAP7_75t_L g12847 ( 
.A(n_12560),
.Y(n_12847)
);

INVx2_ASAP7_75t_L g12848 ( 
.A(n_12622),
.Y(n_12848)
);

AND4x1_ASAP7_75t_L g12849 ( 
.A(n_12766),
.B(n_12391),
.C(n_12229),
.D(n_12416),
.Y(n_12849)
);

INVx2_ASAP7_75t_L g12850 ( 
.A(n_12557),
.Y(n_12850)
);

NAND2xp5_ASAP7_75t_L g12851 ( 
.A(n_12764),
.B(n_12196),
.Y(n_12851)
);

INVx2_ASAP7_75t_L g12852 ( 
.A(n_12554),
.Y(n_12852)
);

AND2x2_ASAP7_75t_L g12853 ( 
.A(n_12628),
.B(n_12472),
.Y(n_12853)
);

INVx2_ASAP7_75t_L g12854 ( 
.A(n_12595),
.Y(n_12854)
);

INVx2_ASAP7_75t_L g12855 ( 
.A(n_12597),
.Y(n_12855)
);

NOR2xp33_ASAP7_75t_L g12856 ( 
.A(n_12698),
.B(n_12246),
.Y(n_12856)
);

NAND2xp5_ASAP7_75t_L g12857 ( 
.A(n_12611),
.B(n_12251),
.Y(n_12857)
);

INVx2_ASAP7_75t_L g12858 ( 
.A(n_12598),
.Y(n_12858)
);

HB1xp67_ASAP7_75t_L g12859 ( 
.A(n_12660),
.Y(n_12859)
);

BUFx2_ASAP7_75t_L g12860 ( 
.A(n_12577),
.Y(n_12860)
);

OR2x2_ASAP7_75t_L g12861 ( 
.A(n_12523),
.B(n_12247),
.Y(n_12861)
);

AOI221xp5_ASAP7_75t_L g12862 ( 
.A1(n_12522),
.A2(n_12249),
.B1(n_12284),
.B2(n_12237),
.C(n_12198),
.Y(n_12862)
);

AND2x2_ASAP7_75t_L g12863 ( 
.A(n_12600),
.B(n_12441),
.Y(n_12863)
);

INVx1_ASAP7_75t_L g12864 ( 
.A(n_12571),
.Y(n_12864)
);

AND2x2_ASAP7_75t_L g12865 ( 
.A(n_12603),
.B(n_12615),
.Y(n_12865)
);

OR2x2_ASAP7_75t_L g12866 ( 
.A(n_12526),
.B(n_12761),
.Y(n_12866)
);

AND2x2_ASAP7_75t_L g12867 ( 
.A(n_12592),
.B(n_12325),
.Y(n_12867)
);

INVx1_ASAP7_75t_L g12868 ( 
.A(n_12572),
.Y(n_12868)
);

AND2x2_ASAP7_75t_L g12869 ( 
.A(n_12602),
.B(n_12380),
.Y(n_12869)
);

AND2x2_ASAP7_75t_L g12870 ( 
.A(n_12618),
.B(n_12283),
.Y(n_12870)
);

INVx1_ASAP7_75t_L g12871 ( 
.A(n_12605),
.Y(n_12871)
);

INVx3_ASAP7_75t_SL g12872 ( 
.A(n_12586),
.Y(n_12872)
);

BUFx2_ASAP7_75t_L g12873 ( 
.A(n_12663),
.Y(n_12873)
);

NAND2xp5_ASAP7_75t_L g12874 ( 
.A(n_12717),
.B(n_12207),
.Y(n_12874)
);

BUFx6f_ASAP7_75t_L g12875 ( 
.A(n_12661),
.Y(n_12875)
);

INVx1_ASAP7_75t_L g12876 ( 
.A(n_12606),
.Y(n_12876)
);

OR2x2_ASAP7_75t_L g12877 ( 
.A(n_12715),
.B(n_12367),
.Y(n_12877)
);

AND2x2_ASAP7_75t_L g12878 ( 
.A(n_12624),
.B(n_12374),
.Y(n_12878)
);

INVx2_ASAP7_75t_L g12879 ( 
.A(n_12518),
.Y(n_12879)
);

AND2x2_ASAP7_75t_L g12880 ( 
.A(n_12691),
.B(n_12411),
.Y(n_12880)
);

AND2x2_ASAP7_75t_L g12881 ( 
.A(n_12679),
.B(n_12405),
.Y(n_12881)
);

NAND2xp5_ASAP7_75t_L g12882 ( 
.A(n_12768),
.B(n_12397),
.Y(n_12882)
);

AND2x2_ASAP7_75t_L g12883 ( 
.A(n_12720),
.B(n_12406),
.Y(n_12883)
);

NAND2x1p5_ASAP7_75t_L g12884 ( 
.A(n_12547),
.B(n_12414),
.Y(n_12884)
);

INVx1_ASAP7_75t_L g12885 ( 
.A(n_12617),
.Y(n_12885)
);

INVx3_ASAP7_75t_L g12886 ( 
.A(n_12696),
.Y(n_12886)
);

AOI21xp33_ASAP7_75t_L g12887 ( 
.A1(n_12719),
.A2(n_12270),
.B(n_12263),
.Y(n_12887)
);

INVx1_ASAP7_75t_L g12888 ( 
.A(n_12621),
.Y(n_12888)
);

AND2x2_ASAP7_75t_L g12889 ( 
.A(n_12724),
.B(n_12398),
.Y(n_12889)
);

INVx2_ASAP7_75t_L g12890 ( 
.A(n_12575),
.Y(n_12890)
);

NAND2xp5_ASAP7_75t_L g12891 ( 
.A(n_12743),
.B(n_12741),
.Y(n_12891)
);

INVx1_ASAP7_75t_L g12892 ( 
.A(n_12625),
.Y(n_12892)
);

INVx2_ASAP7_75t_L g12893 ( 
.A(n_12555),
.Y(n_12893)
);

NAND2xp5_ASAP7_75t_L g12894 ( 
.A(n_12742),
.B(n_12399),
.Y(n_12894)
);

AND2x2_ASAP7_75t_L g12895 ( 
.A(n_12528),
.B(n_12318),
.Y(n_12895)
);

INVx1_ASAP7_75t_L g12896 ( 
.A(n_12635),
.Y(n_12896)
);

AND2x2_ASAP7_75t_L g12897 ( 
.A(n_12723),
.B(n_12335),
.Y(n_12897)
);

AND2x4_ASAP7_75t_L g12898 ( 
.A(n_12562),
.B(n_12305),
.Y(n_12898)
);

INVx8_ASAP7_75t_L g12899 ( 
.A(n_12550),
.Y(n_12899)
);

OR2x2_ASAP7_75t_L g12900 ( 
.A(n_12746),
.B(n_12274),
.Y(n_12900)
);

BUFx2_ASAP7_75t_L g12901 ( 
.A(n_12619),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12637),
.Y(n_12902)
);

AOI21xp5_ASAP7_75t_SL g12903 ( 
.A1(n_12641),
.A2(n_12253),
.B(n_12228),
.Y(n_12903)
);

AOI22xp33_ASAP7_75t_L g12904 ( 
.A1(n_12753),
.A2(n_12271),
.B1(n_12437),
.B2(n_12443),
.Y(n_12904)
);

HB1xp67_ASAP7_75t_L g12905 ( 
.A(n_12726),
.Y(n_12905)
);

BUFx6f_ASAP7_75t_L g12906 ( 
.A(n_12539),
.Y(n_12906)
);

INVx2_ASAP7_75t_L g12907 ( 
.A(n_12567),
.Y(n_12907)
);

NAND2xp5_ASAP7_75t_L g12908 ( 
.A(n_12530),
.B(n_12356),
.Y(n_12908)
);

INVx1_ASAP7_75t_L g12909 ( 
.A(n_12640),
.Y(n_12909)
);

INVx1_ASAP7_75t_L g12910 ( 
.A(n_12642),
.Y(n_12910)
);

HB1xp67_ASAP7_75t_L g12911 ( 
.A(n_12607),
.Y(n_12911)
);

AND2x2_ASAP7_75t_L g12912 ( 
.A(n_12588),
.B(n_12382),
.Y(n_12912)
);

INVx1_ASAP7_75t_L g12913 ( 
.A(n_12643),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_12648),
.Y(n_12914)
);

AND2x4_ASAP7_75t_L g12915 ( 
.A(n_12568),
.B(n_12386),
.Y(n_12915)
);

NAND2xp5_ASAP7_75t_L g12916 ( 
.A(n_12767),
.B(n_12358),
.Y(n_12916)
);

INVxp33_ASAP7_75t_L g12917 ( 
.A(n_12739),
.Y(n_12917)
);

HB1xp67_ASAP7_75t_L g12918 ( 
.A(n_12609),
.Y(n_12918)
);

NAND2xp5_ASAP7_75t_L g12919 ( 
.A(n_12700),
.B(n_1987),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_12656),
.Y(n_12920)
);

NAND2xp5_ASAP7_75t_L g12921 ( 
.A(n_12736),
.B(n_1988),
.Y(n_12921)
);

INVx1_ASAP7_75t_L g12922 ( 
.A(n_12657),
.Y(n_12922)
);

AND2x2_ASAP7_75t_L g12923 ( 
.A(n_12732),
.B(n_1988),
.Y(n_12923)
);

INVx1_ASAP7_75t_SL g12924 ( 
.A(n_12610),
.Y(n_12924)
);

INVx1_ASAP7_75t_L g12925 ( 
.A(n_12659),
.Y(n_12925)
);

INVx2_ASAP7_75t_L g12926 ( 
.A(n_12532),
.Y(n_12926)
);

INVx2_ASAP7_75t_SL g12927 ( 
.A(n_12612),
.Y(n_12927)
);

NAND2xp5_ASAP7_75t_L g12928 ( 
.A(n_12716),
.B(n_1989),
.Y(n_12928)
);

INVx1_ASAP7_75t_L g12929 ( 
.A(n_12664),
.Y(n_12929)
);

INVx1_ASAP7_75t_L g12930 ( 
.A(n_12674),
.Y(n_12930)
);

INVx1_ASAP7_75t_L g12931 ( 
.A(n_12678),
.Y(n_12931)
);

AND2x2_ASAP7_75t_L g12932 ( 
.A(n_12721),
.B(n_12714),
.Y(n_12932)
);

INVx1_ASAP7_75t_L g12933 ( 
.A(n_12688),
.Y(n_12933)
);

INVx2_ASAP7_75t_L g12934 ( 
.A(n_12583),
.Y(n_12934)
);

AND2x4_ASAP7_75t_L g12935 ( 
.A(n_12593),
.B(n_12596),
.Y(n_12935)
);

OAI22xp33_ASAP7_75t_L g12936 ( 
.A1(n_12669),
.A2(n_1991),
.B1(n_1989),
.B2(n_1990),
.Y(n_12936)
);

NAND2xp5_ASAP7_75t_L g12937 ( 
.A(n_12757),
.B(n_1990),
.Y(n_12937)
);

BUFx2_ASAP7_75t_L g12938 ( 
.A(n_12614),
.Y(n_12938)
);

OR2x2_ASAP7_75t_L g12939 ( 
.A(n_12751),
.B(n_1991),
.Y(n_12939)
);

INVx3_ASAP7_75t_L g12940 ( 
.A(n_12601),
.Y(n_12940)
);

INVx2_ASAP7_75t_L g12941 ( 
.A(n_12616),
.Y(n_12941)
);

INVx2_ASAP7_75t_L g12942 ( 
.A(n_12519),
.Y(n_12942)
);

INVx2_ASAP7_75t_L g12943 ( 
.A(n_12549),
.Y(n_12943)
);

AND2x2_ASAP7_75t_L g12944 ( 
.A(n_12712),
.B(n_1993),
.Y(n_12944)
);

INVx2_ASAP7_75t_L g12945 ( 
.A(n_12676),
.Y(n_12945)
);

INVx2_ASAP7_75t_L g12946 ( 
.A(n_12623),
.Y(n_12946)
);

AND2x2_ASAP7_75t_L g12947 ( 
.A(n_12713),
.B(n_1993),
.Y(n_12947)
);

OA21x2_ASAP7_75t_L g12948 ( 
.A1(n_12689),
.A2(n_1994),
.B(n_1995),
.Y(n_12948)
);

INVx3_ASAP7_75t_L g12949 ( 
.A(n_12604),
.Y(n_12949)
);

BUFx6f_ASAP7_75t_SL g12950 ( 
.A(n_12711),
.Y(n_12950)
);

HB1xp67_ASAP7_75t_L g12951 ( 
.A(n_12587),
.Y(n_12951)
);

AND2x2_ASAP7_75t_L g12952 ( 
.A(n_12729),
.B(n_12727),
.Y(n_12952)
);

NAND2xp5_ASAP7_75t_L g12953 ( 
.A(n_12758),
.B(n_12701),
.Y(n_12953)
);

INVx2_ASAP7_75t_L g12954 ( 
.A(n_12638),
.Y(n_12954)
);

INVx2_ASAP7_75t_L g12955 ( 
.A(n_12646),
.Y(n_12955)
);

OR2x2_ASAP7_75t_L g12956 ( 
.A(n_12683),
.B(n_1994),
.Y(n_12956)
);

AND2x2_ASAP7_75t_L g12957 ( 
.A(n_12673),
.B(n_1995),
.Y(n_12957)
);

INVx1_ASAP7_75t_L g12958 ( 
.A(n_12697),
.Y(n_12958)
);

INVx1_ASAP7_75t_L g12959 ( 
.A(n_12704),
.Y(n_12959)
);

AND2x4_ASAP7_75t_L g12960 ( 
.A(n_12654),
.B(n_1996),
.Y(n_12960)
);

INVx1_ASAP7_75t_L g12961 ( 
.A(n_12647),
.Y(n_12961)
);

INVx3_ASAP7_75t_L g12962 ( 
.A(n_12677),
.Y(n_12962)
);

AND2x4_ASAP7_75t_L g12963 ( 
.A(n_12629),
.B(n_1996),
.Y(n_12963)
);

NOR2xp33_ASAP7_75t_L g12964 ( 
.A(n_12599),
.B(n_1997),
.Y(n_12964)
);

AND2x2_ASAP7_75t_L g12965 ( 
.A(n_12653),
.B(n_1997),
.Y(n_12965)
);

AND2x2_ASAP7_75t_L g12966 ( 
.A(n_12668),
.B(n_1998),
.Y(n_12966)
);

INVx1_ASAP7_75t_L g12967 ( 
.A(n_12535),
.Y(n_12967)
);

AND2x2_ASAP7_75t_L g12968 ( 
.A(n_12670),
.B(n_1999),
.Y(n_12968)
);

INVx1_ASAP7_75t_L g12969 ( 
.A(n_12681),
.Y(n_12969)
);

AND2x2_ASAP7_75t_L g12970 ( 
.A(n_12652),
.B(n_1999),
.Y(n_12970)
);

BUFx2_ASAP7_75t_L g12971 ( 
.A(n_12901),
.Y(n_12971)
);

INVx2_ASAP7_75t_L g12972 ( 
.A(n_12775),
.Y(n_12972)
);

AND2x2_ASAP7_75t_L g12973 ( 
.A(n_12837),
.B(n_12699),
.Y(n_12973)
);

INVx1_ASAP7_75t_SL g12974 ( 
.A(n_12872),
.Y(n_12974)
);

INVx1_ASAP7_75t_L g12975 ( 
.A(n_12811),
.Y(n_12975)
);

HB1xp67_ASAP7_75t_L g12976 ( 
.A(n_12860),
.Y(n_12976)
);

INVx1_ASAP7_75t_L g12977 ( 
.A(n_12783),
.Y(n_12977)
);

INVx2_ASAP7_75t_L g12978 ( 
.A(n_12775),
.Y(n_12978)
);

AND2x2_ASAP7_75t_L g12979 ( 
.A(n_12782),
.B(n_12842),
.Y(n_12979)
);

NAND2xp5_ASAP7_75t_L g12980 ( 
.A(n_12845),
.B(n_12762),
.Y(n_12980)
);

INVx1_ASAP7_75t_L g12981 ( 
.A(n_12830),
.Y(n_12981)
);

AND2x2_ASAP7_75t_L g12982 ( 
.A(n_12776),
.B(n_12633),
.Y(n_12982)
);

INVx1_ASAP7_75t_L g12983 ( 
.A(n_12859),
.Y(n_12983)
);

NOR2xp33_ASAP7_75t_L g12984 ( 
.A(n_12808),
.B(n_12725),
.Y(n_12984)
);

OAI22xp5_ASAP7_75t_L g12985 ( 
.A1(n_12795),
.A2(n_12774),
.B1(n_12832),
.B2(n_12814),
.Y(n_12985)
);

INVx2_ASAP7_75t_L g12986 ( 
.A(n_12875),
.Y(n_12986)
);

BUFx3_ASAP7_75t_L g12987 ( 
.A(n_12899),
.Y(n_12987)
);

AND2x2_ASAP7_75t_L g12988 ( 
.A(n_12778),
.B(n_12685),
.Y(n_12988)
);

AND2x2_ASAP7_75t_L g12989 ( 
.A(n_12938),
.B(n_12692),
.Y(n_12989)
);

INVx1_ASAP7_75t_L g12990 ( 
.A(n_12807),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_12824),
.Y(n_12991)
);

INVx2_ASAP7_75t_L g12992 ( 
.A(n_12875),
.Y(n_12992)
);

NAND2xp5_ASAP7_75t_L g12993 ( 
.A(n_12845),
.B(n_12735),
.Y(n_12993)
);

AND2x2_ASAP7_75t_L g12994 ( 
.A(n_12886),
.B(n_12786),
.Y(n_12994)
);

BUFx2_ASAP7_75t_L g12995 ( 
.A(n_12911),
.Y(n_12995)
);

AND2x2_ASAP7_75t_L g12996 ( 
.A(n_12779),
.B(n_12680),
.Y(n_12996)
);

INVx2_ASAP7_75t_L g12997 ( 
.A(n_12828),
.Y(n_12997)
);

NOR2x1_ASAP7_75t_L g12998 ( 
.A(n_12948),
.B(n_12765),
.Y(n_12998)
);

INVx1_ASAP7_75t_L g12999 ( 
.A(n_12905),
.Y(n_12999)
);

BUFx2_ASAP7_75t_L g13000 ( 
.A(n_12918),
.Y(n_13000)
);

INVx2_ASAP7_75t_L g13001 ( 
.A(n_12899),
.Y(n_13001)
);

INVx1_ASAP7_75t_L g13002 ( 
.A(n_12773),
.Y(n_13002)
);

INVx1_ASAP7_75t_L g13003 ( 
.A(n_12781),
.Y(n_13003)
);

AND2x2_ASAP7_75t_L g13004 ( 
.A(n_12789),
.B(n_12690),
.Y(n_13004)
);

BUFx6f_ASAP7_75t_L g13005 ( 
.A(n_12843),
.Y(n_13005)
);

INVx1_ASAP7_75t_L g13006 ( 
.A(n_12844),
.Y(n_13006)
);

HB1xp67_ASAP7_75t_L g13007 ( 
.A(n_12950),
.Y(n_13007)
);

AND2x2_ASAP7_75t_L g13008 ( 
.A(n_12797),
.B(n_12728),
.Y(n_13008)
);

OR2x2_ASAP7_75t_L g13009 ( 
.A(n_12839),
.B(n_12924),
.Y(n_13009)
);

AND2x4_ASAP7_75t_L g13010 ( 
.A(n_12777),
.B(n_12684),
.Y(n_13010)
);

AND2x2_ASAP7_75t_L g13011 ( 
.A(n_12770),
.B(n_12788),
.Y(n_13011)
);

HB1xp67_ASAP7_75t_L g13012 ( 
.A(n_12927),
.Y(n_13012)
);

AND2x2_ASAP7_75t_L g13013 ( 
.A(n_12790),
.B(n_12733),
.Y(n_13013)
);

INVx1_ASAP7_75t_L g13014 ( 
.A(n_12791),
.Y(n_13014)
);

NAND2xp5_ASAP7_75t_L g13015 ( 
.A(n_12845),
.B(n_12754),
.Y(n_13015)
);

INVx1_ASAP7_75t_L g13016 ( 
.A(n_12800),
.Y(n_13016)
);

INVx2_ASAP7_75t_L g13017 ( 
.A(n_12906),
.Y(n_13017)
);

INVx3_ASAP7_75t_SL g13018 ( 
.A(n_12963),
.Y(n_13018)
);

INVx1_ASAP7_75t_L g13019 ( 
.A(n_12801),
.Y(n_13019)
);

INVx5_ASAP7_75t_SL g13020 ( 
.A(n_12960),
.Y(n_13020)
);

NAND2xp5_ASAP7_75t_L g13021 ( 
.A(n_12787),
.B(n_12763),
.Y(n_13021)
);

INVx2_ASAP7_75t_L g13022 ( 
.A(n_12906),
.Y(n_13022)
);

INVx1_ASAP7_75t_L g13023 ( 
.A(n_12816),
.Y(n_13023)
);

AND2x2_ASAP7_75t_L g13024 ( 
.A(n_12771),
.B(n_12686),
.Y(n_13024)
);

INVx1_ASAP7_75t_L g13025 ( 
.A(n_12951),
.Y(n_13025)
);

INVx1_ASAP7_75t_L g13026 ( 
.A(n_12873),
.Y(n_13026)
);

INVx3_ASAP7_75t_L g13027 ( 
.A(n_12780),
.Y(n_13027)
);

AND2x2_ASAP7_75t_L g13028 ( 
.A(n_12796),
.B(n_12687),
.Y(n_13028)
);

BUFx3_ASAP7_75t_L g13029 ( 
.A(n_12785),
.Y(n_13029)
);

AND2x2_ASAP7_75t_L g13030 ( 
.A(n_12941),
.B(n_12675),
.Y(n_13030)
);

HB1xp67_ASAP7_75t_L g13031 ( 
.A(n_12942),
.Y(n_13031)
);

BUFx3_ASAP7_75t_L g13032 ( 
.A(n_12935),
.Y(n_13032)
);

OR2x2_ASAP7_75t_L g13033 ( 
.A(n_12769),
.B(n_12749),
.Y(n_13033)
);

AND2x2_ASAP7_75t_L g13034 ( 
.A(n_12803),
.B(n_12747),
.Y(n_13034)
);

AND2x4_ASAP7_75t_L g13035 ( 
.A(n_12793),
.B(n_12737),
.Y(n_13035)
);

AND2x2_ASAP7_75t_L g13036 ( 
.A(n_12815),
.B(n_12703),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12818),
.Y(n_13037)
);

AND2x2_ASAP7_75t_L g13038 ( 
.A(n_12772),
.B(n_12752),
.Y(n_13038)
);

INVx1_ASAP7_75t_L g13039 ( 
.A(n_12961),
.Y(n_13039)
);

INVx2_ASAP7_75t_L g13040 ( 
.A(n_12838),
.Y(n_13040)
);

INVx1_ASAP7_75t_L g13041 ( 
.A(n_12944),
.Y(n_13041)
);

INVx1_ASAP7_75t_L g13042 ( 
.A(n_12947),
.Y(n_13042)
);

INVx4_ASAP7_75t_L g13043 ( 
.A(n_12848),
.Y(n_13043)
);

AND2x4_ASAP7_75t_SL g13044 ( 
.A(n_12940),
.B(n_12744),
.Y(n_13044)
);

INVx1_ASAP7_75t_L g13045 ( 
.A(n_12923),
.Y(n_13045)
);

AND2x2_ASAP7_75t_L g13046 ( 
.A(n_12865),
.B(n_12750),
.Y(n_13046)
);

OR2x2_ASAP7_75t_SL g13047 ( 
.A(n_12805),
.B(n_12756),
.Y(n_13047)
);

INVx1_ASAP7_75t_L g13048 ( 
.A(n_12821),
.Y(n_13048)
);

INVx1_ASAP7_75t_SL g13049 ( 
.A(n_12794),
.Y(n_13049)
);

OR2x2_ASAP7_75t_L g13050 ( 
.A(n_12804),
.B(n_12564),
.Y(n_13050)
);

AOI22xp5_ASAP7_75t_L g13051 ( 
.A1(n_12806),
.A2(n_12545),
.B1(n_12707),
.B2(n_12644),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12956),
.Y(n_13052)
);

AND2x2_ASAP7_75t_L g13053 ( 
.A(n_12820),
.B(n_12658),
.Y(n_13053)
);

AND2x2_ASAP7_75t_L g13054 ( 
.A(n_12813),
.B(n_12709),
.Y(n_13054)
);

INVx2_ASAP7_75t_SL g13055 ( 
.A(n_12962),
.Y(n_13055)
);

INVx1_ASAP7_75t_L g13056 ( 
.A(n_12893),
.Y(n_13056)
);

INVx2_ASAP7_75t_L g13057 ( 
.A(n_12831),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12907),
.Y(n_13058)
);

INVx2_ASAP7_75t_L g13059 ( 
.A(n_12827),
.Y(n_13059)
);

AND2x2_ASAP7_75t_L g13060 ( 
.A(n_12784),
.B(n_12745),
.Y(n_13060)
);

AND2x2_ASAP7_75t_L g13061 ( 
.A(n_12879),
.B(n_12591),
.Y(n_13061)
);

INVx1_ASAP7_75t_L g13062 ( 
.A(n_12802),
.Y(n_13062)
);

NOR2xp33_ASAP7_75t_L g13063 ( 
.A(n_12917),
.B(n_12620),
.Y(n_13063)
);

INVx2_ASAP7_75t_L g13064 ( 
.A(n_12946),
.Y(n_13064)
);

AND2x2_ASAP7_75t_L g13065 ( 
.A(n_12792),
.B(n_12695),
.Y(n_13065)
);

AOI21xp5_ASAP7_75t_SL g13066 ( 
.A1(n_12819),
.A2(n_12650),
.B(n_12639),
.Y(n_13066)
);

OR2x2_ASAP7_75t_L g13067 ( 
.A(n_12810),
.B(n_12748),
.Y(n_13067)
);

OR2x2_ASAP7_75t_L g13068 ( 
.A(n_12866),
.B(n_12570),
.Y(n_13068)
);

HB1xp67_ASAP7_75t_L g13069 ( 
.A(n_12798),
.Y(n_13069)
);

INVx1_ASAP7_75t_L g13070 ( 
.A(n_12809),
.Y(n_13070)
);

HB1xp67_ASAP7_75t_L g13071 ( 
.A(n_12949),
.Y(n_13071)
);

INVx2_ASAP7_75t_L g13072 ( 
.A(n_12817),
.Y(n_13072)
);

AO21x2_ASAP7_75t_L g13073 ( 
.A1(n_12836),
.A2(n_12671),
.B(n_12755),
.Y(n_13073)
);

INVx1_ASAP7_75t_L g13074 ( 
.A(n_12812),
.Y(n_13074)
);

AND2x2_ASAP7_75t_L g13075 ( 
.A(n_12870),
.B(n_12945),
.Y(n_13075)
);

INVxp67_ASAP7_75t_L g13076 ( 
.A(n_12856),
.Y(n_13076)
);

AND2x2_ASAP7_75t_L g13077 ( 
.A(n_12799),
.B(n_12632),
.Y(n_13077)
);

BUFx2_ASAP7_75t_L g13078 ( 
.A(n_12943),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12954),
.Y(n_13079)
);

INVxp67_ASAP7_75t_L g13080 ( 
.A(n_12867),
.Y(n_13080)
);

OR2x2_ASAP7_75t_L g13081 ( 
.A(n_12953),
.B(n_12926),
.Y(n_13081)
);

INVxp67_ASAP7_75t_SL g13082 ( 
.A(n_12884),
.Y(n_13082)
);

NAND2xp5_ASAP7_75t_L g13083 ( 
.A(n_12829),
.B(n_12895),
.Y(n_13083)
);

HB1xp67_ASAP7_75t_L g13084 ( 
.A(n_12934),
.Y(n_13084)
);

AND2x2_ASAP7_75t_L g13085 ( 
.A(n_12853),
.B(n_12573),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12955),
.Y(n_13086)
);

AND2x2_ASAP7_75t_L g13087 ( 
.A(n_12852),
.B(n_12585),
.Y(n_13087)
);

INVx2_ASAP7_75t_L g13088 ( 
.A(n_12850),
.Y(n_13088)
);

INVxp67_ASAP7_75t_SL g13089 ( 
.A(n_12891),
.Y(n_13089)
);

INVx2_ASAP7_75t_L g13090 ( 
.A(n_12854),
.Y(n_13090)
);

INVx2_ASAP7_75t_SL g13091 ( 
.A(n_12965),
.Y(n_13091)
);

INVx2_ASAP7_75t_L g13092 ( 
.A(n_12855),
.Y(n_13092)
);

AND2x2_ASAP7_75t_L g13093 ( 
.A(n_12858),
.B(n_12833),
.Y(n_13093)
);

NAND2xp5_ASAP7_75t_L g13094 ( 
.A(n_12912),
.B(n_12708),
.Y(n_13094)
);

NAND2xp5_ASAP7_75t_L g13095 ( 
.A(n_12898),
.B(n_12662),
.Y(n_13095)
);

AO21x2_ASAP7_75t_L g13096 ( 
.A1(n_12857),
.A2(n_2000),
.B(n_2001),
.Y(n_13096)
);

BUFx2_ASAP7_75t_L g13097 ( 
.A(n_12890),
.Y(n_13097)
);

INVx2_ASAP7_75t_L g13098 ( 
.A(n_12966),
.Y(n_13098)
);

AO22x1_ASAP7_75t_L g13099 ( 
.A1(n_12851),
.A2(n_2004),
.B1(n_2002),
.B2(n_2003),
.Y(n_13099)
);

INVx1_ASAP7_75t_L g13100 ( 
.A(n_12932),
.Y(n_13100)
);

OR2x2_ASAP7_75t_L g13101 ( 
.A(n_12861),
.B(n_2002),
.Y(n_13101)
);

INVx2_ASAP7_75t_L g13102 ( 
.A(n_12968),
.Y(n_13102)
);

INVx2_ASAP7_75t_L g13103 ( 
.A(n_12970),
.Y(n_13103)
);

AND2x2_ASAP7_75t_L g13104 ( 
.A(n_12835),
.B(n_12863),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12952),
.Y(n_13105)
);

OR2x2_ASAP7_75t_L g13106 ( 
.A(n_12877),
.B(n_12900),
.Y(n_13106)
);

OR2x2_ASAP7_75t_L g13107 ( 
.A(n_12874),
.B(n_2005),
.Y(n_13107)
);

AND2x4_ASAP7_75t_L g13108 ( 
.A(n_12915),
.B(n_2005),
.Y(n_13108)
);

NAND2xp5_ASAP7_75t_L g13109 ( 
.A(n_12869),
.B(n_2006),
.Y(n_13109)
);

AND2x2_ASAP7_75t_L g13110 ( 
.A(n_12880),
.B(n_2006),
.Y(n_13110)
);

INVx1_ASAP7_75t_L g13111 ( 
.A(n_12939),
.Y(n_13111)
);

OR2x2_ASAP7_75t_L g13112 ( 
.A(n_12894),
.B(n_2007),
.Y(n_13112)
);

AND2x4_ASAP7_75t_L g13113 ( 
.A(n_12840),
.B(n_2007),
.Y(n_13113)
);

AND2x2_ASAP7_75t_L g13114 ( 
.A(n_12897),
.B(n_2008),
.Y(n_13114)
);

AND2x2_ASAP7_75t_L g13115 ( 
.A(n_12881),
.B(n_2008),
.Y(n_13115)
);

AND2x2_ASAP7_75t_L g13116 ( 
.A(n_12878),
.B(n_2009),
.Y(n_13116)
);

INVx1_ASAP7_75t_L g13117 ( 
.A(n_12969),
.Y(n_13117)
);

INVx1_ASAP7_75t_L g13118 ( 
.A(n_12822),
.Y(n_13118)
);

HB1xp67_ASAP7_75t_L g13119 ( 
.A(n_12921),
.Y(n_13119)
);

INVx2_ASAP7_75t_L g13120 ( 
.A(n_12957),
.Y(n_13120)
);

AND2x2_ASAP7_75t_L g13121 ( 
.A(n_12889),
.B(n_2009),
.Y(n_13121)
);

AND2x2_ASAP7_75t_L g13122 ( 
.A(n_12883),
.B(n_2010),
.Y(n_13122)
);

INVx1_ASAP7_75t_L g13123 ( 
.A(n_12967),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_12823),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12825),
.Y(n_13125)
);

AND2x2_ASAP7_75t_L g13126 ( 
.A(n_12979),
.B(n_12908),
.Y(n_13126)
);

INVx1_ASAP7_75t_L g13127 ( 
.A(n_12976),
.Y(n_13127)
);

AOI22xp33_ASAP7_75t_L g13128 ( 
.A1(n_12985),
.A2(n_12882),
.B1(n_12846),
.B2(n_12916),
.Y(n_13128)
);

HB1xp67_ASAP7_75t_L g13129 ( 
.A(n_13069),
.Y(n_13129)
);

AO21x2_ASAP7_75t_L g13130 ( 
.A1(n_12980),
.A2(n_13096),
.B(n_13015),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_12995),
.Y(n_13131)
);

OR2x6_ASAP7_75t_L g13132 ( 
.A(n_12971),
.B(n_12972),
.Y(n_13132)
);

AOI22xp33_ASAP7_75t_L g13133 ( 
.A1(n_13073),
.A2(n_12887),
.B1(n_12862),
.B2(n_12904),
.Y(n_13133)
);

INVx1_ASAP7_75t_L g13134 ( 
.A(n_13000),
.Y(n_13134)
);

OAI21x1_ASAP7_75t_L g13135 ( 
.A1(n_13026),
.A2(n_12998),
.B(n_12983),
.Y(n_13135)
);

AOI221xp5_ASAP7_75t_L g13136 ( 
.A1(n_13066),
.A2(n_12903),
.B1(n_12936),
.B2(n_12841),
.C(n_12847),
.Y(n_13136)
);

OAI221xp5_ASAP7_75t_L g13137 ( 
.A1(n_13051),
.A2(n_12849),
.B1(n_12937),
.B2(n_12919),
.C(n_12928),
.Y(n_13137)
);

INVx2_ASAP7_75t_L g13138 ( 
.A(n_12978),
.Y(n_13138)
);

OR2x2_ASAP7_75t_L g13139 ( 
.A(n_13009),
.B(n_12826),
.Y(n_13139)
);

AND2x2_ASAP7_75t_L g13140 ( 
.A(n_12974),
.B(n_12964),
.Y(n_13140)
);

NOR4xp25_ASAP7_75t_SL g13141 ( 
.A(n_13082),
.B(n_12864),
.C(n_12868),
.D(n_12834),
.Y(n_13141)
);

INVx1_ASAP7_75t_SL g13142 ( 
.A(n_13018),
.Y(n_13142)
);

OR2x6_ASAP7_75t_L g13143 ( 
.A(n_13005),
.B(n_12987),
.Y(n_13143)
);

AO21x2_ASAP7_75t_L g13144 ( 
.A1(n_12993),
.A2(n_12876),
.B(n_12871),
.Y(n_13144)
);

AO21x2_ASAP7_75t_L g13145 ( 
.A1(n_13109),
.A2(n_12888),
.B(n_12885),
.Y(n_13145)
);

AOI22xp33_ASAP7_75t_L g13146 ( 
.A1(n_13063),
.A2(n_12896),
.B1(n_12902),
.B2(n_12892),
.Y(n_13146)
);

INVx1_ASAP7_75t_L g13147 ( 
.A(n_13071),
.Y(n_13147)
);

AND2x2_ASAP7_75t_L g13148 ( 
.A(n_12982),
.B(n_12909),
.Y(n_13148)
);

NOR2xp33_ASAP7_75t_R g13149 ( 
.A(n_13005),
.B(n_12910),
.Y(n_13149)
);

OAI221xp5_ASAP7_75t_L g13150 ( 
.A1(n_13076),
.A2(n_12920),
.B1(n_12922),
.B2(n_12914),
.C(n_12913),
.Y(n_13150)
);

OAI211xp5_ASAP7_75t_L g13151 ( 
.A1(n_13094),
.A2(n_13095),
.B(n_13021),
.C(n_13007),
.Y(n_13151)
);

NAND2xp5_ASAP7_75t_L g13152 ( 
.A(n_12989),
.B(n_12925),
.Y(n_13152)
);

BUFx3_ASAP7_75t_L g13153 ( 
.A(n_13032),
.Y(n_13153)
);

AND2x4_ASAP7_75t_L g13154 ( 
.A(n_12994),
.B(n_12929),
.Y(n_13154)
);

HB1xp67_ASAP7_75t_L g13155 ( 
.A(n_13012),
.Y(n_13155)
);

OAI221xp5_ASAP7_75t_L g13156 ( 
.A1(n_13067),
.A2(n_13080),
.B1(n_13068),
.B2(n_13049),
.C(n_13055),
.Y(n_13156)
);

INVx2_ASAP7_75t_L g13157 ( 
.A(n_13020),
.Y(n_13157)
);

OR2x2_ASAP7_75t_L g13158 ( 
.A(n_13033),
.B(n_12930),
.Y(n_13158)
);

AND2x2_ASAP7_75t_L g13159 ( 
.A(n_12973),
.B(n_12931),
.Y(n_13159)
);

OAI221xp5_ASAP7_75t_L g13160 ( 
.A1(n_13106),
.A2(n_12959),
.B1(n_12958),
.B2(n_12933),
.C(n_2013),
.Y(n_13160)
);

OAI22xp5_ASAP7_75t_L g13161 ( 
.A1(n_13047),
.A2(n_13083),
.B1(n_13020),
.B2(n_13050),
.Y(n_13161)
);

INVx2_ASAP7_75t_L g13162 ( 
.A(n_13029),
.Y(n_13162)
);

OAI221xp5_ASAP7_75t_L g13163 ( 
.A1(n_13006),
.A2(n_2013),
.B1(n_2011),
.B2(n_2012),
.C(n_2014),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_12988),
.B(n_2011),
.Y(n_13164)
);

NOR2x2_ASAP7_75t_L g13165 ( 
.A(n_13001),
.B(n_2014),
.Y(n_13165)
);

NAND3xp33_ASAP7_75t_L g13166 ( 
.A(n_12990),
.B(n_12975),
.C(n_13043),
.Y(n_13166)
);

NOR2xp33_ASAP7_75t_R g13167 ( 
.A(n_13027),
.B(n_2015),
.Y(n_13167)
);

OAI22xp5_ASAP7_75t_L g13168 ( 
.A1(n_13089),
.A2(n_12981),
.B1(n_12997),
.B2(n_12992),
.Y(n_13168)
);

NAND4xp25_ASAP7_75t_L g13169 ( 
.A(n_12984),
.B(n_13011),
.C(n_13038),
.D(n_13034),
.Y(n_13169)
);

AOI21xp5_ASAP7_75t_L g13170 ( 
.A1(n_13099),
.A2(n_2015),
.B(n_2016),
.Y(n_13170)
);

OR2x6_ASAP7_75t_L g13171 ( 
.A(n_12986),
.B(n_2016),
.Y(n_13171)
);

AO21x1_ASAP7_75t_SL g13172 ( 
.A1(n_12977),
.A2(n_2017),
.B(n_2018),
.Y(n_13172)
);

OR2x2_ASAP7_75t_L g13173 ( 
.A(n_13101),
.B(n_2017),
.Y(n_13173)
);

INVx1_ASAP7_75t_L g13174 ( 
.A(n_13031),
.Y(n_13174)
);

INVx2_ASAP7_75t_L g13175 ( 
.A(n_13008),
.Y(n_13175)
);

INVx2_ASAP7_75t_L g13176 ( 
.A(n_13004),
.Y(n_13176)
);

INVx2_ASAP7_75t_L g13177 ( 
.A(n_13040),
.Y(n_13177)
);

AOI22xp33_ASAP7_75t_SL g13178 ( 
.A1(n_13085),
.A2(n_2021),
.B1(n_2019),
.B2(n_2020),
.Y(n_13178)
);

INVx2_ASAP7_75t_L g13179 ( 
.A(n_13093),
.Y(n_13179)
);

BUFx3_ASAP7_75t_L g13180 ( 
.A(n_13078),
.Y(n_13180)
);

OR2x2_ASAP7_75t_L g13181 ( 
.A(n_13091),
.B(n_12991),
.Y(n_13181)
);

AND2x2_ASAP7_75t_L g13182 ( 
.A(n_13013),
.B(n_2019),
.Y(n_13182)
);

INVx1_ASAP7_75t_L g13183 ( 
.A(n_13084),
.Y(n_13183)
);

OAI221xp5_ASAP7_75t_L g13184 ( 
.A1(n_13025),
.A2(n_13058),
.B1(n_13056),
.B2(n_13097),
.C(n_13022),
.Y(n_13184)
);

OAI22xp5_ASAP7_75t_L g13185 ( 
.A1(n_13081),
.A2(n_2023),
.B1(n_2020),
.B2(n_2022),
.Y(n_13185)
);

OR2x2_ASAP7_75t_L g13186 ( 
.A(n_12999),
.B(n_2022),
.Y(n_13186)
);

AOI221xp5_ASAP7_75t_L g13187 ( 
.A1(n_13053),
.A2(n_2026),
.B1(n_2024),
.B2(n_2025),
.C(n_2027),
.Y(n_13187)
);

OR2x6_ASAP7_75t_L g13188 ( 
.A(n_13108),
.B(n_2024),
.Y(n_13188)
);

AOI221xp5_ASAP7_75t_L g13189 ( 
.A1(n_13054),
.A2(n_2028),
.B1(n_2026),
.B2(n_2027),
.C(n_2029),
.Y(n_13189)
);

OAI31xp33_ASAP7_75t_L g13190 ( 
.A1(n_13044),
.A2(n_2030),
.A3(n_2028),
.B(n_2029),
.Y(n_13190)
);

INVx1_ASAP7_75t_L g13191 ( 
.A(n_13120),
.Y(n_13191)
);

AND2x2_ASAP7_75t_L g13192 ( 
.A(n_12996),
.B(n_2030),
.Y(n_13192)
);

INVx1_ASAP7_75t_SL g13193 ( 
.A(n_13104),
.Y(n_13193)
);

INVx2_ASAP7_75t_L g13194 ( 
.A(n_13017),
.Y(n_13194)
);

OA21x2_ASAP7_75t_L g13195 ( 
.A1(n_13100),
.A2(n_2031),
.B(n_2032),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_13098),
.Y(n_13196)
);

OAI221xp5_ASAP7_75t_L g13197 ( 
.A1(n_13079),
.A2(n_2033),
.B1(n_2031),
.B2(n_2032),
.C(n_2034),
.Y(n_13197)
);

OAI22xp5_ASAP7_75t_L g13198 ( 
.A1(n_13112),
.A2(n_2036),
.B1(n_2034),
.B2(n_2035),
.Y(n_13198)
);

AOI221xp5_ASAP7_75t_L g13199 ( 
.A1(n_13002),
.A2(n_2037),
.B1(n_2035),
.B2(n_2036),
.C(n_2038),
.Y(n_13199)
);

NAND2xp5_ASAP7_75t_L g13200 ( 
.A(n_13060),
.B(n_13113),
.Y(n_13200)
);

INVx1_ASAP7_75t_L g13201 ( 
.A(n_13102),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_13103),
.Y(n_13202)
);

HB1xp67_ASAP7_75t_L g13203 ( 
.A(n_13114),
.Y(n_13203)
);

NOR2xp33_ASAP7_75t_R g13204 ( 
.A(n_13111),
.B(n_2037),
.Y(n_13204)
);

AND2x2_ASAP7_75t_L g13205 ( 
.A(n_13075),
.B(n_13116),
.Y(n_13205)
);

BUFx2_ASAP7_75t_L g13206 ( 
.A(n_13010),
.Y(n_13206)
);

AOI22xp5_ASAP7_75t_L g13207 ( 
.A1(n_13065),
.A2(n_2040),
.B1(n_2038),
.B2(n_2039),
.Y(n_13207)
);

NOR2xp33_ASAP7_75t_L g13208 ( 
.A(n_13041),
.B(n_2039),
.Y(n_13208)
);

AOI22xp33_ASAP7_75t_L g13209 ( 
.A1(n_13035),
.A2(n_2044),
.B1(n_2040),
.B2(n_2042),
.Y(n_13209)
);

AND2x4_ASAP7_75t_L g13210 ( 
.A(n_13036),
.B(n_2042),
.Y(n_13210)
);

OAI21x1_ASAP7_75t_L g13211 ( 
.A1(n_13024),
.A2(n_2045),
.B(n_2046),
.Y(n_13211)
);

OAI33xp33_ASAP7_75t_L g13212 ( 
.A1(n_13023),
.A2(n_2047),
.A3(n_2049),
.B1(n_2045),
.B2(n_2046),
.B3(n_2048),
.Y(n_13212)
);

NAND3xp33_ASAP7_75t_L g13213 ( 
.A(n_13003),
.B(n_2047),
.C(n_2049),
.Y(n_13213)
);

NAND2xp5_ASAP7_75t_L g13214 ( 
.A(n_13115),
.B(n_2050),
.Y(n_13214)
);

INVx1_ASAP7_75t_L g13215 ( 
.A(n_13042),
.Y(n_13215)
);

OAI31xp33_ASAP7_75t_L g13216 ( 
.A1(n_13077),
.A2(n_2053),
.A3(n_2050),
.B(n_2052),
.Y(n_13216)
);

INVx2_ASAP7_75t_L g13217 ( 
.A(n_13057),
.Y(n_13217)
);

AOI21x1_ASAP7_75t_L g13218 ( 
.A1(n_13110),
.A2(n_2052),
.B(n_2053),
.Y(n_13218)
);

HB1xp67_ASAP7_75t_L g13219 ( 
.A(n_13105),
.Y(n_13219)
);

OAI31xp33_ASAP7_75t_L g13220 ( 
.A1(n_13087),
.A2(n_2056),
.A3(n_2054),
.B(n_2055),
.Y(n_13220)
);

NAND2xp5_ASAP7_75t_L g13221 ( 
.A(n_13046),
.B(n_2056),
.Y(n_13221)
);

AOI22xp33_ASAP7_75t_L g13222 ( 
.A1(n_13028),
.A2(n_2059),
.B1(n_2057),
.B2(n_2058),
.Y(n_13222)
);

NAND2xp33_ASAP7_75t_R g13223 ( 
.A(n_13122),
.B(n_2057),
.Y(n_13223)
);

INVx1_ASAP7_75t_L g13224 ( 
.A(n_13045),
.Y(n_13224)
);

AND2x2_ASAP7_75t_L g13225 ( 
.A(n_13121),
.B(n_2058),
.Y(n_13225)
);

INVx1_ASAP7_75t_L g13226 ( 
.A(n_13030),
.Y(n_13226)
);

OAI33xp33_ASAP7_75t_L g13227 ( 
.A1(n_13014),
.A2(n_2062),
.A3(n_2064),
.B1(n_2059),
.B2(n_2061),
.B3(n_2063),
.Y(n_13227)
);

INVx1_ASAP7_75t_L g13228 ( 
.A(n_13052),
.Y(n_13228)
);

OR2x6_ASAP7_75t_L g13229 ( 
.A(n_13072),
.B(n_2061),
.Y(n_13229)
);

HB1xp67_ASAP7_75t_L g13230 ( 
.A(n_13064),
.Y(n_13230)
);

OAI221xp5_ASAP7_75t_L g13231 ( 
.A1(n_13086),
.A2(n_2064),
.B1(n_2062),
.B2(n_2063),
.C(n_2065),
.Y(n_13231)
);

AND2x2_ASAP7_75t_L g13232 ( 
.A(n_13061),
.B(n_2065),
.Y(n_13232)
);

AO21x1_ASAP7_75t_SL g13233 ( 
.A1(n_13016),
.A2(n_2066),
.B(n_2067),
.Y(n_13233)
);

AND2x2_ASAP7_75t_L g13234 ( 
.A(n_13059),
.B(n_2066),
.Y(n_13234)
);

AND2x4_ASAP7_75t_L g13235 ( 
.A(n_13088),
.B(n_2067),
.Y(n_13235)
);

AND2x4_ASAP7_75t_L g13236 ( 
.A(n_13090),
.B(n_13092),
.Y(n_13236)
);

INVx2_ASAP7_75t_L g13237 ( 
.A(n_13019),
.Y(n_13237)
);

INVx1_ASAP7_75t_L g13238 ( 
.A(n_13048),
.Y(n_13238)
);

AO21x2_ASAP7_75t_L g13239 ( 
.A1(n_13107),
.A2(n_2068),
.B(n_2069),
.Y(n_13239)
);

INVx2_ASAP7_75t_L g13240 ( 
.A(n_13037),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_13039),
.Y(n_13241)
);

NAND2xp5_ASAP7_75t_SL g13242 ( 
.A(n_13119),
.B(n_2068),
.Y(n_13242)
);

INVx1_ASAP7_75t_L g13243 ( 
.A(n_13062),
.Y(n_13243)
);

INVx1_ASAP7_75t_L g13244 ( 
.A(n_13070),
.Y(n_13244)
);

AOI221xp5_ASAP7_75t_L g13245 ( 
.A1(n_13074),
.A2(n_2071),
.B1(n_2069),
.B2(n_2070),
.C(n_2072),
.Y(n_13245)
);

OAI222xp33_ASAP7_75t_L g13246 ( 
.A1(n_13117),
.A2(n_2073),
.B1(n_2075),
.B2(n_2070),
.C1(n_2072),
.C2(n_2074),
.Y(n_13246)
);

OR2x2_ASAP7_75t_L g13247 ( 
.A(n_13118),
.B(n_2073),
.Y(n_13247)
);

OAI22xp5_ASAP7_75t_L g13248 ( 
.A1(n_13123),
.A2(n_2076),
.B1(n_2074),
.B2(n_2075),
.Y(n_13248)
);

INVx2_ASAP7_75t_L g13249 ( 
.A(n_13124),
.Y(n_13249)
);

INVx1_ASAP7_75t_L g13250 ( 
.A(n_13125),
.Y(n_13250)
);

NAND2xp5_ASAP7_75t_L g13251 ( 
.A(n_12974),
.B(n_2076),
.Y(n_13251)
);

INVx1_ASAP7_75t_SL g13252 ( 
.A(n_12974),
.Y(n_13252)
);

OR2x6_ASAP7_75t_L g13253 ( 
.A(n_12971),
.B(n_2077),
.Y(n_13253)
);

NOR2xp33_ASAP7_75t_L g13254 ( 
.A(n_12974),
.B(n_2077),
.Y(n_13254)
);

AND2x2_ASAP7_75t_L g13255 ( 
.A(n_12979),
.B(n_2078),
.Y(n_13255)
);

AND2x2_ASAP7_75t_L g13256 ( 
.A(n_12979),
.B(n_2078),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_12976),
.Y(n_13257)
);

BUFx2_ASAP7_75t_L g13258 ( 
.A(n_13132),
.Y(n_13258)
);

INVx1_ASAP7_75t_L g13259 ( 
.A(n_13129),
.Y(n_13259)
);

OR2x2_ASAP7_75t_L g13260 ( 
.A(n_13193),
.B(n_2079),
.Y(n_13260)
);

AND2x2_ASAP7_75t_L g13261 ( 
.A(n_13142),
.B(n_13252),
.Y(n_13261)
);

INVx2_ASAP7_75t_L g13262 ( 
.A(n_13132),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_13157),
.B(n_2079),
.Y(n_13263)
);

AND2x2_ASAP7_75t_L g13264 ( 
.A(n_13143),
.B(n_2080),
.Y(n_13264)
);

INVx2_ASAP7_75t_L g13265 ( 
.A(n_13165),
.Y(n_13265)
);

HB1xp67_ASAP7_75t_L g13266 ( 
.A(n_13155),
.Y(n_13266)
);

AND2x2_ASAP7_75t_L g13267 ( 
.A(n_13143),
.B(n_2080),
.Y(n_13267)
);

AOI22xp33_ASAP7_75t_L g13268 ( 
.A1(n_13136),
.A2(n_13133),
.B1(n_13153),
.B2(n_13128),
.Y(n_13268)
);

INVx3_ASAP7_75t_L g13269 ( 
.A(n_13180),
.Y(n_13269)
);

HB1xp67_ASAP7_75t_L g13270 ( 
.A(n_13253),
.Y(n_13270)
);

NAND2xp5_ASAP7_75t_L g13271 ( 
.A(n_13205),
.B(n_2081),
.Y(n_13271)
);

INVx1_ASAP7_75t_L g13272 ( 
.A(n_13203),
.Y(n_13272)
);

AND2x2_ASAP7_75t_L g13273 ( 
.A(n_13162),
.B(n_2081),
.Y(n_13273)
);

NAND2xp5_ASAP7_75t_L g13274 ( 
.A(n_13206),
.B(n_2082),
.Y(n_13274)
);

AND2x2_ASAP7_75t_L g13275 ( 
.A(n_13126),
.B(n_2082),
.Y(n_13275)
);

INVx1_ASAP7_75t_L g13276 ( 
.A(n_13253),
.Y(n_13276)
);

INVx1_ASAP7_75t_L g13277 ( 
.A(n_13182),
.Y(n_13277)
);

NAND2xp5_ASAP7_75t_L g13278 ( 
.A(n_13127),
.B(n_2083),
.Y(n_13278)
);

AND2x2_ASAP7_75t_L g13279 ( 
.A(n_13140),
.B(n_2083),
.Y(n_13279)
);

OR2x2_ASAP7_75t_L g13280 ( 
.A(n_13169),
.B(n_2084),
.Y(n_13280)
);

NAND2xp5_ASAP7_75t_L g13281 ( 
.A(n_13257),
.B(n_2084),
.Y(n_13281)
);

INVx1_ASAP7_75t_L g13282 ( 
.A(n_13192),
.Y(n_13282)
);

AND2x4_ASAP7_75t_SL g13283 ( 
.A(n_13154),
.B(n_2085),
.Y(n_13283)
);

INVx1_ASAP7_75t_L g13284 ( 
.A(n_13131),
.Y(n_13284)
);

AND2x2_ASAP7_75t_L g13285 ( 
.A(n_13175),
.B(n_13148),
.Y(n_13285)
);

NAND2xp5_ASAP7_75t_L g13286 ( 
.A(n_13134),
.B(n_2086),
.Y(n_13286)
);

AND2x2_ASAP7_75t_L g13287 ( 
.A(n_13179),
.B(n_2087),
.Y(n_13287)
);

INVx1_ASAP7_75t_L g13288 ( 
.A(n_13251),
.Y(n_13288)
);

NAND4xp25_ASAP7_75t_L g13289 ( 
.A(n_13156),
.B(n_2090),
.C(n_2088),
.D(n_2089),
.Y(n_13289)
);

NAND2xp5_ASAP7_75t_SL g13290 ( 
.A(n_13170),
.B(n_2088),
.Y(n_13290)
);

HB1xp67_ASAP7_75t_L g13291 ( 
.A(n_13167),
.Y(n_13291)
);

AND2x2_ASAP7_75t_L g13292 ( 
.A(n_13176),
.B(n_2089),
.Y(n_13292)
);

AND2x2_ASAP7_75t_L g13293 ( 
.A(n_13138),
.B(n_2090),
.Y(n_13293)
);

NAND2xp5_ASAP7_75t_L g13294 ( 
.A(n_13147),
.B(n_2092),
.Y(n_13294)
);

AND2x4_ASAP7_75t_L g13295 ( 
.A(n_13166),
.B(n_2092),
.Y(n_13295)
);

INVx2_ASAP7_75t_L g13296 ( 
.A(n_13171),
.Y(n_13296)
);

INVx1_ASAP7_75t_L g13297 ( 
.A(n_13219),
.Y(n_13297)
);

AND2x2_ASAP7_75t_L g13298 ( 
.A(n_13159),
.B(n_2093),
.Y(n_13298)
);

NAND2xp5_ASAP7_75t_L g13299 ( 
.A(n_13255),
.B(n_2093),
.Y(n_13299)
);

AND2x2_ASAP7_75t_L g13300 ( 
.A(n_13164),
.B(n_2094),
.Y(n_13300)
);

INVx1_ASAP7_75t_L g13301 ( 
.A(n_13181),
.Y(n_13301)
);

AND2x4_ASAP7_75t_L g13302 ( 
.A(n_13256),
.B(n_2094),
.Y(n_13302)
);

INVx2_ASAP7_75t_L g13303 ( 
.A(n_13171),
.Y(n_13303)
);

AND2x2_ASAP7_75t_L g13304 ( 
.A(n_13254),
.B(n_2095),
.Y(n_13304)
);

HB1xp67_ASAP7_75t_L g13305 ( 
.A(n_13229),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_13225),
.Y(n_13306)
);

INVxp67_ASAP7_75t_SL g13307 ( 
.A(n_13223),
.Y(n_13307)
);

INVx2_ASAP7_75t_L g13308 ( 
.A(n_13188),
.Y(n_13308)
);

NAND2xp5_ASAP7_75t_L g13309 ( 
.A(n_13178),
.B(n_2095),
.Y(n_13309)
);

INVx1_ASAP7_75t_L g13310 ( 
.A(n_13230),
.Y(n_13310)
);

BUFx3_ASAP7_75t_L g13311 ( 
.A(n_13210),
.Y(n_13311)
);

INVx1_ASAP7_75t_L g13312 ( 
.A(n_13158),
.Y(n_13312)
);

INVx1_ASAP7_75t_L g13313 ( 
.A(n_13229),
.Y(n_13313)
);

NOR2x1_ASAP7_75t_R g13314 ( 
.A(n_13242),
.B(n_13200),
.Y(n_13314)
);

OR2x2_ASAP7_75t_L g13315 ( 
.A(n_13139),
.B(n_2096),
.Y(n_13315)
);

INVx2_ASAP7_75t_L g13316 ( 
.A(n_13188),
.Y(n_13316)
);

INVx1_ASAP7_75t_L g13317 ( 
.A(n_13152),
.Y(n_13317)
);

INVxp67_ASAP7_75t_L g13318 ( 
.A(n_13172),
.Y(n_13318)
);

AND2x2_ASAP7_75t_L g13319 ( 
.A(n_13177),
.B(n_2096),
.Y(n_13319)
);

INVx4_ASAP7_75t_L g13320 ( 
.A(n_13236),
.Y(n_13320)
);

OR2x2_ASAP7_75t_L g13321 ( 
.A(n_13174),
.B(n_2097),
.Y(n_13321)
);

AND2x4_ASAP7_75t_L g13322 ( 
.A(n_13183),
.B(n_2097),
.Y(n_13322)
);

HB1xp67_ASAP7_75t_L g13323 ( 
.A(n_13204),
.Y(n_13323)
);

NAND2xp5_ASAP7_75t_L g13324 ( 
.A(n_13130),
.B(n_2098),
.Y(n_13324)
);

INVx1_ASAP7_75t_L g13325 ( 
.A(n_13173),
.Y(n_13325)
);

AND2x2_ASAP7_75t_L g13326 ( 
.A(n_13194),
.B(n_2098),
.Y(n_13326)
);

INVx1_ASAP7_75t_L g13327 ( 
.A(n_13232),
.Y(n_13327)
);

INVx1_ASAP7_75t_L g13328 ( 
.A(n_13214),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_13186),
.Y(n_13329)
);

NAND2xp5_ASAP7_75t_L g13330 ( 
.A(n_13190),
.B(n_13161),
.Y(n_13330)
);

AND2x2_ASAP7_75t_L g13331 ( 
.A(n_13226),
.B(n_2099),
.Y(n_13331)
);

NOR2xp33_ASAP7_75t_L g13332 ( 
.A(n_13151),
.B(n_2101),
.Y(n_13332)
);

AND2x2_ASAP7_75t_L g13333 ( 
.A(n_13191),
.B(n_2102),
.Y(n_13333)
);

INVx2_ASAP7_75t_L g13334 ( 
.A(n_13135),
.Y(n_13334)
);

NAND2xp5_ASAP7_75t_L g13335 ( 
.A(n_13239),
.B(n_2104),
.Y(n_13335)
);

NAND2x1p5_ASAP7_75t_L g13336 ( 
.A(n_13211),
.B(n_2104),
.Y(n_13336)
);

AND2x2_ASAP7_75t_L g13337 ( 
.A(n_13196),
.B(n_13201),
.Y(n_13337)
);

INVx1_ASAP7_75t_L g13338 ( 
.A(n_13247),
.Y(n_13338)
);

AND2x2_ASAP7_75t_L g13339 ( 
.A(n_13202),
.B(n_13149),
.Y(n_13339)
);

INVx1_ASAP7_75t_L g13340 ( 
.A(n_13234),
.Y(n_13340)
);

AND2x2_ASAP7_75t_L g13341 ( 
.A(n_13217),
.B(n_2105),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_13215),
.B(n_2105),
.Y(n_13342)
);

AOI21xp5_ASAP7_75t_L g13343 ( 
.A1(n_13141),
.A2(n_2106),
.B(n_2107),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_13224),
.B(n_2106),
.Y(n_13344)
);

AND2x2_ASAP7_75t_L g13345 ( 
.A(n_13228),
.B(n_2107),
.Y(n_13345)
);

NAND2xp5_ASAP7_75t_L g13346 ( 
.A(n_13216),
.B(n_2108),
.Y(n_13346)
);

INVx2_ASAP7_75t_L g13347 ( 
.A(n_13235),
.Y(n_13347)
);

INVx1_ASAP7_75t_L g13348 ( 
.A(n_13218),
.Y(n_13348)
);

AND2x2_ASAP7_75t_L g13349 ( 
.A(n_13195),
.B(n_13168),
.Y(n_13349)
);

AND2x2_ASAP7_75t_L g13350 ( 
.A(n_13146),
.B(n_13145),
.Y(n_13350)
);

AND2x2_ASAP7_75t_L g13351 ( 
.A(n_13221),
.B(n_2109),
.Y(n_13351)
);

NAND2xp5_ASAP7_75t_L g13352 ( 
.A(n_13220),
.B(n_2109),
.Y(n_13352)
);

INVxp67_ASAP7_75t_SL g13353 ( 
.A(n_13208),
.Y(n_13353)
);

AND2x2_ASAP7_75t_L g13354 ( 
.A(n_13237),
.B(n_2111),
.Y(n_13354)
);

CKINVDCx16_ASAP7_75t_R g13355 ( 
.A(n_13144),
.Y(n_13355)
);

AND2x2_ASAP7_75t_L g13356 ( 
.A(n_13233),
.B(n_2112),
.Y(n_13356)
);

AND2x2_ASAP7_75t_L g13357 ( 
.A(n_13240),
.B(n_2112),
.Y(n_13357)
);

INVx2_ASAP7_75t_L g13358 ( 
.A(n_13238),
.Y(n_13358)
);

OR2x2_ASAP7_75t_L g13359 ( 
.A(n_13184),
.B(n_2113),
.Y(n_13359)
);

INVx1_ASAP7_75t_L g13360 ( 
.A(n_13241),
.Y(n_13360)
);

AND2x2_ASAP7_75t_L g13361 ( 
.A(n_13207),
.B(n_13249),
.Y(n_13361)
);

INVx1_ASAP7_75t_L g13362 ( 
.A(n_13243),
.Y(n_13362)
);

INVx1_ASAP7_75t_L g13363 ( 
.A(n_13250),
.Y(n_13363)
);

AND2x2_ASAP7_75t_L g13364 ( 
.A(n_13244),
.B(n_2113),
.Y(n_13364)
);

NOR2xp33_ASAP7_75t_L g13365 ( 
.A(n_13137),
.B(n_13160),
.Y(n_13365)
);

OAI21xp33_ASAP7_75t_L g13366 ( 
.A1(n_13150),
.A2(n_2115),
.B(n_2116),
.Y(n_13366)
);

INVx1_ASAP7_75t_L g13367 ( 
.A(n_13213),
.Y(n_13367)
);

INVx1_ASAP7_75t_L g13368 ( 
.A(n_13248),
.Y(n_13368)
);

OR2x2_ASAP7_75t_L g13369 ( 
.A(n_13198),
.B(n_2115),
.Y(n_13369)
);

AND2x4_ASAP7_75t_L g13370 ( 
.A(n_13209),
.B(n_2117),
.Y(n_13370)
);

INVxp67_ASAP7_75t_L g13371 ( 
.A(n_13163),
.Y(n_13371)
);

INVx1_ASAP7_75t_L g13372 ( 
.A(n_13185),
.Y(n_13372)
);

INVx1_ASAP7_75t_L g13373 ( 
.A(n_13356),
.Y(n_13373)
);

AND2x2_ASAP7_75t_L g13374 ( 
.A(n_13265),
.B(n_13222),
.Y(n_13374)
);

OR2x2_ASAP7_75t_L g13375 ( 
.A(n_13307),
.B(n_13197),
.Y(n_13375)
);

INVx2_ASAP7_75t_L g13376 ( 
.A(n_13258),
.Y(n_13376)
);

OR2x2_ASAP7_75t_L g13377 ( 
.A(n_13318),
.B(n_13231),
.Y(n_13377)
);

INVx1_ASAP7_75t_L g13378 ( 
.A(n_13266),
.Y(n_13378)
);

AND2x4_ASAP7_75t_L g13379 ( 
.A(n_13261),
.B(n_13212),
.Y(n_13379)
);

AND2x2_ASAP7_75t_L g13380 ( 
.A(n_13262),
.B(n_13187),
.Y(n_13380)
);

NAND2xp5_ASAP7_75t_L g13381 ( 
.A(n_13270),
.B(n_13189),
.Y(n_13381)
);

INVx2_ASAP7_75t_L g13382 ( 
.A(n_13320),
.Y(n_13382)
);

AND2x2_ASAP7_75t_L g13383 ( 
.A(n_13285),
.B(n_13199),
.Y(n_13383)
);

INVx1_ASAP7_75t_L g13384 ( 
.A(n_13323),
.Y(n_13384)
);

INVx1_ASAP7_75t_L g13385 ( 
.A(n_13291),
.Y(n_13385)
);

INVx1_ASAP7_75t_L g13386 ( 
.A(n_13305),
.Y(n_13386)
);

NOR2xp33_ASAP7_75t_L g13387 ( 
.A(n_13269),
.B(n_13296),
.Y(n_13387)
);

HB1xp67_ASAP7_75t_L g13388 ( 
.A(n_13355),
.Y(n_13388)
);

NAND2xp5_ASAP7_75t_L g13389 ( 
.A(n_13349),
.B(n_13245),
.Y(n_13389)
);

INVx1_ASAP7_75t_L g13390 ( 
.A(n_13303),
.Y(n_13390)
);

NAND2xp5_ASAP7_75t_SL g13391 ( 
.A(n_13259),
.B(n_13227),
.Y(n_13391)
);

OR2x2_ASAP7_75t_L g13392 ( 
.A(n_13289),
.B(n_13246),
.Y(n_13392)
);

INVx1_ASAP7_75t_L g13393 ( 
.A(n_13279),
.Y(n_13393)
);

INVx2_ASAP7_75t_L g13394 ( 
.A(n_13311),
.Y(n_13394)
);

INVx2_ASAP7_75t_L g13395 ( 
.A(n_13283),
.Y(n_13395)
);

AND2x4_ASAP7_75t_L g13396 ( 
.A(n_13308),
.B(n_2117),
.Y(n_13396)
);

BUFx2_ASAP7_75t_L g13397 ( 
.A(n_13336),
.Y(n_13397)
);

AND2x2_ASAP7_75t_L g13398 ( 
.A(n_13316),
.B(n_2118),
.Y(n_13398)
);

INVx2_ASAP7_75t_L g13399 ( 
.A(n_13264),
.Y(n_13399)
);

OR2x2_ASAP7_75t_L g13400 ( 
.A(n_13276),
.B(n_2118),
.Y(n_13400)
);

INVx1_ASAP7_75t_L g13401 ( 
.A(n_13298),
.Y(n_13401)
);

NAND2xp5_ASAP7_75t_L g13402 ( 
.A(n_13267),
.B(n_13313),
.Y(n_13402)
);

INVx1_ASAP7_75t_L g13403 ( 
.A(n_13275),
.Y(n_13403)
);

AND2x2_ASAP7_75t_L g13404 ( 
.A(n_13339),
.B(n_2119),
.Y(n_13404)
);

OR2x2_ASAP7_75t_L g13405 ( 
.A(n_13260),
.B(n_2120),
.Y(n_13405)
);

OR2x6_ASAP7_75t_L g13406 ( 
.A(n_13301),
.B(n_2120),
.Y(n_13406)
);

AND2x2_ASAP7_75t_L g13407 ( 
.A(n_13263),
.B(n_13327),
.Y(n_13407)
);

INVx1_ASAP7_75t_L g13408 ( 
.A(n_13272),
.Y(n_13408)
);

AND2x4_ASAP7_75t_L g13409 ( 
.A(n_13277),
.B(n_2121),
.Y(n_13409)
);

AND2x2_ASAP7_75t_L g13410 ( 
.A(n_13282),
.B(n_2121),
.Y(n_13410)
);

AND2x4_ASAP7_75t_SL g13411 ( 
.A(n_13347),
.B(n_2122),
.Y(n_13411)
);

AND2x2_ASAP7_75t_L g13412 ( 
.A(n_13306),
.B(n_2122),
.Y(n_13412)
);

NOR4xp25_ASAP7_75t_SL g13413 ( 
.A(n_13348),
.B(n_2125),
.C(n_2123),
.D(n_2124),
.Y(n_13413)
);

AOI22xp33_ASAP7_75t_L g13414 ( 
.A1(n_13350),
.A2(n_2126),
.B1(n_2123),
.B2(n_2125),
.Y(n_13414)
);

OR2x2_ASAP7_75t_L g13415 ( 
.A(n_13359),
.B(n_2126),
.Y(n_13415)
);

AND2x2_ASAP7_75t_L g13416 ( 
.A(n_13361),
.B(n_13312),
.Y(n_13416)
);

NOR2xp33_ASAP7_75t_L g13417 ( 
.A(n_13366),
.B(n_2127),
.Y(n_13417)
);

INVx2_ASAP7_75t_L g13418 ( 
.A(n_13302),
.Y(n_13418)
);

AND2x2_ASAP7_75t_L g13419 ( 
.A(n_13340),
.B(n_2128),
.Y(n_13419)
);

INVx1_ASAP7_75t_L g13420 ( 
.A(n_13274),
.Y(n_13420)
);

INVx1_ASAP7_75t_L g13421 ( 
.A(n_13300),
.Y(n_13421)
);

OA21x2_ASAP7_75t_L g13422 ( 
.A1(n_13343),
.A2(n_2129),
.B(n_2130),
.Y(n_13422)
);

AND2x4_ASAP7_75t_L g13423 ( 
.A(n_13273),
.B(n_2131),
.Y(n_13423)
);

INVx2_ASAP7_75t_L g13424 ( 
.A(n_13315),
.Y(n_13424)
);

AND2x2_ASAP7_75t_L g13425 ( 
.A(n_13353),
.B(n_2132),
.Y(n_13425)
);

AND2x2_ASAP7_75t_L g13426 ( 
.A(n_13372),
.B(n_2133),
.Y(n_13426)
);

AOI21xp33_ASAP7_75t_L g13427 ( 
.A1(n_13314),
.A2(n_2133),
.B(n_2134),
.Y(n_13427)
);

AND2x2_ASAP7_75t_L g13428 ( 
.A(n_13295),
.B(n_2134),
.Y(n_13428)
);

INVx2_ASAP7_75t_L g13429 ( 
.A(n_13293),
.Y(n_13429)
);

INVx1_ASAP7_75t_L g13430 ( 
.A(n_13297),
.Y(n_13430)
);

INVx1_ASAP7_75t_L g13431 ( 
.A(n_13271),
.Y(n_13431)
);

INVx3_ASAP7_75t_L g13432 ( 
.A(n_13322),
.Y(n_13432)
);

INVxp67_ASAP7_75t_SL g13433 ( 
.A(n_13335),
.Y(n_13433)
);

INVx1_ASAP7_75t_L g13434 ( 
.A(n_13292),
.Y(n_13434)
);

AND2x2_ASAP7_75t_L g13435 ( 
.A(n_13368),
.B(n_2135),
.Y(n_13435)
);

OR2x2_ASAP7_75t_L g13436 ( 
.A(n_13280),
.B(n_2136),
.Y(n_13436)
);

INVx3_ASAP7_75t_L g13437 ( 
.A(n_13310),
.Y(n_13437)
);

AND2x2_ASAP7_75t_L g13438 ( 
.A(n_13367),
.B(n_2136),
.Y(n_13438)
);

INVx2_ASAP7_75t_SL g13439 ( 
.A(n_13326),
.Y(n_13439)
);

INVx1_ASAP7_75t_L g13440 ( 
.A(n_13287),
.Y(n_13440)
);

INVx2_ASAP7_75t_L g13441 ( 
.A(n_13321),
.Y(n_13441)
);

AND2x2_ASAP7_75t_L g13442 ( 
.A(n_13284),
.B(n_2137),
.Y(n_13442)
);

AND2x2_ASAP7_75t_SL g13443 ( 
.A(n_13330),
.B(n_2137),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_13337),
.B(n_2138),
.Y(n_13444)
);

AND2x2_ASAP7_75t_L g13445 ( 
.A(n_13325),
.B(n_2138),
.Y(n_13445)
);

INVx1_ASAP7_75t_L g13446 ( 
.A(n_13331),
.Y(n_13446)
);

NOR2xp33_ASAP7_75t_L g13447 ( 
.A(n_13290),
.B(n_2139),
.Y(n_13447)
);

NOR3xp33_ASAP7_75t_SL g13448 ( 
.A(n_13365),
.B(n_2139),
.C(n_2141),
.Y(n_13448)
);

NOR2xp33_ASAP7_75t_L g13449 ( 
.A(n_13371),
.B(n_2142),
.Y(n_13449)
);

INVx1_ASAP7_75t_L g13450 ( 
.A(n_13299),
.Y(n_13450)
);

AND2x2_ASAP7_75t_L g13451 ( 
.A(n_13329),
.B(n_2142),
.Y(n_13451)
);

INVx1_ASAP7_75t_L g13452 ( 
.A(n_13333),
.Y(n_13452)
);

INVx1_ASAP7_75t_L g13453 ( 
.A(n_13304),
.Y(n_13453)
);

HB1xp67_ASAP7_75t_L g13454 ( 
.A(n_13324),
.Y(n_13454)
);

INVxp67_ASAP7_75t_L g13455 ( 
.A(n_13332),
.Y(n_13455)
);

AND2x2_ASAP7_75t_L g13456 ( 
.A(n_13351),
.B(n_2143),
.Y(n_13456)
);

AND2x2_ASAP7_75t_L g13457 ( 
.A(n_13288),
.B(n_2143),
.Y(n_13457)
);

INVx2_ASAP7_75t_L g13458 ( 
.A(n_13342),
.Y(n_13458)
);

NAND2xp5_ASAP7_75t_L g13459 ( 
.A(n_13268),
.B(n_2144),
.Y(n_13459)
);

INVx4_ASAP7_75t_L g13460 ( 
.A(n_13319),
.Y(n_13460)
);

INVx2_ASAP7_75t_L g13461 ( 
.A(n_13344),
.Y(n_13461)
);

NOR2xp33_ASAP7_75t_L g13462 ( 
.A(n_13309),
.B(n_2144),
.Y(n_13462)
);

INVx2_ASAP7_75t_L g13463 ( 
.A(n_13345),
.Y(n_13463)
);

AND2x2_ASAP7_75t_L g13464 ( 
.A(n_13317),
.B(n_2145),
.Y(n_13464)
);

NAND2xp5_ASAP7_75t_L g13465 ( 
.A(n_13370),
.B(n_2146),
.Y(n_13465)
);

AND2x4_ASAP7_75t_SL g13466 ( 
.A(n_13338),
.B(n_2146),
.Y(n_13466)
);

AND2x2_ASAP7_75t_L g13467 ( 
.A(n_13341),
.B(n_2148),
.Y(n_13467)
);

AND2x2_ASAP7_75t_L g13468 ( 
.A(n_13328),
.B(n_2149),
.Y(n_13468)
);

INVx1_ASAP7_75t_L g13469 ( 
.A(n_13364),
.Y(n_13469)
);

AND2x2_ASAP7_75t_L g13470 ( 
.A(n_13354),
.B(n_2150),
.Y(n_13470)
);

NOR2x1_ASAP7_75t_L g13471 ( 
.A(n_13334),
.B(n_2150),
.Y(n_13471)
);

AND2x2_ASAP7_75t_L g13472 ( 
.A(n_13357),
.B(n_2151),
.Y(n_13472)
);

AND2x2_ASAP7_75t_L g13473 ( 
.A(n_13346),
.B(n_2151),
.Y(n_13473)
);

NAND2xp33_ASAP7_75t_R g13474 ( 
.A(n_13369),
.B(n_2152),
.Y(n_13474)
);

AND2x2_ASAP7_75t_L g13475 ( 
.A(n_13352),
.B(n_2153),
.Y(n_13475)
);

BUFx3_ASAP7_75t_L g13476 ( 
.A(n_13286),
.Y(n_13476)
);

AND2x2_ASAP7_75t_L g13477 ( 
.A(n_13358),
.B(n_2153),
.Y(n_13477)
);

AND2x2_ASAP7_75t_L g13478 ( 
.A(n_13360),
.B(n_2154),
.Y(n_13478)
);

AND2x2_ASAP7_75t_L g13479 ( 
.A(n_13362),
.B(n_2154),
.Y(n_13479)
);

INVx2_ASAP7_75t_L g13480 ( 
.A(n_13278),
.Y(n_13480)
);

AND2x2_ASAP7_75t_L g13481 ( 
.A(n_13363),
.B(n_2155),
.Y(n_13481)
);

INVx1_ASAP7_75t_L g13482 ( 
.A(n_13281),
.Y(n_13482)
);

NAND2xp5_ASAP7_75t_L g13483 ( 
.A(n_13294),
.B(n_2155),
.Y(n_13483)
);

INVx1_ASAP7_75t_L g13484 ( 
.A(n_13356),
.Y(n_13484)
);

INVx2_ASAP7_75t_L g13485 ( 
.A(n_13356),
.Y(n_13485)
);

AND2x2_ASAP7_75t_L g13486 ( 
.A(n_13265),
.B(n_2156),
.Y(n_13486)
);

BUFx6f_ASAP7_75t_L g13487 ( 
.A(n_13261),
.Y(n_13487)
);

OA21x2_ASAP7_75t_L g13488 ( 
.A1(n_13343),
.A2(n_2156),
.B(n_2157),
.Y(n_13488)
);

NAND2xp5_ASAP7_75t_L g13489 ( 
.A(n_13265),
.B(n_2158),
.Y(n_13489)
);

AND2x2_ASAP7_75t_L g13490 ( 
.A(n_13265),
.B(n_2159),
.Y(n_13490)
);

AND2x2_ASAP7_75t_L g13491 ( 
.A(n_13265),
.B(n_2159),
.Y(n_13491)
);

INVx2_ASAP7_75t_L g13492 ( 
.A(n_13356),
.Y(n_13492)
);

INVx1_ASAP7_75t_SL g13493 ( 
.A(n_13356),
.Y(n_13493)
);

INVx1_ASAP7_75t_L g13494 ( 
.A(n_13356),
.Y(n_13494)
);

INVx1_ASAP7_75t_SL g13495 ( 
.A(n_13356),
.Y(n_13495)
);

NAND2xp5_ASAP7_75t_L g13496 ( 
.A(n_13265),
.B(n_2160),
.Y(n_13496)
);

NAND2x1p5_ASAP7_75t_L g13497 ( 
.A(n_13261),
.B(n_2160),
.Y(n_13497)
);

AND2x2_ASAP7_75t_L g13498 ( 
.A(n_13485),
.B(n_2161),
.Y(n_13498)
);

NAND2xp5_ASAP7_75t_SL g13499 ( 
.A(n_13487),
.B(n_2161),
.Y(n_13499)
);

NOR2xp33_ASAP7_75t_L g13500 ( 
.A(n_13493),
.B(n_2162),
.Y(n_13500)
);

AND2x2_ASAP7_75t_L g13501 ( 
.A(n_13492),
.B(n_2162),
.Y(n_13501)
);

INVx1_ASAP7_75t_L g13502 ( 
.A(n_13373),
.Y(n_13502)
);

INVxp67_ASAP7_75t_L g13503 ( 
.A(n_13474),
.Y(n_13503)
);

INVx1_ASAP7_75t_L g13504 ( 
.A(n_13484),
.Y(n_13504)
);

AND2x2_ASAP7_75t_L g13505 ( 
.A(n_13495),
.B(n_13494),
.Y(n_13505)
);

INVx1_ASAP7_75t_L g13506 ( 
.A(n_13486),
.Y(n_13506)
);

INVx2_ASAP7_75t_L g13507 ( 
.A(n_13487),
.Y(n_13507)
);

NAND4xp75_ASAP7_75t_L g13508 ( 
.A(n_13471),
.B(n_2165),
.C(n_2163),
.D(n_2164),
.Y(n_13508)
);

NAND2xp5_ASAP7_75t_L g13509 ( 
.A(n_13490),
.B(n_2164),
.Y(n_13509)
);

INVx1_ASAP7_75t_SL g13510 ( 
.A(n_13397),
.Y(n_13510)
);

AND2x2_ASAP7_75t_L g13511 ( 
.A(n_13376),
.B(n_2165),
.Y(n_13511)
);

INVx2_ASAP7_75t_SL g13512 ( 
.A(n_13411),
.Y(n_13512)
);

NAND2xp33_ASAP7_75t_SL g13513 ( 
.A(n_13413),
.B(n_2166),
.Y(n_13513)
);

INVx1_ASAP7_75t_L g13514 ( 
.A(n_13491),
.Y(n_13514)
);

AOI22x1_ASAP7_75t_SL g13515 ( 
.A1(n_13386),
.A2(n_2168),
.B1(n_2166),
.B2(n_2167),
.Y(n_13515)
);

NOR3xp33_ASAP7_75t_SL g13516 ( 
.A(n_13391),
.B(n_2167),
.C(n_2168),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_13497),
.Y(n_13517)
);

INVx2_ASAP7_75t_SL g13518 ( 
.A(n_13466),
.Y(n_13518)
);

INVx1_ASAP7_75t_SL g13519 ( 
.A(n_13425),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_13388),
.Y(n_13520)
);

XOR2xp5_ASAP7_75t_L g13521 ( 
.A(n_13392),
.B(n_2169),
.Y(n_13521)
);

AND2x4_ASAP7_75t_SL g13522 ( 
.A(n_13382),
.B(n_2169),
.Y(n_13522)
);

INVxp67_ASAP7_75t_SL g13523 ( 
.A(n_13432),
.Y(n_13523)
);

INVxp33_ASAP7_75t_SL g13524 ( 
.A(n_13416),
.Y(n_13524)
);

INVx1_ASAP7_75t_L g13525 ( 
.A(n_13404),
.Y(n_13525)
);

NOR3xp33_ASAP7_75t_SL g13526 ( 
.A(n_13387),
.B(n_2170),
.C(n_2171),
.Y(n_13526)
);

NAND2xp5_ASAP7_75t_L g13527 ( 
.A(n_13379),
.B(n_2170),
.Y(n_13527)
);

INVx2_ASAP7_75t_SL g13528 ( 
.A(n_13409),
.Y(n_13528)
);

NAND2xp5_ASAP7_75t_L g13529 ( 
.A(n_13422),
.B(n_2172),
.Y(n_13529)
);

AND2x2_ASAP7_75t_L g13530 ( 
.A(n_13374),
.B(n_2173),
.Y(n_13530)
);

NOR4xp25_ASAP7_75t_L g13531 ( 
.A(n_13459),
.B(n_2176),
.C(n_2174),
.D(n_2175),
.Y(n_13531)
);

INVx2_ASAP7_75t_SL g13532 ( 
.A(n_13423),
.Y(n_13532)
);

XOR2x2_ASAP7_75t_L g13533 ( 
.A(n_13443),
.B(n_2174),
.Y(n_13533)
);

AND2x2_ASAP7_75t_L g13534 ( 
.A(n_13407),
.B(n_2175),
.Y(n_13534)
);

HB1xp67_ASAP7_75t_L g13535 ( 
.A(n_13406),
.Y(n_13535)
);

XOR2x2_ASAP7_75t_L g13536 ( 
.A(n_13389),
.B(n_2176),
.Y(n_13536)
);

AND2x2_ASAP7_75t_L g13537 ( 
.A(n_13394),
.B(n_2177),
.Y(n_13537)
);

XNOR2xp5_ASAP7_75t_L g13538 ( 
.A(n_13380),
.B(n_2178),
.Y(n_13538)
);

NOR2xp33_ASAP7_75t_L g13539 ( 
.A(n_13460),
.B(n_2178),
.Y(n_13539)
);

NOR2x1_ASAP7_75t_R g13540 ( 
.A(n_13433),
.B(n_13476),
.Y(n_13540)
);

OR2x2_ASAP7_75t_L g13541 ( 
.A(n_13488),
.B(n_2179),
.Y(n_13541)
);

NOR3xp33_ASAP7_75t_SL g13542 ( 
.A(n_13381),
.B(n_2179),
.C(n_2180),
.Y(n_13542)
);

AND2x2_ASAP7_75t_L g13543 ( 
.A(n_13395),
.B(n_2180),
.Y(n_13543)
);

INVx2_ASAP7_75t_SL g13544 ( 
.A(n_13396),
.Y(n_13544)
);

INVx2_ASAP7_75t_L g13545 ( 
.A(n_13406),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_13489),
.Y(n_13546)
);

OAI22xp33_ASAP7_75t_L g13547 ( 
.A1(n_13375),
.A2(n_2183),
.B1(n_2181),
.B2(n_2182),
.Y(n_13547)
);

INVxp67_ASAP7_75t_SL g13548 ( 
.A(n_13437),
.Y(n_13548)
);

NAND4xp75_ASAP7_75t_L g13549 ( 
.A(n_13378),
.B(n_2184),
.C(n_2181),
.D(n_2182),
.Y(n_13549)
);

NAND4xp75_ASAP7_75t_L g13550 ( 
.A(n_13384),
.B(n_2186),
.C(n_2184),
.D(n_2185),
.Y(n_13550)
);

NAND4xp75_ASAP7_75t_L g13551 ( 
.A(n_13385),
.B(n_2187),
.C(n_2185),
.D(n_2186),
.Y(n_13551)
);

XNOR2xp5_ASAP7_75t_L g13552 ( 
.A(n_13383),
.B(n_2187),
.Y(n_13552)
);

INVx3_ASAP7_75t_L g13553 ( 
.A(n_13418),
.Y(n_13553)
);

NAND4xp75_ASAP7_75t_L g13554 ( 
.A(n_13390),
.B(n_2190),
.C(n_2188),
.D(n_2189),
.Y(n_13554)
);

INVxp67_ASAP7_75t_L g13555 ( 
.A(n_13449),
.Y(n_13555)
);

XNOR2x2_ASAP7_75t_L g13556 ( 
.A(n_13496),
.B(n_2188),
.Y(n_13556)
);

INVx3_ASAP7_75t_L g13557 ( 
.A(n_13399),
.Y(n_13557)
);

INVx1_ASAP7_75t_L g13558 ( 
.A(n_13402),
.Y(n_13558)
);

INVx1_ASAP7_75t_L g13559 ( 
.A(n_13444),
.Y(n_13559)
);

AND2x2_ASAP7_75t_L g13560 ( 
.A(n_13435),
.B(n_2189),
.Y(n_13560)
);

NAND2xp5_ASAP7_75t_L g13561 ( 
.A(n_13467),
.B(n_2190),
.Y(n_13561)
);

XNOR2xp5_ASAP7_75t_L g13562 ( 
.A(n_13448),
.B(n_2191),
.Y(n_13562)
);

XNOR2x2_ASAP7_75t_L g13563 ( 
.A(n_13405),
.B(n_2192),
.Y(n_13563)
);

NAND4xp75_ASAP7_75t_L g13564 ( 
.A(n_13408),
.B(n_13430),
.C(n_13393),
.D(n_13421),
.Y(n_13564)
);

AND2x2_ASAP7_75t_L g13565 ( 
.A(n_13426),
.B(n_2192),
.Y(n_13565)
);

NAND2xp5_ASAP7_75t_L g13566 ( 
.A(n_13456),
.B(n_2193),
.Y(n_13566)
);

BUFx2_ASAP7_75t_L g13567 ( 
.A(n_13428),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_13400),
.Y(n_13568)
);

NAND4xp75_ASAP7_75t_L g13569 ( 
.A(n_13453),
.B(n_2195),
.C(n_2193),
.D(n_2194),
.Y(n_13569)
);

INVx1_ASAP7_75t_L g13570 ( 
.A(n_13410),
.Y(n_13570)
);

AND4x1_ASAP7_75t_L g13571 ( 
.A(n_13417),
.B(n_2197),
.C(n_2194),
.D(n_2196),
.Y(n_13571)
);

INVx2_ASAP7_75t_L g13572 ( 
.A(n_13470),
.Y(n_13572)
);

BUFx3_ASAP7_75t_L g13573 ( 
.A(n_13398),
.Y(n_13573)
);

XOR2x2_ASAP7_75t_L g13574 ( 
.A(n_13377),
.B(n_2197),
.Y(n_13574)
);

INVx4_ASAP7_75t_L g13575 ( 
.A(n_13445),
.Y(n_13575)
);

AND2x2_ASAP7_75t_L g13576 ( 
.A(n_13403),
.B(n_2198),
.Y(n_13576)
);

NAND4xp75_ASAP7_75t_L g13577 ( 
.A(n_13439),
.B(n_2200),
.C(n_2198),
.D(n_2199),
.Y(n_13577)
);

NAND4xp75_ASAP7_75t_SL g13578 ( 
.A(n_13438),
.B(n_2202),
.C(n_2199),
.D(n_2201),
.Y(n_13578)
);

AND2x2_ASAP7_75t_L g13579 ( 
.A(n_13401),
.B(n_2201),
.Y(n_13579)
);

INVx1_ASAP7_75t_L g13580 ( 
.A(n_13412),
.Y(n_13580)
);

XNOR2xp5_ASAP7_75t_L g13581 ( 
.A(n_13446),
.B(n_2202),
.Y(n_13581)
);

INVx1_ASAP7_75t_L g13582 ( 
.A(n_13472),
.Y(n_13582)
);

XNOR2x2_ASAP7_75t_L g13583 ( 
.A(n_13462),
.B(n_13447),
.Y(n_13583)
);

OR2x2_ASAP7_75t_L g13584 ( 
.A(n_13415),
.B(n_13436),
.Y(n_13584)
);

NAND4xp75_ASAP7_75t_L g13585 ( 
.A(n_13452),
.B(n_2205),
.C(n_2203),
.D(n_2204),
.Y(n_13585)
);

AND2x2_ASAP7_75t_L g13586 ( 
.A(n_13473),
.B(n_2203),
.Y(n_13586)
);

AND2x2_ASAP7_75t_L g13587 ( 
.A(n_13475),
.B(n_2204),
.Y(n_13587)
);

INVx2_ASAP7_75t_L g13588 ( 
.A(n_13419),
.Y(n_13588)
);

AND2x2_ASAP7_75t_L g13589 ( 
.A(n_13458),
.B(n_2205),
.Y(n_13589)
);

XNOR2xp5_ASAP7_75t_L g13590 ( 
.A(n_13434),
.B(n_2206),
.Y(n_13590)
);

INVx1_ASAP7_75t_L g13591 ( 
.A(n_13451),
.Y(n_13591)
);

NAND2xp33_ASAP7_75t_SL g13592 ( 
.A(n_13424),
.B(n_2206),
.Y(n_13592)
);

AND2x2_ASAP7_75t_L g13593 ( 
.A(n_13461),
.B(n_2208),
.Y(n_13593)
);

INVx1_ASAP7_75t_L g13594 ( 
.A(n_13442),
.Y(n_13594)
);

INVx1_ASAP7_75t_L g13595 ( 
.A(n_13478),
.Y(n_13595)
);

XNOR2xp5_ASAP7_75t_L g13596 ( 
.A(n_13440),
.B(n_2209),
.Y(n_13596)
);

INVx1_ASAP7_75t_SL g13597 ( 
.A(n_13457),
.Y(n_13597)
);

NAND3xp33_ASAP7_75t_L g13598 ( 
.A(n_13414),
.B(n_2210),
.C(n_2211),
.Y(n_13598)
);

NAND2xp5_ASAP7_75t_L g13599 ( 
.A(n_13469),
.B(n_2210),
.Y(n_13599)
);

XNOR2xp5_ASAP7_75t_L g13600 ( 
.A(n_13463),
.B(n_2212),
.Y(n_13600)
);

NAND4xp75_ASAP7_75t_SL g13601 ( 
.A(n_13464),
.B(n_2214),
.C(n_2212),
.D(n_2213),
.Y(n_13601)
);

AND2x2_ASAP7_75t_L g13602 ( 
.A(n_13429),
.B(n_2214),
.Y(n_13602)
);

INVx4_ASAP7_75t_L g13603 ( 
.A(n_13477),
.Y(n_13603)
);

NAND2xp5_ASAP7_75t_L g13604 ( 
.A(n_13479),
.B(n_2215),
.Y(n_13604)
);

NOR3xp33_ASAP7_75t_L g13605 ( 
.A(n_13455),
.B(n_2215),
.C(n_2216),
.Y(n_13605)
);

NAND2xp5_ASAP7_75t_L g13606 ( 
.A(n_13481),
.B(n_2216),
.Y(n_13606)
);

NOR2xp33_ASAP7_75t_L g13607 ( 
.A(n_13427),
.B(n_2217),
.Y(n_13607)
);

NAND4xp75_ASAP7_75t_L g13608 ( 
.A(n_13420),
.B(n_13431),
.C(n_13450),
.D(n_13482),
.Y(n_13608)
);

AND2x2_ASAP7_75t_L g13609 ( 
.A(n_13441),
.B(n_2217),
.Y(n_13609)
);

XOR2x2_ASAP7_75t_L g13610 ( 
.A(n_13465),
.B(n_2219),
.Y(n_13610)
);

INVx1_ASAP7_75t_L g13611 ( 
.A(n_13468),
.Y(n_13611)
);

NAND2xp5_ASAP7_75t_L g13612 ( 
.A(n_13454),
.B(n_2219),
.Y(n_13612)
);

NAND4xp75_ASAP7_75t_L g13613 ( 
.A(n_13480),
.B(n_2222),
.C(n_2220),
.D(n_2221),
.Y(n_13613)
);

NOR4xp25_ASAP7_75t_L g13614 ( 
.A(n_13483),
.B(n_2222),
.C(n_2220),
.D(n_2221),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_13373),
.Y(n_13615)
);

INVx2_ASAP7_75t_L g13616 ( 
.A(n_13487),
.Y(n_13616)
);

NAND4xp25_ASAP7_75t_L g13617 ( 
.A(n_13387),
.B(n_2225),
.C(n_2223),
.D(n_2224),
.Y(n_13617)
);

NOR3xp33_ASAP7_75t_L g13618 ( 
.A(n_13387),
.B(n_2224),
.C(n_2225),
.Y(n_13618)
);

HB1xp67_ASAP7_75t_L g13619 ( 
.A(n_13388),
.Y(n_13619)
);

INVxp67_ASAP7_75t_L g13620 ( 
.A(n_13474),
.Y(n_13620)
);

NAND4xp75_ASAP7_75t_SL g13621 ( 
.A(n_13387),
.B(n_2228),
.C(n_2226),
.D(n_2227),
.Y(n_13621)
);

AOI21xp5_ASAP7_75t_L g13622 ( 
.A1(n_13388),
.A2(n_2226),
.B(n_2229),
.Y(n_13622)
);

INVx1_ASAP7_75t_L g13623 ( 
.A(n_13373),
.Y(n_13623)
);

OAI22x1_ASAP7_75t_L g13624 ( 
.A1(n_13485),
.A2(n_2231),
.B1(n_2229),
.B2(n_2230),
.Y(n_13624)
);

XOR2x2_ASAP7_75t_L g13625 ( 
.A(n_13387),
.B(n_2230),
.Y(n_13625)
);

XOR2x2_ASAP7_75t_L g13626 ( 
.A(n_13387),
.B(n_2231),
.Y(n_13626)
);

INVx1_ASAP7_75t_L g13627 ( 
.A(n_13373),
.Y(n_13627)
);

HB1xp67_ASAP7_75t_L g13628 ( 
.A(n_13388),
.Y(n_13628)
);

XOR2xp5_ASAP7_75t_L g13629 ( 
.A(n_13487),
.B(n_2232),
.Y(n_13629)
);

BUFx3_ASAP7_75t_L g13630 ( 
.A(n_13397),
.Y(n_13630)
);

INVx1_ASAP7_75t_L g13631 ( 
.A(n_13373),
.Y(n_13631)
);

NOR3xp33_ASAP7_75t_SL g13632 ( 
.A(n_13391),
.B(n_2232),
.C(n_2233),
.Y(n_13632)
);

INVx4_ASAP7_75t_L g13633 ( 
.A(n_13487),
.Y(n_13633)
);

XOR2x2_ASAP7_75t_L g13634 ( 
.A(n_13387),
.B(n_2234),
.Y(n_13634)
);

NAND2x1_ASAP7_75t_SL g13635 ( 
.A(n_13388),
.B(n_2234),
.Y(n_13635)
);

NAND4xp75_ASAP7_75t_SL g13636 ( 
.A(n_13387),
.B(n_2237),
.C(n_2235),
.D(n_2236),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_13373),
.Y(n_13637)
);

INVx1_ASAP7_75t_SL g13638 ( 
.A(n_13493),
.Y(n_13638)
);

NAND2xp5_ASAP7_75t_L g13639 ( 
.A(n_13493),
.B(n_2236),
.Y(n_13639)
);

INVx1_ASAP7_75t_L g13640 ( 
.A(n_13373),
.Y(n_13640)
);

NAND2xp5_ASAP7_75t_L g13641 ( 
.A(n_13493),
.B(n_2237),
.Y(n_13641)
);

NAND3xp33_ASAP7_75t_L g13642 ( 
.A(n_13388),
.B(n_2238),
.C(n_2239),
.Y(n_13642)
);

OR2x2_ASAP7_75t_L g13643 ( 
.A(n_13493),
.B(n_2238),
.Y(n_13643)
);

INVx2_ASAP7_75t_L g13644 ( 
.A(n_13487),
.Y(n_13644)
);

AND2x2_ASAP7_75t_L g13645 ( 
.A(n_13485),
.B(n_2239),
.Y(n_13645)
);

AND2x2_ASAP7_75t_L g13646 ( 
.A(n_13485),
.B(n_2240),
.Y(n_13646)
);

INVx1_ASAP7_75t_L g13647 ( 
.A(n_13373),
.Y(n_13647)
);

OR2x2_ASAP7_75t_L g13648 ( 
.A(n_13493),
.B(n_2240),
.Y(n_13648)
);

NOR2xp33_ASAP7_75t_L g13649 ( 
.A(n_13524),
.B(n_2241),
.Y(n_13649)
);

NAND3xp33_ASAP7_75t_L g13650 ( 
.A(n_13513),
.B(n_2241),
.C(n_2242),
.Y(n_13650)
);

INVx1_ASAP7_75t_L g13651 ( 
.A(n_13635),
.Y(n_13651)
);

NOR2x1_ASAP7_75t_L g13652 ( 
.A(n_13508),
.B(n_2242),
.Y(n_13652)
);

XNOR2xp5_ASAP7_75t_L g13653 ( 
.A(n_13536),
.B(n_2243),
.Y(n_13653)
);

OAI221xp5_ASAP7_75t_L g13654 ( 
.A1(n_13523),
.A2(n_2246),
.B1(n_2244),
.B2(n_2245),
.C(n_2247),
.Y(n_13654)
);

NAND2xp5_ASAP7_75t_SL g13655 ( 
.A(n_13633),
.B(n_13512),
.Y(n_13655)
);

OAI221xp5_ASAP7_75t_L g13656 ( 
.A1(n_13548),
.A2(n_2246),
.B1(n_2244),
.B2(n_2245),
.C(n_2247),
.Y(n_13656)
);

NAND2xp5_ASAP7_75t_L g13657 ( 
.A(n_13518),
.B(n_2248),
.Y(n_13657)
);

NAND2xp5_ASAP7_75t_L g13658 ( 
.A(n_13638),
.B(n_2248),
.Y(n_13658)
);

NOR2x1_ASAP7_75t_L g13659 ( 
.A(n_13577),
.B(n_2249),
.Y(n_13659)
);

OAI22xp33_ASAP7_75t_L g13660 ( 
.A1(n_13510),
.A2(n_2251),
.B1(n_2249),
.B2(n_2250),
.Y(n_13660)
);

NAND2xp5_ASAP7_75t_L g13661 ( 
.A(n_13535),
.B(n_2251),
.Y(n_13661)
);

OAI22xp33_ASAP7_75t_L g13662 ( 
.A1(n_13619),
.A2(n_2254),
.B1(n_2252),
.B2(n_2253),
.Y(n_13662)
);

OAI22xp33_ASAP7_75t_L g13663 ( 
.A1(n_13628),
.A2(n_2254),
.B1(n_2252),
.B2(n_2253),
.Y(n_13663)
);

AO221x2_ASAP7_75t_L g13664 ( 
.A1(n_13521),
.A2(n_2257),
.B1(n_2255),
.B2(n_2256),
.C(n_2258),
.Y(n_13664)
);

NAND2xp5_ASAP7_75t_L g13665 ( 
.A(n_13553),
.B(n_2255),
.Y(n_13665)
);

OAI22xp33_ASAP7_75t_L g13666 ( 
.A1(n_13503),
.A2(n_2259),
.B1(n_2256),
.B2(n_2257),
.Y(n_13666)
);

AND2x4_ASAP7_75t_L g13667 ( 
.A(n_13630),
.B(n_2259),
.Y(n_13667)
);

NOR4xp25_ASAP7_75t_SL g13668 ( 
.A(n_13592),
.B(n_2262),
.C(n_2260),
.D(n_2261),
.Y(n_13668)
);

AOI21xp5_ASAP7_75t_L g13669 ( 
.A1(n_13620),
.A2(n_2260),
.B(n_2261),
.Y(n_13669)
);

AOI22xp5_ASAP7_75t_L g13670 ( 
.A1(n_13520),
.A2(n_2264),
.B1(n_2262),
.B2(n_2263),
.Y(n_13670)
);

NAND2xp5_ASAP7_75t_L g13671 ( 
.A(n_13505),
.B(n_2263),
.Y(n_13671)
);

BUFx3_ASAP7_75t_L g13672 ( 
.A(n_13567),
.Y(n_13672)
);

AO221x2_ASAP7_75t_L g13673 ( 
.A1(n_13502),
.A2(n_2266),
.B1(n_2264),
.B2(n_2265),
.C(n_2267),
.Y(n_13673)
);

AO221x2_ASAP7_75t_L g13674 ( 
.A1(n_13504),
.A2(n_2267),
.B1(n_2265),
.B2(n_2266),
.C(n_2268),
.Y(n_13674)
);

OR2x2_ASAP7_75t_L g13675 ( 
.A(n_13541),
.B(n_2268),
.Y(n_13675)
);

CKINVDCx5p33_ASAP7_75t_R g13676 ( 
.A(n_13515),
.Y(n_13676)
);

AND2x2_ASAP7_75t_L g13677 ( 
.A(n_13530),
.B(n_2269),
.Y(n_13677)
);

AND2x4_ASAP7_75t_L g13678 ( 
.A(n_13528),
.B(n_2269),
.Y(n_13678)
);

INVx2_ASAP7_75t_SL g13679 ( 
.A(n_13522),
.Y(n_13679)
);

NAND2xp5_ASAP7_75t_L g13680 ( 
.A(n_13519),
.B(n_2270),
.Y(n_13680)
);

NOR2xp33_ASAP7_75t_L g13681 ( 
.A(n_13575),
.B(n_2271),
.Y(n_13681)
);

NAND2xp5_ASAP7_75t_L g13682 ( 
.A(n_13544),
.B(n_2271),
.Y(n_13682)
);

OAI221xp5_ASAP7_75t_L g13683 ( 
.A1(n_13527),
.A2(n_2274),
.B1(n_2272),
.B2(n_2273),
.C(n_2275),
.Y(n_13683)
);

AOI22xp5_ASAP7_75t_L g13684 ( 
.A1(n_13507),
.A2(n_2276),
.B1(n_2273),
.B2(n_2274),
.Y(n_13684)
);

NAND2xp33_ASAP7_75t_SL g13685 ( 
.A(n_13542),
.B(n_2276),
.Y(n_13685)
);

CKINVDCx20_ASAP7_75t_R g13686 ( 
.A(n_13574),
.Y(n_13686)
);

NOR2xp33_ASAP7_75t_L g13687 ( 
.A(n_13603),
.B(n_2277),
.Y(n_13687)
);

OAI22xp33_ASAP7_75t_L g13688 ( 
.A1(n_13517),
.A2(n_2279),
.B1(n_2277),
.B2(n_2278),
.Y(n_13688)
);

NAND2xp5_ASAP7_75t_L g13689 ( 
.A(n_13534),
.B(n_2278),
.Y(n_13689)
);

NOR4xp25_ASAP7_75t_SL g13690 ( 
.A(n_13525),
.B(n_2281),
.C(n_2279),
.D(n_2280),
.Y(n_13690)
);

NOR2xp33_ASAP7_75t_L g13691 ( 
.A(n_13617),
.B(n_2280),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_13629),
.Y(n_13692)
);

OAI22xp33_ASAP7_75t_L g13693 ( 
.A1(n_13616),
.A2(n_2283),
.B1(n_2281),
.B2(n_2282),
.Y(n_13693)
);

NAND2xp5_ASAP7_75t_L g13694 ( 
.A(n_13532),
.B(n_2282),
.Y(n_13694)
);

AOI22xp5_ASAP7_75t_L g13695 ( 
.A1(n_13644),
.A2(n_2286),
.B1(n_2283),
.B2(n_2284),
.Y(n_13695)
);

OAI22xp33_ASAP7_75t_L g13696 ( 
.A1(n_13545),
.A2(n_2287),
.B1(n_2284),
.B2(n_2286),
.Y(n_13696)
);

AO221x2_ASAP7_75t_L g13697 ( 
.A1(n_13615),
.A2(n_2289),
.B1(n_2287),
.B2(n_2288),
.C(n_2290),
.Y(n_13697)
);

INVx1_ASAP7_75t_SL g13698 ( 
.A(n_13578),
.Y(n_13698)
);

OAI22xp33_ASAP7_75t_L g13699 ( 
.A1(n_13643),
.A2(n_2290),
.B1(n_2288),
.B2(n_2289),
.Y(n_13699)
);

AND2x4_ASAP7_75t_SL g13700 ( 
.A(n_13572),
.B(n_2291),
.Y(n_13700)
);

NAND2xp5_ASAP7_75t_L g13701 ( 
.A(n_13557),
.B(n_2291),
.Y(n_13701)
);

AOI22xp5_ASAP7_75t_SL g13702 ( 
.A1(n_13624),
.A2(n_2294),
.B1(n_2292),
.B2(n_2293),
.Y(n_13702)
);

NOR2x1_ASAP7_75t_L g13703 ( 
.A(n_13569),
.B(n_2292),
.Y(n_13703)
);

NOR2xp33_ASAP7_75t_L g13704 ( 
.A(n_13571),
.B(n_2294),
.Y(n_13704)
);

CKINVDCx20_ASAP7_75t_R g13705 ( 
.A(n_13625),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13538),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_13600),
.Y(n_13707)
);

NAND2xp5_ASAP7_75t_L g13708 ( 
.A(n_13560),
.B(n_2295),
.Y(n_13708)
);

AND2x4_ASAP7_75t_SL g13709 ( 
.A(n_13582),
.B(n_2295),
.Y(n_13709)
);

AOI22xp5_ASAP7_75t_L g13710 ( 
.A1(n_13558),
.A2(n_2298),
.B1(n_2296),
.B2(n_2297),
.Y(n_13710)
);

OAI22xp33_ASAP7_75t_L g13711 ( 
.A1(n_13648),
.A2(n_2299),
.B1(n_2296),
.B2(n_2298),
.Y(n_13711)
);

OAI221xp5_ASAP7_75t_L g13712 ( 
.A1(n_13516),
.A2(n_2302),
.B1(n_2300),
.B2(n_2301),
.C(n_2303),
.Y(n_13712)
);

INVx3_ASAP7_75t_L g13713 ( 
.A(n_13573),
.Y(n_13713)
);

INVx3_ASAP7_75t_L g13714 ( 
.A(n_13564),
.Y(n_13714)
);

OAI221xp5_ASAP7_75t_L g13715 ( 
.A1(n_13632),
.A2(n_2302),
.B1(n_2300),
.B2(n_2301),
.C(n_2303),
.Y(n_13715)
);

NAND2xp5_ASAP7_75t_L g13716 ( 
.A(n_13565),
.B(n_2304),
.Y(n_13716)
);

NAND2xp5_ASAP7_75t_L g13717 ( 
.A(n_13511),
.B(n_2305),
.Y(n_13717)
);

AO221x1_ASAP7_75t_L g13718 ( 
.A1(n_13547),
.A2(n_13631),
.B1(n_13637),
.B2(n_13627),
.C(n_13623),
.Y(n_13718)
);

AOI22xp5_ASAP7_75t_L g13719 ( 
.A1(n_13597),
.A2(n_13559),
.B1(n_13514),
.B2(n_13506),
.Y(n_13719)
);

NAND2xp5_ASAP7_75t_L g13720 ( 
.A(n_13498),
.B(n_13501),
.Y(n_13720)
);

NOR2x1_ASAP7_75t_L g13721 ( 
.A(n_13549),
.B(n_2305),
.Y(n_13721)
);

INVx2_ASAP7_75t_L g13722 ( 
.A(n_13563),
.Y(n_13722)
);

NAND2xp5_ASAP7_75t_L g13723 ( 
.A(n_13645),
.B(n_2306),
.Y(n_13723)
);

NAND2xp5_ASAP7_75t_L g13724 ( 
.A(n_13646),
.B(n_2308),
.Y(n_13724)
);

OAI22xp33_ASAP7_75t_L g13725 ( 
.A1(n_13639),
.A2(n_13641),
.B1(n_13647),
.B2(n_13640),
.Y(n_13725)
);

NAND2xp5_ASAP7_75t_L g13726 ( 
.A(n_13543),
.B(n_2308),
.Y(n_13726)
);

AO221x2_ASAP7_75t_L g13727 ( 
.A1(n_13570),
.A2(n_2312),
.B1(n_2310),
.B2(n_2311),
.C(n_2313),
.Y(n_13727)
);

NAND2xp5_ASAP7_75t_L g13728 ( 
.A(n_13576),
.B(n_2310),
.Y(n_13728)
);

INVx2_ASAP7_75t_SL g13729 ( 
.A(n_13537),
.Y(n_13729)
);

NAND2xp5_ASAP7_75t_L g13730 ( 
.A(n_13579),
.B(n_2311),
.Y(n_13730)
);

HB1xp67_ASAP7_75t_L g13731 ( 
.A(n_13601),
.Y(n_13731)
);

AND2x2_ASAP7_75t_L g13732 ( 
.A(n_13588),
.B(n_2312),
.Y(n_13732)
);

INVx2_ASAP7_75t_L g13733 ( 
.A(n_13584),
.Y(n_13733)
);

NOR2xp33_ASAP7_75t_L g13734 ( 
.A(n_13580),
.B(n_13591),
.Y(n_13734)
);

NAND2xp5_ASAP7_75t_L g13735 ( 
.A(n_13614),
.B(n_2314),
.Y(n_13735)
);

AND2x4_ASAP7_75t_L g13736 ( 
.A(n_13594),
.B(n_2314),
.Y(n_13736)
);

AND2x4_ASAP7_75t_L g13737 ( 
.A(n_13595),
.B(n_2315),
.Y(n_13737)
);

NOR2x1_ASAP7_75t_L g13738 ( 
.A(n_13550),
.B(n_2315),
.Y(n_13738)
);

OAI22xp33_ASAP7_75t_L g13739 ( 
.A1(n_13598),
.A2(n_2319),
.B1(n_2320),
.B2(n_2318),
.Y(n_13739)
);

NAND2xp33_ASAP7_75t_SL g13740 ( 
.A(n_13526),
.B(n_2316),
.Y(n_13740)
);

AND2x4_ASAP7_75t_L g13741 ( 
.A(n_13568),
.B(n_2318),
.Y(n_13741)
);

NAND2xp33_ASAP7_75t_SL g13742 ( 
.A(n_13529),
.B(n_2319),
.Y(n_13742)
);

NAND2xp5_ASAP7_75t_L g13743 ( 
.A(n_13586),
.B(n_2320),
.Y(n_13743)
);

AO221x2_ASAP7_75t_L g13744 ( 
.A1(n_13611),
.A2(n_2323),
.B1(n_2321),
.B2(n_2322),
.C(n_2324),
.Y(n_13744)
);

OR2x2_ASAP7_75t_L g13745 ( 
.A(n_13531),
.B(n_2321),
.Y(n_13745)
);

OR2x2_ASAP7_75t_L g13746 ( 
.A(n_13599),
.B(n_2322),
.Y(n_13746)
);

NAND2xp5_ASAP7_75t_L g13747 ( 
.A(n_13587),
.B(n_2324),
.Y(n_13747)
);

AO221x2_ASAP7_75t_L g13748 ( 
.A1(n_13546),
.A2(n_2327),
.B1(n_2325),
.B2(n_2326),
.C(n_2328),
.Y(n_13748)
);

INVxp67_ASAP7_75t_SL g13749 ( 
.A(n_13556),
.Y(n_13749)
);

OAI22xp5_ASAP7_75t_L g13750 ( 
.A1(n_13552),
.A2(n_2327),
.B1(n_2325),
.B2(n_2326),
.Y(n_13750)
);

NAND2xp5_ASAP7_75t_L g13751 ( 
.A(n_13500),
.B(n_2328),
.Y(n_13751)
);

AND2x2_ASAP7_75t_L g13752 ( 
.A(n_13589),
.B(n_2329),
.Y(n_13752)
);

INVxp33_ASAP7_75t_SL g13753 ( 
.A(n_13540),
.Y(n_13753)
);

OR2x2_ASAP7_75t_L g13754 ( 
.A(n_13612),
.B(n_2329),
.Y(n_13754)
);

AND2x2_ASAP7_75t_L g13755 ( 
.A(n_13593),
.B(n_2330),
.Y(n_13755)
);

AND2x2_ASAP7_75t_L g13756 ( 
.A(n_13602),
.B(n_2330),
.Y(n_13756)
);

AO221x2_ASAP7_75t_L g13757 ( 
.A1(n_13642),
.A2(n_2333),
.B1(n_2331),
.B2(n_2332),
.C(n_2334),
.Y(n_13757)
);

NOR2x1_ASAP7_75t_L g13758 ( 
.A(n_13551),
.B(n_2332),
.Y(n_13758)
);

INVx2_ASAP7_75t_SL g13759 ( 
.A(n_13609),
.Y(n_13759)
);

NAND2xp5_ASAP7_75t_L g13760 ( 
.A(n_13622),
.B(n_2333),
.Y(n_13760)
);

AO221x2_ASAP7_75t_L g13761 ( 
.A1(n_13509),
.A2(n_2338),
.B1(n_2334),
.B2(n_2336),
.C(n_2339),
.Y(n_13761)
);

AND2x2_ASAP7_75t_L g13762 ( 
.A(n_13533),
.B(n_2336),
.Y(n_13762)
);

NAND2xp5_ASAP7_75t_L g13763 ( 
.A(n_13590),
.B(n_2338),
.Y(n_13763)
);

OAI22xp33_ASAP7_75t_L g13764 ( 
.A1(n_13604),
.A2(n_2341),
.B1(n_2342),
.B2(n_2340),
.Y(n_13764)
);

NAND2xp33_ASAP7_75t_R g13765 ( 
.A(n_13539),
.B(n_2339),
.Y(n_13765)
);

NAND2xp5_ASAP7_75t_L g13766 ( 
.A(n_13596),
.B(n_2341),
.Y(n_13766)
);

NAND2xp33_ASAP7_75t_SL g13767 ( 
.A(n_13562),
.B(n_2343),
.Y(n_13767)
);

NAND2xp5_ASAP7_75t_L g13768 ( 
.A(n_13581),
.B(n_2343),
.Y(n_13768)
);

INVx1_ASAP7_75t_L g13769 ( 
.A(n_13626),
.Y(n_13769)
);

CKINVDCx20_ASAP7_75t_R g13770 ( 
.A(n_13634),
.Y(n_13770)
);

AOI22xp5_ASAP7_75t_L g13771 ( 
.A1(n_13555),
.A2(n_3371),
.B1(n_3372),
.B2(n_3370),
.Y(n_13771)
);

NAND2xp5_ASAP7_75t_L g13772 ( 
.A(n_13618),
.B(n_2344),
.Y(n_13772)
);

BUFx2_ASAP7_75t_L g13773 ( 
.A(n_13566),
.Y(n_13773)
);

NAND2xp5_ASAP7_75t_L g13774 ( 
.A(n_13585),
.B(n_2344),
.Y(n_13774)
);

NAND2xp5_ASAP7_75t_L g13775 ( 
.A(n_13554),
.B(n_2345),
.Y(n_13775)
);

NOR2x1_ASAP7_75t_L g13776 ( 
.A(n_13613),
.B(n_2345),
.Y(n_13776)
);

NAND2xp5_ASAP7_75t_L g13777 ( 
.A(n_13605),
.B(n_2346),
.Y(n_13777)
);

NAND2xp33_ASAP7_75t_SL g13778 ( 
.A(n_13499),
.B(n_2346),
.Y(n_13778)
);

AO221x2_ASAP7_75t_L g13779 ( 
.A1(n_13561),
.A2(n_2350),
.B1(n_2347),
.B2(n_2349),
.C(n_2351),
.Y(n_13779)
);

CKINVDCx5p33_ASAP7_75t_R g13780 ( 
.A(n_13610),
.Y(n_13780)
);

INVx1_ASAP7_75t_L g13781 ( 
.A(n_13606),
.Y(n_13781)
);

AO221x2_ASAP7_75t_L g13782 ( 
.A1(n_13583),
.A2(n_2350),
.B1(n_2347),
.B2(n_2349),
.C(n_2351),
.Y(n_13782)
);

OAI22xp33_ASAP7_75t_L g13783 ( 
.A1(n_13607),
.A2(n_2354),
.B1(n_2355),
.B2(n_2353),
.Y(n_13783)
);

NAND2xp5_ASAP7_75t_L g13784 ( 
.A(n_13608),
.B(n_2352),
.Y(n_13784)
);

INVx1_ASAP7_75t_L g13785 ( 
.A(n_13621),
.Y(n_13785)
);

NAND2xp5_ASAP7_75t_L g13786 ( 
.A(n_13636),
.B(n_2352),
.Y(n_13786)
);

CKINVDCx20_ASAP7_75t_R g13787 ( 
.A(n_13536),
.Y(n_13787)
);

AO221x2_ASAP7_75t_L g13788 ( 
.A1(n_13521),
.A2(n_2355),
.B1(n_2353),
.B2(n_2354),
.C(n_2356),
.Y(n_13788)
);

NAND2xp5_ASAP7_75t_L g13789 ( 
.A(n_13523),
.B(n_2357),
.Y(n_13789)
);

OAI22xp33_ASAP7_75t_L g13790 ( 
.A1(n_13633),
.A2(n_2359),
.B1(n_2360),
.B2(n_2358),
.Y(n_13790)
);

OAI221xp5_ASAP7_75t_L g13791 ( 
.A1(n_13513),
.A2(n_2359),
.B1(n_2357),
.B2(n_2358),
.C(n_2361),
.Y(n_13791)
);

NOR2x1_ASAP7_75t_L g13792 ( 
.A(n_13650),
.B(n_2361),
.Y(n_13792)
);

INVx1_ASAP7_75t_SL g13793 ( 
.A(n_13702),
.Y(n_13793)
);

NAND4xp25_ASAP7_75t_SL g13794 ( 
.A(n_13719),
.B(n_2364),
.C(n_2362),
.D(n_2363),
.Y(n_13794)
);

NAND2xp5_ASAP7_75t_L g13795 ( 
.A(n_13676),
.B(n_2362),
.Y(n_13795)
);

OR2x2_ASAP7_75t_L g13796 ( 
.A(n_13651),
.B(n_2364),
.Y(n_13796)
);

OR2x6_ASAP7_75t_L g13797 ( 
.A(n_13679),
.B(n_2365),
.Y(n_13797)
);

NOR2x1_ASAP7_75t_L g13798 ( 
.A(n_13672),
.B(n_2365),
.Y(n_13798)
);

OR2x2_ASAP7_75t_L g13799 ( 
.A(n_13722),
.B(n_2366),
.Y(n_13799)
);

NAND3xp33_ASAP7_75t_L g13800 ( 
.A(n_13685),
.B(n_2366),
.C(n_2367),
.Y(n_13800)
);

NAND2xp5_ASAP7_75t_L g13801 ( 
.A(n_13678),
.B(n_2368),
.Y(n_13801)
);

NAND2xp5_ASAP7_75t_L g13802 ( 
.A(n_13749),
.B(n_2369),
.Y(n_13802)
);

INVxp67_ASAP7_75t_SL g13803 ( 
.A(n_13659),
.Y(n_13803)
);

INVxp67_ASAP7_75t_L g13804 ( 
.A(n_13704),
.Y(n_13804)
);

NOR2xp33_ASAP7_75t_L g13805 ( 
.A(n_13791),
.B(n_2370),
.Y(n_13805)
);

AND2x2_ASAP7_75t_L g13806 ( 
.A(n_13762),
.B(n_2371),
.Y(n_13806)
);

NAND2xp33_ASAP7_75t_SL g13807 ( 
.A(n_13668),
.B(n_2371),
.Y(n_13807)
);

AND2x2_ASAP7_75t_L g13808 ( 
.A(n_13733),
.B(n_2372),
.Y(n_13808)
);

NAND2xp5_ASAP7_75t_L g13809 ( 
.A(n_13782),
.B(n_13700),
.Y(n_13809)
);

OR2x2_ASAP7_75t_L g13810 ( 
.A(n_13745),
.B(n_2372),
.Y(n_13810)
);

NAND2xp5_ASAP7_75t_L g13811 ( 
.A(n_13782),
.B(n_2373),
.Y(n_13811)
);

OR2x2_ASAP7_75t_L g13812 ( 
.A(n_13675),
.B(n_2373),
.Y(n_13812)
);

AND2x2_ASAP7_75t_L g13813 ( 
.A(n_13698),
.B(n_2374),
.Y(n_13813)
);

BUFx2_ASAP7_75t_L g13814 ( 
.A(n_13652),
.Y(n_13814)
);

CKINVDCx16_ASAP7_75t_R g13815 ( 
.A(n_13787),
.Y(n_13815)
);

AND2x2_ASAP7_75t_L g13816 ( 
.A(n_13731),
.B(n_13713),
.Y(n_13816)
);

INVx1_ASAP7_75t_L g13817 ( 
.A(n_13677),
.Y(n_13817)
);

NOR2xp33_ASAP7_75t_L g13818 ( 
.A(n_13753),
.B(n_2374),
.Y(n_13818)
);

AND2x2_ASAP7_75t_L g13819 ( 
.A(n_13714),
.B(n_2375),
.Y(n_13819)
);

AND2x2_ASAP7_75t_L g13820 ( 
.A(n_13785),
.B(n_2376),
.Y(n_13820)
);

INVx1_ASAP7_75t_L g13821 ( 
.A(n_13673),
.Y(n_13821)
);

AOI22xp33_ASAP7_75t_L g13822 ( 
.A1(n_13718),
.A2(n_2378),
.B1(n_2376),
.B2(n_2377),
.Y(n_13822)
);

NAND4xp25_ASAP7_75t_L g13823 ( 
.A(n_13734),
.B(n_2379),
.C(n_2377),
.D(n_2378),
.Y(n_13823)
);

NAND2xp5_ASAP7_75t_L g13824 ( 
.A(n_13709),
.B(n_2379),
.Y(n_13824)
);

INVx1_ASAP7_75t_L g13825 ( 
.A(n_13673),
.Y(n_13825)
);

NAND2xp5_ASAP7_75t_L g13826 ( 
.A(n_13667),
.B(n_2380),
.Y(n_13826)
);

AND2x2_ASAP7_75t_L g13827 ( 
.A(n_13732),
.B(n_2380),
.Y(n_13827)
);

CKINVDCx20_ASAP7_75t_R g13828 ( 
.A(n_13705),
.Y(n_13828)
);

AOI31xp67_ASAP7_75t_SL g13829 ( 
.A1(n_13784),
.A2(n_2383),
.A3(n_2381),
.B(n_2382),
.Y(n_13829)
);

AND2x2_ASAP7_75t_L g13830 ( 
.A(n_13729),
.B(n_2381),
.Y(n_13830)
);

OR2x2_ASAP7_75t_L g13831 ( 
.A(n_13735),
.B(n_2382),
.Y(n_13831)
);

BUFx2_ASAP7_75t_L g13832 ( 
.A(n_13721),
.Y(n_13832)
);

INVx1_ASAP7_75t_L g13833 ( 
.A(n_13674),
.Y(n_13833)
);

OR2x4_ASAP7_75t_L g13834 ( 
.A(n_13691),
.B(n_2383),
.Y(n_13834)
);

AOI21xp5_ASAP7_75t_L g13835 ( 
.A1(n_13655),
.A2(n_2384),
.B(n_2385),
.Y(n_13835)
);

AND2x2_ASAP7_75t_L g13836 ( 
.A(n_13738),
.B(n_2384),
.Y(n_13836)
);

NAND2xp5_ASAP7_75t_L g13837 ( 
.A(n_13664),
.B(n_2385),
.Y(n_13837)
);

AND2x2_ASAP7_75t_L g13838 ( 
.A(n_13758),
.B(n_2386),
.Y(n_13838)
);

AND2x2_ASAP7_75t_L g13839 ( 
.A(n_13703),
.B(n_2387),
.Y(n_13839)
);

INVx1_ASAP7_75t_L g13840 ( 
.A(n_13674),
.Y(n_13840)
);

AND2x4_ASAP7_75t_L g13841 ( 
.A(n_13752),
.B(n_2388),
.Y(n_13841)
);

AND2x2_ASAP7_75t_L g13842 ( 
.A(n_13759),
.B(n_2387),
.Y(n_13842)
);

INVx2_ASAP7_75t_L g13843 ( 
.A(n_13755),
.Y(n_13843)
);

NAND2xp33_ASAP7_75t_SL g13844 ( 
.A(n_13690),
.B(n_2390),
.Y(n_13844)
);

INVx1_ASAP7_75t_SL g13845 ( 
.A(n_13740),
.Y(n_13845)
);

INVx1_ASAP7_75t_L g13846 ( 
.A(n_13697),
.Y(n_13846)
);

NAND2x1_ASAP7_75t_L g13847 ( 
.A(n_13776),
.B(n_2392),
.Y(n_13847)
);

NOR3xp33_ASAP7_75t_L g13848 ( 
.A(n_13767),
.B(n_2395),
.C(n_2394),
.Y(n_13848)
);

NAND2xp67_ASAP7_75t_L g13849 ( 
.A(n_13756),
.B(n_2393),
.Y(n_13849)
);

NOR2xp33_ASAP7_75t_R g13850 ( 
.A(n_13765),
.B(n_2396),
.Y(n_13850)
);

INVx1_ASAP7_75t_L g13851 ( 
.A(n_13697),
.Y(n_13851)
);

INVx1_ASAP7_75t_L g13852 ( 
.A(n_13727),
.Y(n_13852)
);

OAI21xp33_ASAP7_75t_SL g13853 ( 
.A1(n_13720),
.A2(n_2395),
.B(n_2396),
.Y(n_13853)
);

HB1xp67_ASAP7_75t_L g13854 ( 
.A(n_13664),
.Y(n_13854)
);

NAND2xp5_ASAP7_75t_L g13855 ( 
.A(n_13788),
.B(n_2397),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_13769),
.B(n_2397),
.Y(n_13856)
);

AND2x2_ASAP7_75t_L g13857 ( 
.A(n_13692),
.B(n_2398),
.Y(n_13857)
);

INVx1_ASAP7_75t_L g13858 ( 
.A(n_13727),
.Y(n_13858)
);

INVx2_ASAP7_75t_L g13859 ( 
.A(n_13736),
.Y(n_13859)
);

HB1xp67_ASAP7_75t_L g13860 ( 
.A(n_13788),
.Y(n_13860)
);

OR2x2_ASAP7_75t_L g13861 ( 
.A(n_13657),
.B(n_2398),
.Y(n_13861)
);

AND2x2_ASAP7_75t_L g13862 ( 
.A(n_13706),
.B(n_2399),
.Y(n_13862)
);

AND2x2_ASAP7_75t_L g13863 ( 
.A(n_13707),
.B(n_2399),
.Y(n_13863)
);

NOR2xp33_ASAP7_75t_L g13864 ( 
.A(n_13712),
.B(n_2401),
.Y(n_13864)
);

NAND2xp33_ASAP7_75t_R g13865 ( 
.A(n_13780),
.B(n_3376),
.Y(n_13865)
);

INVx1_ASAP7_75t_L g13866 ( 
.A(n_13744),
.Y(n_13866)
);

OAI221xp5_ASAP7_75t_L g13867 ( 
.A1(n_13661),
.A2(n_13789),
.B1(n_13658),
.B2(n_13653),
.C(n_13778),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_13744),
.Y(n_13868)
);

OAI31xp33_ASAP7_75t_L g13869 ( 
.A1(n_13742),
.A2(n_2403),
.A3(n_2401),
.B(n_2402),
.Y(n_13869)
);

AND2x2_ASAP7_75t_L g13870 ( 
.A(n_13773),
.B(n_2403),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_13748),
.Y(n_13871)
);

AND5x1_ASAP7_75t_L g13872 ( 
.A(n_13649),
.B(n_2406),
.C(n_2404),
.D(n_2405),
.E(n_2408),
.Y(n_13872)
);

NAND2xp5_ASAP7_75t_L g13873 ( 
.A(n_13660),
.B(n_2404),
.Y(n_13873)
);

NAND2xp5_ASAP7_75t_L g13874 ( 
.A(n_13669),
.B(n_13662),
.Y(n_13874)
);

NAND2xp33_ASAP7_75t_R g13875 ( 
.A(n_13760),
.B(n_3364),
.Y(n_13875)
);

NAND2xp5_ASAP7_75t_L g13876 ( 
.A(n_13663),
.B(n_13761),
.Y(n_13876)
);

CKINVDCx16_ASAP7_75t_R g13877 ( 
.A(n_13770),
.Y(n_13877)
);

NAND2xp5_ASAP7_75t_L g13878 ( 
.A(n_13761),
.B(n_2405),
.Y(n_13878)
);

AND2x2_ASAP7_75t_L g13879 ( 
.A(n_13757),
.B(n_2408),
.Y(n_13879)
);

HB1xp67_ASAP7_75t_L g13880 ( 
.A(n_13779),
.Y(n_13880)
);

INVx1_ASAP7_75t_L g13881 ( 
.A(n_13748),
.Y(n_13881)
);

AND2x2_ASAP7_75t_L g13882 ( 
.A(n_13757),
.B(n_2409),
.Y(n_13882)
);

OR2x2_ASAP7_75t_L g13883 ( 
.A(n_13694),
.B(n_2409),
.Y(n_13883)
);

OR2x2_ASAP7_75t_L g13884 ( 
.A(n_13671),
.B(n_2410),
.Y(n_13884)
);

NAND2xp5_ASAP7_75t_L g13885 ( 
.A(n_13681),
.B(n_2410),
.Y(n_13885)
);

INVx1_ASAP7_75t_L g13886 ( 
.A(n_13786),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_13781),
.B(n_2411),
.Y(n_13887)
);

INVx1_ASAP7_75t_L g13888 ( 
.A(n_13779),
.Y(n_13888)
);

NAND2xp5_ASAP7_75t_L g13889 ( 
.A(n_13687),
.B(n_13688),
.Y(n_13889)
);

INVx1_ASAP7_75t_L g13890 ( 
.A(n_13689),
.Y(n_13890)
);

AND2x2_ASAP7_75t_L g13891 ( 
.A(n_13763),
.B(n_2412),
.Y(n_13891)
);

NAND2xp5_ASAP7_75t_L g13892 ( 
.A(n_13666),
.B(n_2412),
.Y(n_13892)
);

NOR2xp33_ASAP7_75t_R g13893 ( 
.A(n_13686),
.B(n_2414),
.Y(n_13893)
);

AND2x2_ASAP7_75t_L g13894 ( 
.A(n_13766),
.B(n_2413),
.Y(n_13894)
);

AND2x2_ASAP7_75t_L g13895 ( 
.A(n_13768),
.B(n_2413),
.Y(n_13895)
);

AND2x2_ASAP7_75t_L g13896 ( 
.A(n_13743),
.B(n_2414),
.Y(n_13896)
);

INVx1_ASAP7_75t_SL g13897 ( 
.A(n_13737),
.Y(n_13897)
);

AND2x2_ASAP7_75t_L g13898 ( 
.A(n_13747),
.B(n_2415),
.Y(n_13898)
);

NAND2xp33_ASAP7_75t_SL g13899 ( 
.A(n_13774),
.B(n_2415),
.Y(n_13899)
);

AOI31xp33_ASAP7_75t_L g13900 ( 
.A1(n_13680),
.A2(n_2424),
.A3(n_2432),
.B(n_2416),
.Y(n_13900)
);

INVx1_ASAP7_75t_L g13901 ( 
.A(n_13665),
.Y(n_13901)
);

NAND2xp5_ASAP7_75t_L g13902 ( 
.A(n_13790),
.B(n_2416),
.Y(n_13902)
);

INVx2_ASAP7_75t_L g13903 ( 
.A(n_13741),
.Y(n_13903)
);

NAND2xp5_ASAP7_75t_L g13904 ( 
.A(n_13696),
.B(n_13699),
.Y(n_13904)
);

INVx1_ASAP7_75t_L g13905 ( 
.A(n_13775),
.Y(n_13905)
);

NAND3xp33_ASAP7_75t_L g13906 ( 
.A(n_13715),
.B(n_2417),
.C(n_2418),
.Y(n_13906)
);

AND2x2_ASAP7_75t_L g13907 ( 
.A(n_13708),
.B(n_2417),
.Y(n_13907)
);

NOR2x1_ASAP7_75t_SL g13908 ( 
.A(n_13754),
.B(n_2418),
.Y(n_13908)
);

INVx2_ASAP7_75t_SL g13909 ( 
.A(n_13682),
.Y(n_13909)
);

INVx1_ASAP7_75t_SL g13910 ( 
.A(n_13701),
.Y(n_13910)
);

INVx1_ASAP7_75t_SL g13911 ( 
.A(n_13716),
.Y(n_13911)
);

NAND2xp5_ASAP7_75t_L g13912 ( 
.A(n_13711),
.B(n_2419),
.Y(n_13912)
);

INVx1_ASAP7_75t_L g13913 ( 
.A(n_13726),
.Y(n_13913)
);

INVx1_ASAP7_75t_L g13914 ( 
.A(n_13728),
.Y(n_13914)
);

NOR2xp67_ASAP7_75t_SL g13915 ( 
.A(n_13654),
.B(n_3361),
.Y(n_13915)
);

NAND2xp5_ASAP7_75t_L g13916 ( 
.A(n_13693),
.B(n_2420),
.Y(n_13916)
);

NAND2x1_ASAP7_75t_L g13917 ( 
.A(n_13717),
.B(n_2420),
.Y(n_13917)
);

HB1xp67_ASAP7_75t_L g13918 ( 
.A(n_13750),
.Y(n_13918)
);

NOR2xp33_ASAP7_75t_L g13919 ( 
.A(n_13730),
.B(n_2421),
.Y(n_13919)
);

OR2x2_ASAP7_75t_L g13920 ( 
.A(n_13746),
.B(n_2421),
.Y(n_13920)
);

INVx1_ASAP7_75t_SL g13921 ( 
.A(n_13723),
.Y(n_13921)
);

INVx1_ASAP7_75t_L g13922 ( 
.A(n_13724),
.Y(n_13922)
);

INVx1_ASAP7_75t_L g13923 ( 
.A(n_13751),
.Y(n_13923)
);

NAND2x1p5_ASAP7_75t_L g13924 ( 
.A(n_13670),
.B(n_2423),
.Y(n_13924)
);

NOR2xp33_ASAP7_75t_L g13925 ( 
.A(n_13683),
.B(n_2422),
.Y(n_13925)
);

INVx4_ASAP7_75t_L g13926 ( 
.A(n_13725),
.Y(n_13926)
);

AND2x4_ASAP7_75t_SL g13927 ( 
.A(n_13828),
.B(n_13710),
.Y(n_13927)
);

OR2x2_ASAP7_75t_L g13928 ( 
.A(n_13815),
.B(n_13772),
.Y(n_13928)
);

INVx1_ASAP7_75t_L g13929 ( 
.A(n_13880),
.Y(n_13929)
);

INVx1_ASAP7_75t_L g13930 ( 
.A(n_13854),
.Y(n_13930)
);

INVx1_ASAP7_75t_L g13931 ( 
.A(n_13860),
.Y(n_13931)
);

HB1xp67_ASAP7_75t_L g13932 ( 
.A(n_13797),
.Y(n_13932)
);

AND2x2_ASAP7_75t_L g13933 ( 
.A(n_13877),
.B(n_13777),
.Y(n_13933)
);

AND3x2_ASAP7_75t_L g13934 ( 
.A(n_13814),
.B(n_13764),
.C(n_13783),
.Y(n_13934)
);

INVx2_ASAP7_75t_L g13935 ( 
.A(n_13797),
.Y(n_13935)
);

INVx1_ASAP7_75t_SL g13936 ( 
.A(n_13807),
.Y(n_13936)
);

NAND2xp5_ASAP7_75t_L g13937 ( 
.A(n_13879),
.B(n_13882),
.Y(n_13937)
);

AND2x2_ASAP7_75t_L g13938 ( 
.A(n_13813),
.B(n_13684),
.Y(n_13938)
);

AOI22xp33_ASAP7_75t_L g13939 ( 
.A1(n_13926),
.A2(n_13739),
.B1(n_13656),
.B2(n_13695),
.Y(n_13939)
);

NAND2xp5_ASAP7_75t_L g13940 ( 
.A(n_13793),
.B(n_13771),
.Y(n_13940)
);

NOR2xp33_ASAP7_75t_L g13941 ( 
.A(n_13926),
.B(n_2422),
.Y(n_13941)
);

OR2x2_ASAP7_75t_L g13942 ( 
.A(n_13844),
.B(n_2423),
.Y(n_13942)
);

INVx2_ASAP7_75t_L g13943 ( 
.A(n_13799),
.Y(n_13943)
);

OA21x2_ASAP7_75t_L g13944 ( 
.A1(n_13822),
.A2(n_2424),
.B(n_2425),
.Y(n_13944)
);

AND2x2_ASAP7_75t_L g13945 ( 
.A(n_13806),
.B(n_2425),
.Y(n_13945)
);

AOI22xp33_ASAP7_75t_L g13946 ( 
.A1(n_13832),
.A2(n_2428),
.B1(n_2426),
.B2(n_2427),
.Y(n_13946)
);

AND2x2_ASAP7_75t_L g13947 ( 
.A(n_13856),
.B(n_2426),
.Y(n_13947)
);

INVx1_ASAP7_75t_L g13948 ( 
.A(n_13849),
.Y(n_13948)
);

NAND2xp5_ASAP7_75t_L g13949 ( 
.A(n_13852),
.B(n_13858),
.Y(n_13949)
);

INVx1_ASAP7_75t_L g13950 ( 
.A(n_13795),
.Y(n_13950)
);

INVx1_ASAP7_75t_L g13951 ( 
.A(n_13809),
.Y(n_13951)
);

CKINVDCx14_ASAP7_75t_R g13952 ( 
.A(n_13850),
.Y(n_13952)
);

INVx1_ASAP7_75t_SL g13953 ( 
.A(n_13893),
.Y(n_13953)
);

INVxp67_ASAP7_75t_SL g13954 ( 
.A(n_13798),
.Y(n_13954)
);

NOR2x1p5_ASAP7_75t_L g13955 ( 
.A(n_13847),
.B(n_3368),
.Y(n_13955)
);

INVx1_ASAP7_75t_L g13956 ( 
.A(n_13837),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_13855),
.Y(n_13957)
);

INVx1_ASAP7_75t_L g13958 ( 
.A(n_13802),
.Y(n_13958)
);

AND2x2_ASAP7_75t_L g13959 ( 
.A(n_13863),
.B(n_2427),
.Y(n_13959)
);

INVx2_ASAP7_75t_L g13960 ( 
.A(n_13841),
.Y(n_13960)
);

AND2x2_ASAP7_75t_L g13961 ( 
.A(n_13862),
.B(n_2428),
.Y(n_13961)
);

AOI22xp5_ASAP7_75t_L g13962 ( 
.A1(n_13816),
.A2(n_2431),
.B1(n_2429),
.B2(n_2430),
.Y(n_13962)
);

INVx1_ASAP7_75t_SL g13963 ( 
.A(n_13836),
.Y(n_13963)
);

AND2x2_ASAP7_75t_L g13964 ( 
.A(n_13820),
.B(n_2430),
.Y(n_13964)
);

NAND3x1_ASAP7_75t_L g13965 ( 
.A(n_13811),
.B(n_2431),
.C(n_2432),
.Y(n_13965)
);

INVx1_ASAP7_75t_L g13966 ( 
.A(n_13878),
.Y(n_13966)
);

HB1xp67_ASAP7_75t_L g13967 ( 
.A(n_13888),
.Y(n_13967)
);

INVx1_ASAP7_75t_L g13968 ( 
.A(n_13908),
.Y(n_13968)
);

CKINVDCx16_ASAP7_75t_R g13969 ( 
.A(n_13865),
.Y(n_13969)
);

AND2x4_ASAP7_75t_L g13970 ( 
.A(n_13859),
.B(n_2433),
.Y(n_13970)
);

INVx2_ASAP7_75t_L g13971 ( 
.A(n_13841),
.Y(n_13971)
);

AND2x2_ASAP7_75t_L g13972 ( 
.A(n_13857),
.B(n_2433),
.Y(n_13972)
);

INVxp67_ASAP7_75t_L g13973 ( 
.A(n_13818),
.Y(n_13973)
);

OR2x2_ASAP7_75t_L g13974 ( 
.A(n_13866),
.B(n_13868),
.Y(n_13974)
);

INVx1_ASAP7_75t_SL g13975 ( 
.A(n_13838),
.Y(n_13975)
);

INVx1_ASAP7_75t_L g13976 ( 
.A(n_13796),
.Y(n_13976)
);

INVxp67_ASAP7_75t_L g13977 ( 
.A(n_13821),
.Y(n_13977)
);

INVx1_ASAP7_75t_L g13978 ( 
.A(n_13839),
.Y(n_13978)
);

HB1xp67_ASAP7_75t_L g13979 ( 
.A(n_13825),
.Y(n_13979)
);

INVxp67_ASAP7_75t_L g13980 ( 
.A(n_13833),
.Y(n_13980)
);

INVx1_ASAP7_75t_SL g13981 ( 
.A(n_13840),
.Y(n_13981)
);

AOI22xp5_ASAP7_75t_L g13982 ( 
.A1(n_13845),
.A2(n_2436),
.B1(n_2434),
.B2(n_2435),
.Y(n_13982)
);

AND2x2_ASAP7_75t_L g13983 ( 
.A(n_13897),
.B(n_2435),
.Y(n_13983)
);

AND2x2_ASAP7_75t_SL g13984 ( 
.A(n_13846),
.B(n_2437),
.Y(n_13984)
);

INVx1_ASAP7_75t_L g13985 ( 
.A(n_13808),
.Y(n_13985)
);

INVx1_ASAP7_75t_L g13986 ( 
.A(n_13851),
.Y(n_13986)
);

OAI22xp5_ASAP7_75t_L g13987 ( 
.A1(n_13800),
.A2(n_2439),
.B1(n_2437),
.B2(n_2438),
.Y(n_13987)
);

AOI22xp33_ASAP7_75t_L g13988 ( 
.A1(n_13871),
.A2(n_2442),
.B1(n_2438),
.B2(n_2441),
.Y(n_13988)
);

NAND2xp5_ASAP7_75t_L g13989 ( 
.A(n_13881),
.B(n_2442),
.Y(n_13989)
);

INVx1_ASAP7_75t_L g13990 ( 
.A(n_13827),
.Y(n_13990)
);

AOI22xp33_ASAP7_75t_L g13991 ( 
.A1(n_13848),
.A2(n_2445),
.B1(n_2443),
.B2(n_2444),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13830),
.Y(n_13992)
);

AOI22xp33_ASAP7_75t_L g13993 ( 
.A1(n_13886),
.A2(n_2445),
.B1(n_2443),
.B2(n_2444),
.Y(n_13993)
);

NAND2xp5_ASAP7_75t_L g13994 ( 
.A(n_13803),
.B(n_2446),
.Y(n_13994)
);

AOI22xp33_ASAP7_75t_L g13995 ( 
.A1(n_13819),
.A2(n_2449),
.B1(n_2447),
.B2(n_2448),
.Y(n_13995)
);

INVx1_ASAP7_75t_L g13996 ( 
.A(n_13842),
.Y(n_13996)
);

INVx1_ASAP7_75t_SL g13997 ( 
.A(n_13812),
.Y(n_13997)
);

INVx1_ASAP7_75t_L g13998 ( 
.A(n_13824),
.Y(n_13998)
);

AND2x2_ASAP7_75t_L g13999 ( 
.A(n_13843),
.B(n_2447),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_13870),
.B(n_2448),
.Y(n_14000)
);

INVx1_ASAP7_75t_L g14001 ( 
.A(n_13810),
.Y(n_14001)
);

AOI22xp33_ASAP7_75t_L g14002 ( 
.A1(n_13918),
.A2(n_2452),
.B1(n_2450),
.B2(n_2451),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13801),
.Y(n_14003)
);

INVx1_ASAP7_75t_SL g14004 ( 
.A(n_13876),
.Y(n_14004)
);

AND2x2_ASAP7_75t_L g14005 ( 
.A(n_13903),
.B(n_2450),
.Y(n_14005)
);

INVx1_ASAP7_75t_L g14006 ( 
.A(n_13826),
.Y(n_14006)
);

NAND2xp5_ASAP7_75t_L g14007 ( 
.A(n_13817),
.B(n_2451),
.Y(n_14007)
);

INVx1_ASAP7_75t_L g14008 ( 
.A(n_13900),
.Y(n_14008)
);

NOR3xp33_ASAP7_75t_L g14009 ( 
.A(n_13867),
.B(n_2452),
.C(n_2453),
.Y(n_14009)
);

NAND2xp5_ASAP7_75t_L g14010 ( 
.A(n_13887),
.B(n_2453),
.Y(n_14010)
);

NAND2xp5_ASAP7_75t_L g14011 ( 
.A(n_13896),
.B(n_2454),
.Y(n_14011)
);

AND2x4_ASAP7_75t_L g14012 ( 
.A(n_13872),
.B(n_2455),
.Y(n_14012)
);

OR2x2_ASAP7_75t_L g14013 ( 
.A(n_13794),
.B(n_2455),
.Y(n_14013)
);

NAND3xp33_ASAP7_75t_SL g14014 ( 
.A(n_13869),
.B(n_2456),
.C(n_2457),
.Y(n_14014)
);

CKINVDCx16_ASAP7_75t_R g14015 ( 
.A(n_13875),
.Y(n_14015)
);

INVx1_ASAP7_75t_L g14016 ( 
.A(n_13831),
.Y(n_14016)
);

NOR2xp33_ASAP7_75t_L g14017 ( 
.A(n_13823),
.B(n_2457),
.Y(n_14017)
);

INVx2_ASAP7_75t_SL g14018 ( 
.A(n_13917),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_13891),
.B(n_2458),
.Y(n_14019)
);

HB1xp67_ASAP7_75t_L g14020 ( 
.A(n_13792),
.Y(n_14020)
);

AOI22xp33_ASAP7_75t_L g14021 ( 
.A1(n_13899),
.A2(n_2461),
.B1(n_2459),
.B2(n_2460),
.Y(n_14021)
);

AND2x2_ASAP7_75t_L g14022 ( 
.A(n_13894),
.B(n_2459),
.Y(n_14022)
);

NOR2xp33_ASAP7_75t_L g14023 ( 
.A(n_13853),
.B(n_2460),
.Y(n_14023)
);

AOI22xp33_ASAP7_75t_L g14024 ( 
.A1(n_13905),
.A2(n_2464),
.B1(n_2461),
.B2(n_2463),
.Y(n_14024)
);

OAI22xp5_ASAP7_75t_L g14025 ( 
.A1(n_13829),
.A2(n_2466),
.B1(n_2463),
.B2(n_2465),
.Y(n_14025)
);

OR2x2_ASAP7_75t_L g14026 ( 
.A(n_13920),
.B(n_2465),
.Y(n_14026)
);

AND2x2_ASAP7_75t_L g14027 ( 
.A(n_13895),
.B(n_2466),
.Y(n_14027)
);

INVxp67_ASAP7_75t_L g14028 ( 
.A(n_13915),
.Y(n_14028)
);

INVx2_ASAP7_75t_L g14029 ( 
.A(n_13884),
.Y(n_14029)
);

INVx1_ASAP7_75t_L g14030 ( 
.A(n_13873),
.Y(n_14030)
);

INVx1_ASAP7_75t_SL g14031 ( 
.A(n_13861),
.Y(n_14031)
);

AND2x4_ASAP7_75t_L g14032 ( 
.A(n_13898),
.B(n_2467),
.Y(n_14032)
);

INVx2_ASAP7_75t_L g14033 ( 
.A(n_13883),
.Y(n_14033)
);

AND2x2_ASAP7_75t_L g14034 ( 
.A(n_13907),
.B(n_2468),
.Y(n_14034)
);

INVx1_ASAP7_75t_L g14035 ( 
.A(n_13902),
.Y(n_14035)
);

INVx1_ASAP7_75t_L g14036 ( 
.A(n_13892),
.Y(n_14036)
);

NAND2xp5_ASAP7_75t_L g14037 ( 
.A(n_13835),
.B(n_13919),
.Y(n_14037)
);

NOR2xp33_ASAP7_75t_L g14038 ( 
.A(n_13804),
.B(n_2468),
.Y(n_14038)
);

AND2x2_ASAP7_75t_L g14039 ( 
.A(n_13864),
.B(n_2469),
.Y(n_14039)
);

AND2x2_ASAP7_75t_L g14040 ( 
.A(n_13924),
.B(n_2470),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_13912),
.Y(n_14041)
);

AOI222xp33_ASAP7_75t_L g14042 ( 
.A1(n_13874),
.A2(n_2473),
.B1(n_2475),
.B2(n_2471),
.C1(n_2472),
.C2(n_2474),
.Y(n_14042)
);

INVx2_ASAP7_75t_L g14043 ( 
.A(n_13834),
.Y(n_14043)
);

NAND2x1_ASAP7_75t_L g14044 ( 
.A(n_13909),
.B(n_13890),
.Y(n_14044)
);

AND2x2_ASAP7_75t_L g14045 ( 
.A(n_13911),
.B(n_2472),
.Y(n_14045)
);

NAND2xp5_ASAP7_75t_SL g14046 ( 
.A(n_13916),
.B(n_2473),
.Y(n_14046)
);

INVx1_ASAP7_75t_L g14047 ( 
.A(n_13904),
.Y(n_14047)
);

INVx1_ASAP7_75t_L g14048 ( 
.A(n_13885),
.Y(n_14048)
);

NAND2xp5_ASAP7_75t_L g14049 ( 
.A(n_13921),
.B(n_2476),
.Y(n_14049)
);

NAND2xp5_ASAP7_75t_L g14050 ( 
.A(n_13805),
.B(n_2477),
.Y(n_14050)
);

AND2x4_ASAP7_75t_L g14051 ( 
.A(n_13913),
.B(n_2478),
.Y(n_14051)
);

INVx1_ASAP7_75t_L g14052 ( 
.A(n_13889),
.Y(n_14052)
);

OAI222xp33_ASAP7_75t_L g14053 ( 
.A1(n_13936),
.A2(n_13910),
.B1(n_13901),
.B2(n_13914),
.C1(n_13922),
.C2(n_13923),
.Y(n_14053)
);

AOI222xp33_ASAP7_75t_L g14054 ( 
.A1(n_13941),
.A2(n_13906),
.B1(n_13925),
.B2(n_2480),
.C1(n_2482),
.C2(n_2478),
.Y(n_14054)
);

INVx2_ASAP7_75t_SL g14055 ( 
.A(n_13955),
.Y(n_14055)
);

INVx1_ASAP7_75t_L g14056 ( 
.A(n_13942),
.Y(n_14056)
);

NOR2xp33_ASAP7_75t_L g14057 ( 
.A(n_13969),
.B(n_2479),
.Y(n_14057)
);

INVx1_ASAP7_75t_L g14058 ( 
.A(n_13932),
.Y(n_14058)
);

HB1xp67_ASAP7_75t_L g14059 ( 
.A(n_13944),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13944),
.Y(n_14060)
);

INVx1_ASAP7_75t_L g14061 ( 
.A(n_13945),
.Y(n_14061)
);

INVx1_ASAP7_75t_SL g14062 ( 
.A(n_13984),
.Y(n_14062)
);

OAI22xp33_ASAP7_75t_L g14063 ( 
.A1(n_14015),
.A2(n_2482),
.B1(n_2479),
.B2(n_2481),
.Y(n_14063)
);

NAND2xp5_ASAP7_75t_L g14064 ( 
.A(n_13970),
.B(n_14012),
.Y(n_14064)
);

INVxp67_ASAP7_75t_SL g14065 ( 
.A(n_13965),
.Y(n_14065)
);

AOI21xp5_ASAP7_75t_L g14066 ( 
.A1(n_13954),
.A2(n_2481),
.B(n_2483),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13983),
.B(n_2484),
.Y(n_14067)
);

OR2x2_ASAP7_75t_L g14068 ( 
.A(n_13968),
.B(n_2484),
.Y(n_14068)
);

NOR2xp67_ASAP7_75t_SL g14069 ( 
.A(n_14020),
.B(n_2485),
.Y(n_14069)
);

INVxp67_ASAP7_75t_L g14070 ( 
.A(n_14023),
.Y(n_14070)
);

INVx1_ASAP7_75t_L g14071 ( 
.A(n_13937),
.Y(n_14071)
);

OAI22xp5_ASAP7_75t_L g14072 ( 
.A1(n_13952),
.A2(n_2488),
.B1(n_2486),
.B2(n_2487),
.Y(n_14072)
);

AOI22xp5_ASAP7_75t_L g14073 ( 
.A1(n_13981),
.A2(n_2491),
.B1(n_2489),
.B2(n_2490),
.Y(n_14073)
);

O2A1O1Ixp33_ASAP7_75t_L g14074 ( 
.A1(n_13979),
.A2(n_2491),
.B(n_2489),
.C(n_2490),
.Y(n_14074)
);

OR2x2_ASAP7_75t_L g14075 ( 
.A(n_14018),
.B(n_2492),
.Y(n_14075)
);

AOI22xp5_ASAP7_75t_L g14076 ( 
.A1(n_14004),
.A2(n_2495),
.B1(n_2493),
.B2(n_2494),
.Y(n_14076)
);

OAI21xp5_ASAP7_75t_L g14077 ( 
.A1(n_13977),
.A2(n_2493),
.B(n_2494),
.Y(n_14077)
);

INVx1_ASAP7_75t_L g14078 ( 
.A(n_14005),
.Y(n_14078)
);

OR4x1_ASAP7_75t_L g14079 ( 
.A(n_13929),
.B(n_2497),
.C(n_2495),
.D(n_2496),
.Y(n_14079)
);

NAND2xp5_ASAP7_75t_SL g14080 ( 
.A(n_13960),
.B(n_2497),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13999),
.B(n_2498),
.Y(n_14081)
);

NOR2xp33_ASAP7_75t_L g14082 ( 
.A(n_13971),
.B(n_2498),
.Y(n_14082)
);

INVx2_ASAP7_75t_L g14083 ( 
.A(n_14026),
.Y(n_14083)
);

INVx1_ASAP7_75t_L g14084 ( 
.A(n_13967),
.Y(n_14084)
);

AOI22xp5_ASAP7_75t_L g14085 ( 
.A1(n_13930),
.A2(n_2501),
.B1(n_2499),
.B2(n_2500),
.Y(n_14085)
);

AND2x2_ASAP7_75t_L g14086 ( 
.A(n_13964),
.B(n_2499),
.Y(n_14086)
);

INVx1_ASAP7_75t_L g14087 ( 
.A(n_13947),
.Y(n_14087)
);

AND2x2_ASAP7_75t_L g14088 ( 
.A(n_13935),
.B(n_2501),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13959),
.Y(n_14089)
);

AOI22xp33_ASAP7_75t_L g14090 ( 
.A1(n_13931),
.A2(n_13986),
.B1(n_13951),
.B2(n_14047),
.Y(n_14090)
);

INVx1_ASAP7_75t_L g14091 ( 
.A(n_13961),
.Y(n_14091)
);

NAND2xp5_ASAP7_75t_L g14092 ( 
.A(n_13972),
.B(n_2503),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_14013),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13974),
.Y(n_14094)
);

INVx1_ASAP7_75t_L g14095 ( 
.A(n_13989),
.Y(n_14095)
);

NAND2xp5_ASAP7_75t_L g14096 ( 
.A(n_14032),
.B(n_2503),
.Y(n_14096)
);

AOI22xp5_ASAP7_75t_L g14097 ( 
.A1(n_13980),
.A2(n_2506),
.B1(n_2504),
.B2(n_2505),
.Y(n_14097)
);

OAI21xp5_ASAP7_75t_L g14098 ( 
.A1(n_13949),
.A2(n_2504),
.B(n_2505),
.Y(n_14098)
);

OR2x2_ASAP7_75t_L g14099 ( 
.A(n_13953),
.B(n_2506),
.Y(n_14099)
);

OAI22xp33_ASAP7_75t_L g14100 ( 
.A1(n_13994),
.A2(n_2509),
.B1(n_2507),
.B2(n_2508),
.Y(n_14100)
);

OAI22xp5_ASAP7_75t_L g14101 ( 
.A1(n_13939),
.A2(n_2510),
.B1(n_2507),
.B2(n_2508),
.Y(n_14101)
);

INVx1_ASAP7_75t_L g14102 ( 
.A(n_14000),
.Y(n_14102)
);

NAND2xp33_ASAP7_75t_L g14103 ( 
.A(n_14009),
.B(n_2510),
.Y(n_14103)
);

AOI22xp33_ASAP7_75t_L g14104 ( 
.A1(n_14014),
.A2(n_2513),
.B1(n_2511),
.B2(n_2512),
.Y(n_14104)
);

AOI21xp5_ASAP7_75t_SL g14105 ( 
.A1(n_14025),
.A2(n_2511),
.B(n_2514),
.Y(n_14105)
);

AOI32xp33_ASAP7_75t_L g14106 ( 
.A1(n_13927),
.A2(n_2533),
.A3(n_2541),
.B1(n_2525),
.B2(n_2515),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_L g14107 ( 
.A(n_13934),
.B(n_2515),
.Y(n_14107)
);

INVx1_ASAP7_75t_L g14108 ( 
.A(n_14034),
.Y(n_14108)
);

INVxp67_ASAP7_75t_L g14109 ( 
.A(n_14038),
.Y(n_14109)
);

INVx1_ASAP7_75t_L g14110 ( 
.A(n_14019),
.Y(n_14110)
);

AOI222xp33_ASAP7_75t_L g14111 ( 
.A1(n_14028),
.A2(n_2520),
.B1(n_2522),
.B2(n_2516),
.C1(n_2518),
.C2(n_2521),
.Y(n_14111)
);

INVx2_ASAP7_75t_L g14112 ( 
.A(n_14051),
.Y(n_14112)
);

NAND2xp5_ASAP7_75t_L g14113 ( 
.A(n_13988),
.B(n_2521),
.Y(n_14113)
);

NAND2xp5_ASAP7_75t_L g14114 ( 
.A(n_13948),
.B(n_14022),
.Y(n_14114)
);

OR2x6_ASAP7_75t_L g14115 ( 
.A(n_14044),
.B(n_2523),
.Y(n_14115)
);

OAI22xp5_ASAP7_75t_L g14116 ( 
.A1(n_14002),
.A2(n_2526),
.B1(n_2524),
.B2(n_2525),
.Y(n_14116)
);

INVx2_ASAP7_75t_L g14117 ( 
.A(n_14027),
.Y(n_14117)
);

OR2x2_ASAP7_75t_L g14118 ( 
.A(n_14007),
.B(n_2524),
.Y(n_14118)
);

NAND2xp5_ASAP7_75t_SL g14119 ( 
.A(n_14042),
.B(n_2527),
.Y(n_14119)
);

O2A1O1Ixp5_ASAP7_75t_L g14120 ( 
.A1(n_13940),
.A2(n_2530),
.B(n_2528),
.C(n_2529),
.Y(n_14120)
);

AOI222xp33_ASAP7_75t_L g14121 ( 
.A1(n_14052),
.A2(n_2531),
.B1(n_2533),
.B2(n_2528),
.C1(n_2529),
.C2(n_2532),
.Y(n_14121)
);

NAND2xp5_ASAP7_75t_L g14122 ( 
.A(n_14040),
.B(n_2531),
.Y(n_14122)
);

OAI22xp5_ASAP7_75t_SL g14123 ( 
.A1(n_14021),
.A2(n_2535),
.B1(n_2532),
.B2(n_2534),
.Y(n_14123)
);

OAI322xp33_ASAP7_75t_L g14124 ( 
.A1(n_13928),
.A2(n_2539),
.A3(n_2538),
.B1(n_2536),
.B2(n_2534),
.C1(n_2535),
.C2(n_2537),
.Y(n_14124)
);

OAI22xp5_ASAP7_75t_L g14125 ( 
.A1(n_13991),
.A2(n_2539),
.B1(n_2537),
.B2(n_2538),
.Y(n_14125)
);

INVx1_ASAP7_75t_SL g14126 ( 
.A(n_14045),
.Y(n_14126)
);

INVx2_ASAP7_75t_L g14127 ( 
.A(n_14039),
.Y(n_14127)
);

NAND2xp33_ASAP7_75t_L g14128 ( 
.A(n_14008),
.B(n_2540),
.Y(n_14128)
);

AO22x1_ASAP7_75t_L g14129 ( 
.A1(n_13990),
.A2(n_2543),
.B1(n_2540),
.B2(n_2542),
.Y(n_14129)
);

OAI22xp33_ASAP7_75t_L g14130 ( 
.A1(n_13982),
.A2(n_2544),
.B1(n_2542),
.B2(n_2543),
.Y(n_14130)
);

INVx1_ASAP7_75t_L g14131 ( 
.A(n_14010),
.Y(n_14131)
);

INVx2_ASAP7_75t_L g14132 ( 
.A(n_13938),
.Y(n_14132)
);

INVx1_ASAP7_75t_L g14133 ( 
.A(n_14049),
.Y(n_14133)
);

AND2x2_ASAP7_75t_L g14134 ( 
.A(n_13933),
.B(n_13963),
.Y(n_14134)
);

INVxp67_ASAP7_75t_SL g14135 ( 
.A(n_14011),
.Y(n_14135)
);

AOI221xp5_ASAP7_75t_L g14136 ( 
.A1(n_13975),
.A2(n_2546),
.B1(n_2544),
.B2(n_2545),
.C(n_2547),
.Y(n_14136)
);

INVxp67_ASAP7_75t_L g14137 ( 
.A(n_14017),
.Y(n_14137)
);

INVx2_ASAP7_75t_L g14138 ( 
.A(n_13992),
.Y(n_14138)
);

NAND2xp5_ASAP7_75t_L g14139 ( 
.A(n_13995),
.B(n_2545),
.Y(n_14139)
);

NAND2xp5_ASAP7_75t_L g14140 ( 
.A(n_13946),
.B(n_2546),
.Y(n_14140)
);

AOI22xp5_ASAP7_75t_L g14141 ( 
.A1(n_13996),
.A2(n_2550),
.B1(n_2548),
.B2(n_2549),
.Y(n_14141)
);

OAI21xp5_ASAP7_75t_L g14142 ( 
.A1(n_13973),
.A2(n_2549),
.B(n_2550),
.Y(n_14142)
);

AOI22xp33_ASAP7_75t_L g14143 ( 
.A1(n_14043),
.A2(n_2553),
.B1(n_2551),
.B2(n_2552),
.Y(n_14143)
);

NOR2xp33_ASAP7_75t_L g14144 ( 
.A(n_13997),
.B(n_2551),
.Y(n_14144)
);

OR2x2_ASAP7_75t_L g14145 ( 
.A(n_13978),
.B(n_2552),
.Y(n_14145)
);

OAI21xp33_ASAP7_75t_SL g14146 ( 
.A1(n_14046),
.A2(n_3369),
.B(n_3361),
.Y(n_14146)
);

INVx2_ASAP7_75t_L g14147 ( 
.A(n_13943),
.Y(n_14147)
);

AOI222xp33_ASAP7_75t_L g14148 ( 
.A1(n_13966),
.A2(n_2555),
.B1(n_2557),
.B2(n_2553),
.C1(n_2554),
.C2(n_2556),
.Y(n_14148)
);

A2O1A1Ixp33_ASAP7_75t_L g14149 ( 
.A1(n_13976),
.A2(n_2556),
.B(n_2554),
.C(n_2555),
.Y(n_14149)
);

INVx1_ASAP7_75t_SL g14150 ( 
.A(n_14031),
.Y(n_14150)
);

INVx1_ASAP7_75t_L g14151 ( 
.A(n_14050),
.Y(n_14151)
);

INVx1_ASAP7_75t_L g14152 ( 
.A(n_13987),
.Y(n_14152)
);

INVx1_ASAP7_75t_SL g14153 ( 
.A(n_14001),
.Y(n_14153)
);

INVxp67_ASAP7_75t_SL g14154 ( 
.A(n_13962),
.Y(n_14154)
);

OAI22xp5_ASAP7_75t_L g14155 ( 
.A1(n_13985),
.A2(n_2559),
.B1(n_2557),
.B2(n_2558),
.Y(n_14155)
);

NOR2xp33_ASAP7_75t_L g14156 ( 
.A(n_13956),
.B(n_2558),
.Y(n_14156)
);

OAI22xp33_ASAP7_75t_L g14157 ( 
.A1(n_13957),
.A2(n_2562),
.B1(n_2560),
.B2(n_2561),
.Y(n_14157)
);

INVx1_ASAP7_75t_L g14158 ( 
.A(n_14037),
.Y(n_14158)
);

OR2x2_ASAP7_75t_L g14159 ( 
.A(n_13950),
.B(n_13958),
.Y(n_14159)
);

AOI31xp33_ASAP7_75t_L g14160 ( 
.A1(n_14016),
.A2(n_2568),
.A3(n_2576),
.B(n_2560),
.Y(n_14160)
);

OAI21xp33_ASAP7_75t_L g14161 ( 
.A1(n_14030),
.A2(n_2561),
.B(n_2562),
.Y(n_14161)
);

NAND2xp5_ASAP7_75t_L g14162 ( 
.A(n_14024),
.B(n_2563),
.Y(n_14162)
);

OAI22xp5_ASAP7_75t_L g14163 ( 
.A1(n_14041),
.A2(n_2565),
.B1(n_2563),
.B2(n_2564),
.Y(n_14163)
);

OAI21xp33_ASAP7_75t_L g14164 ( 
.A1(n_14036),
.A2(n_2564),
.B(n_2565),
.Y(n_14164)
);

NAND2xp5_ASAP7_75t_L g14165 ( 
.A(n_13993),
.B(n_14029),
.Y(n_14165)
);

AOI222xp33_ASAP7_75t_L g14166 ( 
.A1(n_14035),
.A2(n_2568),
.B1(n_2570),
.B2(n_2566),
.C1(n_2567),
.C2(n_2569),
.Y(n_14166)
);

OAI322xp33_ASAP7_75t_L g14167 ( 
.A1(n_13998),
.A2(n_2575),
.A3(n_2574),
.B1(n_2572),
.B2(n_2569),
.C1(n_2571),
.C2(n_2573),
.Y(n_14167)
);

INVxp67_ASAP7_75t_L g14168 ( 
.A(n_14033),
.Y(n_14168)
);

INVx1_ASAP7_75t_L g14169 ( 
.A(n_14006),
.Y(n_14169)
);

INVxp67_ASAP7_75t_L g14170 ( 
.A(n_14003),
.Y(n_14170)
);

OR2x2_ASAP7_75t_L g14171 ( 
.A(n_14048),
.B(n_2571),
.Y(n_14171)
);

INVx1_ASAP7_75t_L g14172 ( 
.A(n_13942),
.Y(n_14172)
);

AND2x2_ASAP7_75t_L g14173 ( 
.A(n_13936),
.B(n_2572),
.Y(n_14173)
);

INVx1_ASAP7_75t_L g14174 ( 
.A(n_13942),
.Y(n_14174)
);

NAND2xp5_ASAP7_75t_L g14175 ( 
.A(n_13936),
.B(n_2574),
.Y(n_14175)
);

NOR2xp33_ASAP7_75t_L g14176 ( 
.A(n_13969),
.B(n_2575),
.Y(n_14176)
);

OR2x2_ASAP7_75t_L g14177 ( 
.A(n_13969),
.B(n_2576),
.Y(n_14177)
);

INVx3_ASAP7_75t_L g14178 ( 
.A(n_13970),
.Y(n_14178)
);

OAI22xp5_ASAP7_75t_L g14179 ( 
.A1(n_13936),
.A2(n_2579),
.B1(n_2577),
.B2(n_2578),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13936),
.B(n_2577),
.Y(n_14180)
);

OAI21xp33_ASAP7_75t_L g14181 ( 
.A1(n_14004),
.A2(n_2579),
.B(n_2580),
.Y(n_14181)
);

OAI32xp33_ASAP7_75t_L g14182 ( 
.A1(n_13942),
.A2(n_2582),
.A3(n_2580),
.B1(n_2581),
.B2(n_2583),
.Y(n_14182)
);

INVx1_ASAP7_75t_L g14183 ( 
.A(n_13942),
.Y(n_14183)
);

AOI22xp33_ASAP7_75t_L g14184 ( 
.A1(n_14084),
.A2(n_2584),
.B1(n_2585),
.B2(n_2582),
.Y(n_14184)
);

NOR2xp33_ASAP7_75t_L g14185 ( 
.A(n_14177),
.B(n_2581),
.Y(n_14185)
);

NAND2xp5_ASAP7_75t_L g14186 ( 
.A(n_14059),
.B(n_2585),
.Y(n_14186)
);

AND2x4_ASAP7_75t_L g14187 ( 
.A(n_14094),
.B(n_2584),
.Y(n_14187)
);

NAND2xp5_ASAP7_75t_SL g14188 ( 
.A(n_14060),
.B(n_2586),
.Y(n_14188)
);

AND2x2_ASAP7_75t_L g14189 ( 
.A(n_14173),
.B(n_2587),
.Y(n_14189)
);

INVx1_ASAP7_75t_L g14190 ( 
.A(n_14068),
.Y(n_14190)
);

OAI22xp5_ASAP7_75t_L g14191 ( 
.A1(n_14090),
.A2(n_2589),
.B1(n_2587),
.B2(n_2588),
.Y(n_14191)
);

INVx1_ASAP7_75t_L g14192 ( 
.A(n_14107),
.Y(n_14192)
);

INVxp67_ASAP7_75t_SL g14193 ( 
.A(n_14069),
.Y(n_14193)
);

O2A1O1Ixp33_ASAP7_75t_L g14194 ( 
.A1(n_14128),
.A2(n_14115),
.B(n_14120),
.C(n_14065),
.Y(n_14194)
);

AOI22xp5_ASAP7_75t_L g14195 ( 
.A1(n_14058),
.A2(n_2590),
.B1(n_2588),
.B2(n_2589),
.Y(n_14195)
);

INVx1_ASAP7_75t_L g14196 ( 
.A(n_14075),
.Y(n_14196)
);

NAND4xp75_ASAP7_75t_L g14197 ( 
.A(n_14180),
.B(n_2592),
.C(n_2590),
.D(n_2591),
.Y(n_14197)
);

INVxp67_ASAP7_75t_SL g14198 ( 
.A(n_14057),
.Y(n_14198)
);

A2O1A1Ixp33_ASAP7_75t_L g14199 ( 
.A1(n_14074),
.A2(n_2593),
.B(n_2591),
.C(n_2592),
.Y(n_14199)
);

OR2x2_ASAP7_75t_L g14200 ( 
.A(n_14115),
.B(n_2593),
.Y(n_14200)
);

OAI22xp5_ASAP7_75t_L g14201 ( 
.A1(n_14104),
.A2(n_2596),
.B1(n_2594),
.B2(n_2595),
.Y(n_14201)
);

OAI22xp33_ASAP7_75t_L g14202 ( 
.A1(n_14175),
.A2(n_2597),
.B1(n_2598),
.B2(n_2596),
.Y(n_14202)
);

AND4x1_ASAP7_75t_L g14203 ( 
.A(n_14176),
.B(n_2599),
.C(n_2595),
.D(n_2598),
.Y(n_14203)
);

INVx1_ASAP7_75t_L g14204 ( 
.A(n_14086),
.Y(n_14204)
);

INVx1_ASAP7_75t_L g14205 ( 
.A(n_14067),
.Y(n_14205)
);

OAI21xp33_ASAP7_75t_L g14206 ( 
.A1(n_14150),
.A2(n_2600),
.B(n_2601),
.Y(n_14206)
);

INVx2_ASAP7_75t_L g14207 ( 
.A(n_14079),
.Y(n_14207)
);

INVxp67_ASAP7_75t_L g14208 ( 
.A(n_14082),
.Y(n_14208)
);

NAND2xp5_ASAP7_75t_SL g14209 ( 
.A(n_14106),
.B(n_2600),
.Y(n_14209)
);

INVx2_ASAP7_75t_L g14210 ( 
.A(n_14145),
.Y(n_14210)
);

AOI22xp5_ASAP7_75t_L g14211 ( 
.A1(n_14153),
.A2(n_2603),
.B1(n_2601),
.B2(n_2602),
.Y(n_14211)
);

AND2x2_ASAP7_75t_L g14212 ( 
.A(n_14183),
.B(n_2603),
.Y(n_14212)
);

INVx2_ASAP7_75t_L g14213 ( 
.A(n_14171),
.Y(n_14213)
);

AOI221xp5_ASAP7_75t_L g14214 ( 
.A1(n_14053),
.A2(n_2606),
.B1(n_2604),
.B2(n_2605),
.C(n_2607),
.Y(n_14214)
);

OAI21xp5_ASAP7_75t_L g14215 ( 
.A1(n_14168),
.A2(n_2604),
.B(n_2605),
.Y(n_14215)
);

AOI22xp5_ASAP7_75t_L g14216 ( 
.A1(n_14132),
.A2(n_2609),
.B1(n_2607),
.B2(n_2608),
.Y(n_14216)
);

INVx2_ASAP7_75t_SL g14217 ( 
.A(n_14178),
.Y(n_14217)
);

NAND2xp5_ASAP7_75t_L g14218 ( 
.A(n_14129),
.B(n_2609),
.Y(n_14218)
);

NAND2xp5_ASAP7_75t_L g14219 ( 
.A(n_14088),
.B(n_2610),
.Y(n_14219)
);

NAND3xp33_ASAP7_75t_L g14220 ( 
.A(n_14054),
.B(n_2608),
.C(n_2610),
.Y(n_14220)
);

OAI22xp33_ASAP7_75t_L g14221 ( 
.A1(n_14099),
.A2(n_2613),
.B1(n_2614),
.B2(n_2612),
.Y(n_14221)
);

INVx1_ASAP7_75t_L g14222 ( 
.A(n_14064),
.Y(n_14222)
);

NOR2x1_ASAP7_75t_L g14223 ( 
.A(n_14178),
.B(n_14167),
.Y(n_14223)
);

INVx1_ASAP7_75t_L g14224 ( 
.A(n_14092),
.Y(n_14224)
);

AOI21xp5_ASAP7_75t_L g14225 ( 
.A1(n_14103),
.A2(n_2611),
.B(n_2612),
.Y(n_14225)
);

OAI221xp5_ASAP7_75t_L g14226 ( 
.A1(n_14181),
.A2(n_14146),
.B1(n_14062),
.B2(n_14144),
.C(n_14055),
.Y(n_14226)
);

NAND2xp5_ASAP7_75t_L g14227 ( 
.A(n_14160),
.B(n_2613),
.Y(n_14227)
);

INVx1_ASAP7_75t_L g14228 ( 
.A(n_14096),
.Y(n_14228)
);

AOI22xp33_ASAP7_75t_L g14229 ( 
.A1(n_14138),
.A2(n_2615),
.B1(n_2616),
.B2(n_2614),
.Y(n_14229)
);

AO32x1_ASAP7_75t_L g14230 ( 
.A1(n_14134),
.A2(n_2616),
.A3(n_2611),
.B1(n_2615),
.B2(n_2617),
.Y(n_14230)
);

OAI22xp33_ASAP7_75t_SL g14231 ( 
.A1(n_14056),
.A2(n_2625),
.B1(n_2633),
.B2(n_2617),
.Y(n_14231)
);

INVx2_ASAP7_75t_L g14232 ( 
.A(n_14118),
.Y(n_14232)
);

NAND2xp5_ASAP7_75t_L g14233 ( 
.A(n_14063),
.B(n_2619),
.Y(n_14233)
);

OR2x2_ASAP7_75t_L g14234 ( 
.A(n_14081),
.B(n_2618),
.Y(n_14234)
);

INVx2_ASAP7_75t_L g14235 ( 
.A(n_14117),
.Y(n_14235)
);

OR2x2_ASAP7_75t_L g14236 ( 
.A(n_14122),
.B(n_2618),
.Y(n_14236)
);

NOR3xp33_ASAP7_75t_L g14237 ( 
.A(n_14114),
.B(n_2621),
.C(n_2620),
.Y(n_14237)
);

INVx2_ASAP7_75t_L g14238 ( 
.A(n_14112),
.Y(n_14238)
);

CKINVDCx16_ASAP7_75t_R g14239 ( 
.A(n_14126),
.Y(n_14239)
);

NOR2xp33_ASAP7_75t_L g14240 ( 
.A(n_14161),
.B(n_2619),
.Y(n_14240)
);

AOI22xp5_ASAP7_75t_L g14241 ( 
.A1(n_14147),
.A2(n_2623),
.B1(n_2621),
.B2(n_2622),
.Y(n_14241)
);

INVx1_ASAP7_75t_L g14242 ( 
.A(n_14123),
.Y(n_14242)
);

INVxp67_ASAP7_75t_L g14243 ( 
.A(n_14156),
.Y(n_14243)
);

INVx1_ASAP7_75t_L g14244 ( 
.A(n_14172),
.Y(n_14244)
);

NOR2x1_ASAP7_75t_L g14245 ( 
.A(n_14124),
.B(n_3368),
.Y(n_14245)
);

OA21x2_ASAP7_75t_L g14246 ( 
.A1(n_14071),
.A2(n_2622),
.B(n_2623),
.Y(n_14246)
);

AOI221x1_ASAP7_75t_L g14247 ( 
.A1(n_14174),
.A2(n_2627),
.B1(n_2624),
.B2(n_2626),
.C(n_2628),
.Y(n_14247)
);

OAI32xp33_ASAP7_75t_L g14248 ( 
.A1(n_14113),
.A2(n_14140),
.A3(n_14162),
.B1(n_14139),
.B2(n_14165),
.Y(n_14248)
);

AOI211xp5_ASAP7_75t_SL g14249 ( 
.A1(n_14105),
.A2(n_2627),
.B(n_2624),
.C(n_2626),
.Y(n_14249)
);

NAND2xp5_ASAP7_75t_L g14250 ( 
.A(n_14066),
.B(n_2630),
.Y(n_14250)
);

INVx1_ASAP7_75t_L g14251 ( 
.A(n_14061),
.Y(n_14251)
);

OR2x2_ASAP7_75t_L g14252 ( 
.A(n_14087),
.B(n_2629),
.Y(n_14252)
);

INVx1_ASAP7_75t_L g14253 ( 
.A(n_14080),
.Y(n_14253)
);

HB1xp67_ASAP7_75t_L g14254 ( 
.A(n_14072),
.Y(n_14254)
);

AOI22xp33_ASAP7_75t_L g14255 ( 
.A1(n_14083),
.A2(n_2631),
.B1(n_2632),
.B2(n_2630),
.Y(n_14255)
);

NAND2xp5_ASAP7_75t_L g14256 ( 
.A(n_14073),
.B(n_2631),
.Y(n_14256)
);

OAI31xp33_ASAP7_75t_L g14257 ( 
.A1(n_14130),
.A2(n_14093),
.A3(n_14101),
.B(n_14125),
.Y(n_14257)
);

AOI21xp5_ASAP7_75t_L g14258 ( 
.A1(n_14119),
.A2(n_14154),
.B(n_14182),
.Y(n_14258)
);

OAI22xp5_ASAP7_75t_L g14259 ( 
.A1(n_14076),
.A2(n_2633),
.B1(n_2629),
.B2(n_2632),
.Y(n_14259)
);

INVxp67_ASAP7_75t_L g14260 ( 
.A(n_14111),
.Y(n_14260)
);

INVx2_ASAP7_75t_L g14261 ( 
.A(n_14089),
.Y(n_14261)
);

INVx1_ASAP7_75t_L g14262 ( 
.A(n_14091),
.Y(n_14262)
);

NAND2xp5_ASAP7_75t_L g14263 ( 
.A(n_14108),
.B(n_14110),
.Y(n_14263)
);

NOR2xp33_ASAP7_75t_L g14264 ( 
.A(n_14164),
.B(n_2634),
.Y(n_14264)
);

INVx1_ASAP7_75t_L g14265 ( 
.A(n_14078),
.Y(n_14265)
);

INVxp67_ASAP7_75t_SL g14266 ( 
.A(n_14157),
.Y(n_14266)
);

AOI221xp5_ASAP7_75t_L g14267 ( 
.A1(n_14070),
.A2(n_2637),
.B1(n_2635),
.B2(n_2636),
.C(n_2638),
.Y(n_14267)
);

INVx1_ASAP7_75t_L g14268 ( 
.A(n_14127),
.Y(n_14268)
);

OAI22xp5_ASAP7_75t_L g14269 ( 
.A1(n_14170),
.A2(n_2638),
.B1(n_2636),
.B2(n_2637),
.Y(n_14269)
);

NAND3xp33_ASAP7_75t_L g14270 ( 
.A(n_14098),
.B(n_2639),
.C(n_2640),
.Y(n_14270)
);

INVx1_ASAP7_75t_L g14271 ( 
.A(n_14077),
.Y(n_14271)
);

OAI21xp33_ASAP7_75t_L g14272 ( 
.A1(n_14152),
.A2(n_2639),
.B(n_2640),
.Y(n_14272)
);

INVx1_ASAP7_75t_L g14273 ( 
.A(n_14179),
.Y(n_14273)
);

INVx1_ASAP7_75t_L g14274 ( 
.A(n_14142),
.Y(n_14274)
);

AOI211xp5_ASAP7_75t_L g14275 ( 
.A1(n_14116),
.A2(n_14169),
.B(n_14100),
.C(n_14158),
.Y(n_14275)
);

INVx1_ASAP7_75t_L g14276 ( 
.A(n_14159),
.Y(n_14276)
);

INVx1_ASAP7_75t_L g14277 ( 
.A(n_14085),
.Y(n_14277)
);

INVx1_ASAP7_75t_L g14278 ( 
.A(n_14097),
.Y(n_14278)
);

NOR2x1_ASAP7_75t_L g14279 ( 
.A(n_14149),
.B(n_3371),
.Y(n_14279)
);

INVx1_ASAP7_75t_L g14280 ( 
.A(n_14135),
.Y(n_14280)
);

HB1xp67_ASAP7_75t_L g14281 ( 
.A(n_14155),
.Y(n_14281)
);

AND2x2_ASAP7_75t_SL g14282 ( 
.A(n_14133),
.B(n_14095),
.Y(n_14282)
);

AOI22xp33_ASAP7_75t_L g14283 ( 
.A1(n_14102),
.A2(n_2643),
.B1(n_2644),
.B2(n_2642),
.Y(n_14283)
);

INVx2_ASAP7_75t_L g14284 ( 
.A(n_14131),
.Y(n_14284)
);

NAND2xp5_ASAP7_75t_L g14285 ( 
.A(n_14121),
.B(n_2642),
.Y(n_14285)
);

INVx2_ASAP7_75t_L g14286 ( 
.A(n_14151),
.Y(n_14286)
);

INVx1_ASAP7_75t_L g14287 ( 
.A(n_14163),
.Y(n_14287)
);

AND2x2_ASAP7_75t_L g14288 ( 
.A(n_14109),
.B(n_2641),
.Y(n_14288)
);

OAI22xp33_ASAP7_75t_L g14289 ( 
.A1(n_14137),
.A2(n_2645),
.B1(n_2646),
.B2(n_2644),
.Y(n_14289)
);

INVx1_ASAP7_75t_L g14290 ( 
.A(n_14141),
.Y(n_14290)
);

OAI22xp5_ASAP7_75t_L g14291 ( 
.A1(n_14143),
.A2(n_2646),
.B1(n_2641),
.B2(n_2645),
.Y(n_14291)
);

INVx1_ASAP7_75t_L g14292 ( 
.A(n_14166),
.Y(n_14292)
);

INVx1_ASAP7_75t_L g14293 ( 
.A(n_14148),
.Y(n_14293)
);

OR2x2_ASAP7_75t_L g14294 ( 
.A(n_14136),
.B(n_2647),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_14200),
.Y(n_14295)
);

NAND2xp5_ASAP7_75t_L g14296 ( 
.A(n_14212),
.B(n_2647),
.Y(n_14296)
);

NAND2xp5_ASAP7_75t_L g14297 ( 
.A(n_14189),
.B(n_2648),
.Y(n_14297)
);

NAND2xp5_ASAP7_75t_L g14298 ( 
.A(n_14249),
.B(n_2648),
.Y(n_14298)
);

INVx1_ASAP7_75t_L g14299 ( 
.A(n_14186),
.Y(n_14299)
);

BUFx2_ASAP7_75t_L g14300 ( 
.A(n_14246),
.Y(n_14300)
);

INVx2_ASAP7_75t_L g14301 ( 
.A(n_14246),
.Y(n_14301)
);

NAND2xp5_ASAP7_75t_L g14302 ( 
.A(n_14239),
.B(n_2649),
.Y(n_14302)
);

AND2x2_ASAP7_75t_L g14303 ( 
.A(n_14193),
.B(n_2649),
.Y(n_14303)
);

INVx1_ASAP7_75t_SL g14304 ( 
.A(n_14197),
.Y(n_14304)
);

AOI22xp5_ASAP7_75t_L g14305 ( 
.A1(n_14217),
.A2(n_2658),
.B1(n_2666),
.B2(n_2650),
.Y(n_14305)
);

NAND2xp5_ASAP7_75t_L g14306 ( 
.A(n_14203),
.B(n_2651),
.Y(n_14306)
);

NAND2xp5_ASAP7_75t_L g14307 ( 
.A(n_14185),
.B(n_2651),
.Y(n_14307)
);

NAND2xp5_ASAP7_75t_L g14308 ( 
.A(n_14221),
.B(n_2652),
.Y(n_14308)
);

NOR2xp33_ASAP7_75t_L g14309 ( 
.A(n_14206),
.B(n_2653),
.Y(n_14309)
);

INVx1_ASAP7_75t_L g14310 ( 
.A(n_14218),
.Y(n_14310)
);

AND2x4_ASAP7_75t_SL g14311 ( 
.A(n_14238),
.B(n_2653),
.Y(n_14311)
);

NAND2x1_ASAP7_75t_L g14312 ( 
.A(n_14279),
.B(n_2654),
.Y(n_14312)
);

AND2x2_ASAP7_75t_L g14313 ( 
.A(n_14207),
.B(n_2654),
.Y(n_14313)
);

AND2x4_ASAP7_75t_L g14314 ( 
.A(n_14288),
.B(n_2655),
.Y(n_14314)
);

AND2x2_ASAP7_75t_L g14315 ( 
.A(n_14204),
.B(n_14235),
.Y(n_14315)
);

OR2x2_ASAP7_75t_L g14316 ( 
.A(n_14227),
.B(n_2656),
.Y(n_14316)
);

INVx1_ASAP7_75t_L g14317 ( 
.A(n_14252),
.Y(n_14317)
);

NOR2xp33_ASAP7_75t_L g14318 ( 
.A(n_14272),
.B(n_2656),
.Y(n_14318)
);

INVx1_ASAP7_75t_SL g14319 ( 
.A(n_14187),
.Y(n_14319)
);

OR2x2_ASAP7_75t_L g14320 ( 
.A(n_14219),
.B(n_14236),
.Y(n_14320)
);

INVx1_ASAP7_75t_L g14321 ( 
.A(n_14230),
.Y(n_14321)
);

INVx1_ASAP7_75t_L g14322 ( 
.A(n_14230),
.Y(n_14322)
);

INVx1_ASAP7_75t_L g14323 ( 
.A(n_14188),
.Y(n_14323)
);

INVx1_ASAP7_75t_SL g14324 ( 
.A(n_14234),
.Y(n_14324)
);

NAND2xp5_ASAP7_75t_L g14325 ( 
.A(n_14231),
.B(n_2657),
.Y(n_14325)
);

NAND2xp5_ASAP7_75t_L g14326 ( 
.A(n_14214),
.B(n_2657),
.Y(n_14326)
);

INVx1_ASAP7_75t_L g14327 ( 
.A(n_14285),
.Y(n_14327)
);

INVx1_ASAP7_75t_L g14328 ( 
.A(n_14233),
.Y(n_14328)
);

NAND2xp5_ASAP7_75t_L g14329 ( 
.A(n_14202),
.B(n_2658),
.Y(n_14329)
);

NAND2xp5_ASAP7_75t_L g14330 ( 
.A(n_14237),
.B(n_2659),
.Y(n_14330)
);

NOR2xp33_ASAP7_75t_L g14331 ( 
.A(n_14205),
.B(n_2660),
.Y(n_14331)
);

NOR2x1_ASAP7_75t_L g14332 ( 
.A(n_14194),
.B(n_2661),
.Y(n_14332)
);

INVx1_ASAP7_75t_SL g14333 ( 
.A(n_14250),
.Y(n_14333)
);

AND2x2_ASAP7_75t_L g14334 ( 
.A(n_14223),
.B(n_2660),
.Y(n_14334)
);

NAND2xp5_ASAP7_75t_L g14335 ( 
.A(n_14276),
.B(n_14211),
.Y(n_14335)
);

NAND2xp5_ASAP7_75t_L g14336 ( 
.A(n_14191),
.B(n_2662),
.Y(n_14336)
);

NOR2x1_ASAP7_75t_L g14337 ( 
.A(n_14289),
.B(n_3360),
.Y(n_14337)
);

HB1xp67_ASAP7_75t_L g14338 ( 
.A(n_14247),
.Y(n_14338)
);

AND2x2_ASAP7_75t_L g14339 ( 
.A(n_14261),
.B(n_2662),
.Y(n_14339)
);

NOR2x1_ASAP7_75t_L g14340 ( 
.A(n_14220),
.B(n_3362),
.Y(n_14340)
);

NOR2x1_ASAP7_75t_L g14341 ( 
.A(n_14215),
.B(n_3362),
.Y(n_14341)
);

NAND2xp5_ASAP7_75t_L g14342 ( 
.A(n_14266),
.B(n_2663),
.Y(n_14342)
);

AND2x2_ASAP7_75t_L g14343 ( 
.A(n_14245),
.B(n_2663),
.Y(n_14343)
);

INVx1_ASAP7_75t_SL g14344 ( 
.A(n_14294),
.Y(n_14344)
);

NOR2xp33_ASAP7_75t_L g14345 ( 
.A(n_14260),
.B(n_14268),
.Y(n_14345)
);

HB1xp67_ASAP7_75t_L g14346 ( 
.A(n_14269),
.Y(n_14346)
);

INVx1_ASAP7_75t_L g14347 ( 
.A(n_14254),
.Y(n_14347)
);

NAND2xp5_ASAP7_75t_L g14348 ( 
.A(n_14251),
.B(n_14262),
.Y(n_14348)
);

CKINVDCx20_ASAP7_75t_R g14349 ( 
.A(n_14281),
.Y(n_14349)
);

OR2x2_ASAP7_75t_L g14350 ( 
.A(n_14256),
.B(n_2664),
.Y(n_14350)
);

HB1xp67_ASAP7_75t_L g14351 ( 
.A(n_14190),
.Y(n_14351)
);

HB1xp67_ASAP7_75t_L g14352 ( 
.A(n_14196),
.Y(n_14352)
);

NAND2xp33_ASAP7_75t_L g14353 ( 
.A(n_14244),
.B(n_2665),
.Y(n_14353)
);

NAND2xp5_ASAP7_75t_L g14354 ( 
.A(n_14199),
.B(n_2665),
.Y(n_14354)
);

INVx1_ASAP7_75t_L g14355 ( 
.A(n_14263),
.Y(n_14355)
);

INVx2_ASAP7_75t_L g14356 ( 
.A(n_14210),
.Y(n_14356)
);

INVx1_ASAP7_75t_L g14357 ( 
.A(n_14222),
.Y(n_14357)
);

INVx1_ASAP7_75t_L g14358 ( 
.A(n_14270),
.Y(n_14358)
);

NOR2xp33_ASAP7_75t_L g14359 ( 
.A(n_14226),
.B(n_2667),
.Y(n_14359)
);

OR2x2_ASAP7_75t_L g14360 ( 
.A(n_14291),
.B(n_2667),
.Y(n_14360)
);

NAND2xp5_ASAP7_75t_L g14361 ( 
.A(n_14184),
.B(n_2668),
.Y(n_14361)
);

INVx1_ASAP7_75t_L g14362 ( 
.A(n_14240),
.Y(n_14362)
);

AND2x2_ASAP7_75t_L g14363 ( 
.A(n_14292),
.B(n_2668),
.Y(n_14363)
);

NAND2xp5_ASAP7_75t_L g14364 ( 
.A(n_14264),
.B(n_14216),
.Y(n_14364)
);

OR2x2_ASAP7_75t_L g14365 ( 
.A(n_14201),
.B(n_2669),
.Y(n_14365)
);

NAND2xp5_ASAP7_75t_L g14366 ( 
.A(n_14195),
.B(n_2669),
.Y(n_14366)
);

HB1xp67_ASAP7_75t_L g14367 ( 
.A(n_14259),
.Y(n_14367)
);

INVx1_ASAP7_75t_L g14368 ( 
.A(n_14198),
.Y(n_14368)
);

NAND2xp5_ASAP7_75t_L g14369 ( 
.A(n_14229),
.B(n_2670),
.Y(n_14369)
);

INVx1_ASAP7_75t_L g14370 ( 
.A(n_14293),
.Y(n_14370)
);

INVx1_ASAP7_75t_L g14371 ( 
.A(n_14242),
.Y(n_14371)
);

AND2x2_ASAP7_75t_L g14372 ( 
.A(n_14213),
.B(n_2670),
.Y(n_14372)
);

NAND2xp5_ASAP7_75t_L g14373 ( 
.A(n_14225),
.B(n_2671),
.Y(n_14373)
);

HB1xp67_ASAP7_75t_L g14374 ( 
.A(n_14253),
.Y(n_14374)
);

INVx1_ASAP7_75t_L g14375 ( 
.A(n_14265),
.Y(n_14375)
);

HB1xp67_ASAP7_75t_L g14376 ( 
.A(n_14192),
.Y(n_14376)
);

INVx1_ASAP7_75t_L g14377 ( 
.A(n_14209),
.Y(n_14377)
);

INVxp67_ASAP7_75t_L g14378 ( 
.A(n_14287),
.Y(n_14378)
);

INVx2_ASAP7_75t_L g14379 ( 
.A(n_14232),
.Y(n_14379)
);

INVx1_ASAP7_75t_L g14380 ( 
.A(n_14273),
.Y(n_14380)
);

NOR2xp33_ASAP7_75t_L g14381 ( 
.A(n_14208),
.B(n_2671),
.Y(n_14381)
);

NAND2x1_ASAP7_75t_SL g14382 ( 
.A(n_14271),
.B(n_2672),
.Y(n_14382)
);

INVx1_ASAP7_75t_L g14383 ( 
.A(n_14282),
.Y(n_14383)
);

NAND2xp5_ASAP7_75t_L g14384 ( 
.A(n_14255),
.B(n_2672),
.Y(n_14384)
);

OR2x6_ASAP7_75t_L g14385 ( 
.A(n_14258),
.B(n_2674),
.Y(n_14385)
);

AND2x4_ASAP7_75t_SL g14386 ( 
.A(n_14284),
.B(n_2673),
.Y(n_14386)
);

INVx1_ASAP7_75t_L g14387 ( 
.A(n_14280),
.Y(n_14387)
);

INVx1_ASAP7_75t_L g14388 ( 
.A(n_14274),
.Y(n_14388)
);

INVx1_ASAP7_75t_SL g14389 ( 
.A(n_14241),
.Y(n_14389)
);

INVx1_ASAP7_75t_SL g14390 ( 
.A(n_14290),
.Y(n_14390)
);

INVxp33_ASAP7_75t_L g14391 ( 
.A(n_14359),
.Y(n_14391)
);

INVx1_ASAP7_75t_L g14392 ( 
.A(n_14300),
.Y(n_14392)
);

OR2x2_ASAP7_75t_L g14393 ( 
.A(n_14302),
.B(n_14298),
.Y(n_14393)
);

INVxp67_ASAP7_75t_L g14394 ( 
.A(n_14331),
.Y(n_14394)
);

AND2x2_ASAP7_75t_L g14395 ( 
.A(n_14334),
.B(n_14277),
.Y(n_14395)
);

HB1xp67_ASAP7_75t_L g14396 ( 
.A(n_14301),
.Y(n_14396)
);

CKINVDCx20_ASAP7_75t_R g14397 ( 
.A(n_14349),
.Y(n_14397)
);

AND2x2_ASAP7_75t_L g14398 ( 
.A(n_14363),
.B(n_14286),
.Y(n_14398)
);

INVx1_ASAP7_75t_L g14399 ( 
.A(n_14382),
.Y(n_14399)
);

INVx1_ASAP7_75t_L g14400 ( 
.A(n_14311),
.Y(n_14400)
);

INVx1_ASAP7_75t_L g14401 ( 
.A(n_14303),
.Y(n_14401)
);

AND2x2_ASAP7_75t_L g14402 ( 
.A(n_14313),
.B(n_14278),
.Y(n_14402)
);

INVx2_ASAP7_75t_L g14403 ( 
.A(n_14314),
.Y(n_14403)
);

INVx1_ASAP7_75t_L g14404 ( 
.A(n_14386),
.Y(n_14404)
);

INVx1_ASAP7_75t_L g14405 ( 
.A(n_14314),
.Y(n_14405)
);

AOI21xp5_ASAP7_75t_L g14406 ( 
.A1(n_14312),
.A2(n_14248),
.B(n_14257),
.Y(n_14406)
);

AOI21xp33_ASAP7_75t_SL g14407 ( 
.A1(n_14321),
.A2(n_14243),
.B(n_14224),
.Y(n_14407)
);

INVx1_ASAP7_75t_L g14408 ( 
.A(n_14338),
.Y(n_14408)
);

NAND2xp5_ASAP7_75t_L g14409 ( 
.A(n_14339),
.B(n_14228),
.Y(n_14409)
);

AND2x2_ASAP7_75t_L g14410 ( 
.A(n_14343),
.B(n_14275),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_14306),
.Y(n_14411)
);

INVx1_ASAP7_75t_L g14412 ( 
.A(n_14342),
.Y(n_14412)
);

A2O1A1Ixp33_ASAP7_75t_L g14413 ( 
.A1(n_14345),
.A2(n_14267),
.B(n_14283),
.C(n_2676),
.Y(n_14413)
);

INVx1_ASAP7_75t_L g14414 ( 
.A(n_14297),
.Y(n_14414)
);

INVx1_ASAP7_75t_L g14415 ( 
.A(n_14325),
.Y(n_14415)
);

NAND2xp5_ASAP7_75t_SL g14416 ( 
.A(n_14383),
.B(n_2674),
.Y(n_14416)
);

A2O1A1Ixp33_ASAP7_75t_L g14417 ( 
.A1(n_14309),
.A2(n_14318),
.B(n_14347),
.C(n_14381),
.Y(n_14417)
);

INVx1_ASAP7_75t_L g14418 ( 
.A(n_14296),
.Y(n_14418)
);

BUFx2_ASAP7_75t_L g14419 ( 
.A(n_14385),
.Y(n_14419)
);

OR2x2_ASAP7_75t_L g14420 ( 
.A(n_14385),
.B(n_14316),
.Y(n_14420)
);

AND2x2_ASAP7_75t_L g14421 ( 
.A(n_14315),
.B(n_14352),
.Y(n_14421)
);

OR2x2_ASAP7_75t_L g14422 ( 
.A(n_14373),
.B(n_2675),
.Y(n_14422)
);

OAI221xp5_ASAP7_75t_L g14423 ( 
.A1(n_14378),
.A2(n_3377),
.B1(n_2677),
.B2(n_2675),
.C(n_2676),
.Y(n_14423)
);

INVx1_ASAP7_75t_L g14424 ( 
.A(n_14351),
.Y(n_14424)
);

INVx2_ASAP7_75t_L g14425 ( 
.A(n_14372),
.Y(n_14425)
);

NOR3xp33_ASAP7_75t_SL g14426 ( 
.A(n_14348),
.B(n_2677),
.C(n_2678),
.Y(n_14426)
);

NAND2xp33_ASAP7_75t_R g14427 ( 
.A(n_14322),
.B(n_3359),
.Y(n_14427)
);

NAND2xp33_ASAP7_75t_R g14428 ( 
.A(n_14323),
.B(n_3359),
.Y(n_14428)
);

NOR2xp67_ASAP7_75t_L g14429 ( 
.A(n_14374),
.B(n_2678),
.Y(n_14429)
);

INVx1_ASAP7_75t_L g14430 ( 
.A(n_14332),
.Y(n_14430)
);

OAI21xp33_ASAP7_75t_SL g14431 ( 
.A1(n_14341),
.A2(n_2679),
.B(n_2680),
.Y(n_14431)
);

A2O1A1Ixp33_ASAP7_75t_L g14432 ( 
.A1(n_14375),
.A2(n_2683),
.B(n_2679),
.C(n_2681),
.Y(n_14432)
);

NAND2xp5_ASAP7_75t_SL g14433 ( 
.A(n_14356),
.B(n_2681),
.Y(n_14433)
);

INVx2_ASAP7_75t_L g14434 ( 
.A(n_14350),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_14353),
.Y(n_14435)
);

INVx1_ASAP7_75t_L g14436 ( 
.A(n_14308),
.Y(n_14436)
);

INVx1_ASAP7_75t_L g14437 ( 
.A(n_14336),
.Y(n_14437)
);

AND2x2_ASAP7_75t_L g14438 ( 
.A(n_14319),
.B(n_2684),
.Y(n_14438)
);

NAND2xp5_ASAP7_75t_L g14439 ( 
.A(n_14304),
.B(n_2683),
.Y(n_14439)
);

NAND2xp5_ASAP7_75t_SL g14440 ( 
.A(n_14370),
.B(n_2684),
.Y(n_14440)
);

OAI31xp33_ASAP7_75t_L g14441 ( 
.A1(n_14390),
.A2(n_2687),
.A3(n_2685),
.B(n_2686),
.Y(n_14441)
);

NAND2xp5_ASAP7_75t_L g14442 ( 
.A(n_14295),
.B(n_2685),
.Y(n_14442)
);

NOR4xp25_ASAP7_75t_SL g14443 ( 
.A(n_14357),
.B(n_3373),
.C(n_3374),
.D(n_3370),
.Y(n_14443)
);

INVx1_ASAP7_75t_L g14444 ( 
.A(n_14330),
.Y(n_14444)
);

INVx1_ASAP7_75t_L g14445 ( 
.A(n_14329),
.Y(n_14445)
);

INVx2_ASAP7_75t_L g14446 ( 
.A(n_14360),
.Y(n_14446)
);

INVx1_ASAP7_75t_L g14447 ( 
.A(n_14307),
.Y(n_14447)
);

AOI22xp5_ASAP7_75t_L g14448 ( 
.A1(n_14355),
.A2(n_2689),
.B1(n_2686),
.B2(n_2688),
.Y(n_14448)
);

INVx3_ASAP7_75t_L g14449 ( 
.A(n_14379),
.Y(n_14449)
);

NAND2xp5_ASAP7_75t_L g14450 ( 
.A(n_14317),
.B(n_2689),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_14376),
.Y(n_14451)
);

AOI21xp5_ASAP7_75t_L g14452 ( 
.A1(n_14335),
.A2(n_2690),
.B(n_2691),
.Y(n_14452)
);

NAND2xp5_ASAP7_75t_L g14453 ( 
.A(n_14337),
.B(n_2690),
.Y(n_14453)
);

NOR4xp25_ASAP7_75t_SL g14454 ( 
.A(n_14380),
.B(n_3355),
.C(n_3356),
.D(n_3354),
.Y(n_14454)
);

NAND2xp5_ASAP7_75t_L g14455 ( 
.A(n_14368),
.B(n_2691),
.Y(n_14455)
);

NAND2xp5_ASAP7_75t_L g14456 ( 
.A(n_14387),
.B(n_2692),
.Y(n_14456)
);

AOI21xp5_ASAP7_75t_L g14457 ( 
.A1(n_14326),
.A2(n_14354),
.B(n_14366),
.Y(n_14457)
);

NAND4xp25_ASAP7_75t_L g14458 ( 
.A(n_14371),
.B(n_2694),
.C(n_2692),
.D(n_2693),
.Y(n_14458)
);

NOR2xp33_ASAP7_75t_L g14459 ( 
.A(n_14365),
.B(n_2693),
.Y(n_14459)
);

NAND2xp5_ASAP7_75t_L g14460 ( 
.A(n_14324),
.B(n_14305),
.Y(n_14460)
);

AOI22xp33_ASAP7_75t_L g14461 ( 
.A1(n_14388),
.A2(n_2697),
.B1(n_2695),
.B2(n_2696),
.Y(n_14461)
);

NAND2xp5_ASAP7_75t_SL g14462 ( 
.A(n_14361),
.B(n_2695),
.Y(n_14462)
);

A2O1A1Ixp33_ASAP7_75t_L g14463 ( 
.A1(n_14340),
.A2(n_2699),
.B(n_2696),
.C(n_2698),
.Y(n_14463)
);

OAI22xp33_ASAP7_75t_L g14464 ( 
.A1(n_14384),
.A2(n_2701),
.B1(n_2699),
.B2(n_2700),
.Y(n_14464)
);

NAND2xp5_ASAP7_75t_L g14465 ( 
.A(n_14346),
.B(n_2701),
.Y(n_14465)
);

NOR3xp33_ASAP7_75t_SL g14466 ( 
.A(n_14364),
.B(n_2702),
.C(n_2703),
.Y(n_14466)
);

NAND2xp5_ASAP7_75t_L g14467 ( 
.A(n_14333),
.B(n_2702),
.Y(n_14467)
);

NOR2xp33_ASAP7_75t_L g14468 ( 
.A(n_14369),
.B(n_2704),
.Y(n_14468)
);

INVx1_ASAP7_75t_L g14469 ( 
.A(n_14438),
.Y(n_14469)
);

INVx1_ASAP7_75t_L g14470 ( 
.A(n_14456),
.Y(n_14470)
);

HB1xp67_ASAP7_75t_L g14471 ( 
.A(n_14429),
.Y(n_14471)
);

INVx1_ASAP7_75t_L g14472 ( 
.A(n_14455),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_14421),
.Y(n_14473)
);

HB1xp67_ASAP7_75t_L g14474 ( 
.A(n_14428),
.Y(n_14474)
);

NOR2xp33_ASAP7_75t_L g14475 ( 
.A(n_14431),
.B(n_14389),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_14450),
.Y(n_14476)
);

BUFx2_ASAP7_75t_L g14477 ( 
.A(n_14426),
.Y(n_14477)
);

INVx2_ASAP7_75t_L g14478 ( 
.A(n_14397),
.Y(n_14478)
);

INVx2_ASAP7_75t_L g14479 ( 
.A(n_14449),
.Y(n_14479)
);

BUFx2_ASAP7_75t_L g14480 ( 
.A(n_14466),
.Y(n_14480)
);

INVx1_ASAP7_75t_L g14481 ( 
.A(n_14465),
.Y(n_14481)
);

INVx2_ASAP7_75t_L g14482 ( 
.A(n_14449),
.Y(n_14482)
);

INVx1_ASAP7_75t_L g14483 ( 
.A(n_14442),
.Y(n_14483)
);

INVx2_ASAP7_75t_SL g14484 ( 
.A(n_14403),
.Y(n_14484)
);

INVxp33_ASAP7_75t_SL g14485 ( 
.A(n_14395),
.Y(n_14485)
);

INVxp67_ASAP7_75t_L g14486 ( 
.A(n_14427),
.Y(n_14486)
);

INVx3_ASAP7_75t_L g14487 ( 
.A(n_14399),
.Y(n_14487)
);

INVx2_ASAP7_75t_L g14488 ( 
.A(n_14422),
.Y(n_14488)
);

INVx2_ASAP7_75t_L g14489 ( 
.A(n_14392),
.Y(n_14489)
);

NOR2x1_ASAP7_75t_L g14490 ( 
.A(n_14430),
.B(n_14320),
.Y(n_14490)
);

INVx2_ASAP7_75t_L g14491 ( 
.A(n_14424),
.Y(n_14491)
);

INVx1_ASAP7_75t_L g14492 ( 
.A(n_14396),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_14439),
.Y(n_14493)
);

INVx1_ASAP7_75t_L g14494 ( 
.A(n_14453),
.Y(n_14494)
);

INVx2_ASAP7_75t_L g14495 ( 
.A(n_14405),
.Y(n_14495)
);

INVx1_ASAP7_75t_L g14496 ( 
.A(n_14467),
.Y(n_14496)
);

INVx1_ASAP7_75t_SL g14497 ( 
.A(n_14419),
.Y(n_14497)
);

INVxp33_ASAP7_75t_SL g14498 ( 
.A(n_14402),
.Y(n_14498)
);

INVx1_ASAP7_75t_L g14499 ( 
.A(n_14416),
.Y(n_14499)
);

INVx5_ASAP7_75t_L g14500 ( 
.A(n_14398),
.Y(n_14500)
);

INVx2_ASAP7_75t_SL g14501 ( 
.A(n_14433),
.Y(n_14501)
);

INVx1_ASAP7_75t_SL g14502 ( 
.A(n_14440),
.Y(n_14502)
);

INVx2_ASAP7_75t_L g14503 ( 
.A(n_14420),
.Y(n_14503)
);

INVx2_ASAP7_75t_L g14504 ( 
.A(n_14451),
.Y(n_14504)
);

INVxp67_ASAP7_75t_L g14505 ( 
.A(n_14459),
.Y(n_14505)
);

INVx2_ASAP7_75t_L g14506 ( 
.A(n_14425),
.Y(n_14506)
);

INVx1_ASAP7_75t_L g14507 ( 
.A(n_14408),
.Y(n_14507)
);

INVx5_ASAP7_75t_SL g14508 ( 
.A(n_14434),
.Y(n_14508)
);

INVx1_ASAP7_75t_L g14509 ( 
.A(n_14401),
.Y(n_14509)
);

NOR2xp33_ASAP7_75t_L g14510 ( 
.A(n_14400),
.B(n_14310),
.Y(n_14510)
);

INVx1_ASAP7_75t_L g14511 ( 
.A(n_14463),
.Y(n_14511)
);

INVx2_ASAP7_75t_L g14512 ( 
.A(n_14393),
.Y(n_14512)
);

INVx1_ASAP7_75t_L g14513 ( 
.A(n_14410),
.Y(n_14513)
);

INVx1_ASAP7_75t_L g14514 ( 
.A(n_14404),
.Y(n_14514)
);

INVx2_ASAP7_75t_L g14515 ( 
.A(n_14446),
.Y(n_14515)
);

AND2x2_ASAP7_75t_L g14516 ( 
.A(n_14454),
.B(n_14367),
.Y(n_14516)
);

CKINVDCx20_ASAP7_75t_R g14517 ( 
.A(n_14460),
.Y(n_14517)
);

NOR2xp33_ASAP7_75t_L g14518 ( 
.A(n_14391),
.B(n_14358),
.Y(n_14518)
);

NAND2xp5_ASAP7_75t_SL g14519 ( 
.A(n_14441),
.B(n_14377),
.Y(n_14519)
);

BUFx2_ASAP7_75t_L g14520 ( 
.A(n_14458),
.Y(n_14520)
);

INVx1_ASAP7_75t_L g14521 ( 
.A(n_14435),
.Y(n_14521)
);

INVx1_ASAP7_75t_L g14522 ( 
.A(n_14468),
.Y(n_14522)
);

CKINVDCx5p33_ASAP7_75t_R g14523 ( 
.A(n_14406),
.Y(n_14523)
);

INVx1_ASAP7_75t_L g14524 ( 
.A(n_14409),
.Y(n_14524)
);

INVx1_ASAP7_75t_L g14525 ( 
.A(n_14462),
.Y(n_14525)
);

INVxp67_ASAP7_75t_L g14526 ( 
.A(n_14423),
.Y(n_14526)
);

INVx2_ASAP7_75t_L g14527 ( 
.A(n_14414),
.Y(n_14527)
);

CKINVDCx20_ASAP7_75t_R g14528 ( 
.A(n_14394),
.Y(n_14528)
);

HB1xp67_ASAP7_75t_L g14529 ( 
.A(n_14432),
.Y(n_14529)
);

CKINVDCx20_ASAP7_75t_R g14530 ( 
.A(n_14411),
.Y(n_14530)
);

INVx1_ASAP7_75t_L g14531 ( 
.A(n_14464),
.Y(n_14531)
);

INVx1_ASAP7_75t_L g14532 ( 
.A(n_14452),
.Y(n_14532)
);

INVxp67_ASAP7_75t_L g14533 ( 
.A(n_14448),
.Y(n_14533)
);

INVx1_ASAP7_75t_L g14534 ( 
.A(n_14418),
.Y(n_14534)
);

INVx1_ASAP7_75t_L g14535 ( 
.A(n_14413),
.Y(n_14535)
);

INVx2_ASAP7_75t_L g14536 ( 
.A(n_14412),
.Y(n_14536)
);

INVx1_ASAP7_75t_L g14537 ( 
.A(n_14415),
.Y(n_14537)
);

INVx2_ASAP7_75t_L g14538 ( 
.A(n_14447),
.Y(n_14538)
);

INVx1_ASAP7_75t_L g14539 ( 
.A(n_14436),
.Y(n_14539)
);

INVx2_ASAP7_75t_L g14540 ( 
.A(n_14444),
.Y(n_14540)
);

CKINVDCx6p67_ASAP7_75t_R g14541 ( 
.A(n_14445),
.Y(n_14541)
);

INVx2_ASAP7_75t_SL g14542 ( 
.A(n_14437),
.Y(n_14542)
);

INVx2_ASAP7_75t_SL g14543 ( 
.A(n_14443),
.Y(n_14543)
);

BUFx2_ASAP7_75t_L g14544 ( 
.A(n_14417),
.Y(n_14544)
);

INVx2_ASAP7_75t_L g14545 ( 
.A(n_14461),
.Y(n_14545)
);

HB1xp67_ASAP7_75t_L g14546 ( 
.A(n_14457),
.Y(n_14546)
);

INVx2_ASAP7_75t_L g14547 ( 
.A(n_14407),
.Y(n_14547)
);

INVx1_ASAP7_75t_L g14548 ( 
.A(n_14438),
.Y(n_14548)
);

INVxp33_ASAP7_75t_L g14549 ( 
.A(n_14438),
.Y(n_14549)
);

INVx2_ASAP7_75t_L g14550 ( 
.A(n_14478),
.Y(n_14550)
);

AOI221xp5_ASAP7_75t_L g14551 ( 
.A1(n_14473),
.A2(n_14344),
.B1(n_14327),
.B2(n_14328),
.C(n_14362),
.Y(n_14551)
);

AOI22xp5_ASAP7_75t_L g14552 ( 
.A1(n_14517),
.A2(n_14299),
.B1(n_2707),
.B2(n_2705),
.Y(n_14552)
);

INVx1_ASAP7_75t_L g14553 ( 
.A(n_14516),
.Y(n_14553)
);

INVxp67_ASAP7_75t_L g14554 ( 
.A(n_14471),
.Y(n_14554)
);

AOI22xp5_ASAP7_75t_L g14555 ( 
.A1(n_14498),
.A2(n_2707),
.B1(n_2705),
.B2(n_2706),
.Y(n_14555)
);

INVx2_ASAP7_75t_L g14556 ( 
.A(n_14500),
.Y(n_14556)
);

AOI22xp5_ASAP7_75t_L g14557 ( 
.A1(n_14485),
.A2(n_2709),
.B1(n_2706),
.B2(n_2708),
.Y(n_14557)
);

AOI31xp33_ASAP7_75t_L g14558 ( 
.A1(n_14543),
.A2(n_2711),
.A3(n_2708),
.B(n_2710),
.Y(n_14558)
);

OA22x2_ASAP7_75t_L g14559 ( 
.A1(n_14497),
.A2(n_2713),
.B1(n_2711),
.B2(n_2712),
.Y(n_14559)
);

INVx1_ASAP7_75t_L g14560 ( 
.A(n_14495),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_14474),
.Y(n_14561)
);

INVx1_ASAP7_75t_L g14562 ( 
.A(n_14500),
.Y(n_14562)
);

O2A1O1Ixp33_ASAP7_75t_SL g14563 ( 
.A1(n_14486),
.A2(n_14519),
.B(n_14492),
.C(n_14507),
.Y(n_14563)
);

INVx1_ASAP7_75t_L g14564 ( 
.A(n_14484),
.Y(n_14564)
);

INVx1_ASAP7_75t_L g14565 ( 
.A(n_14479),
.Y(n_14565)
);

OAI221xp5_ASAP7_75t_SL g14566 ( 
.A1(n_14489),
.A2(n_3366),
.B1(n_3367),
.B2(n_3365),
.C(n_3364),
.Y(n_14566)
);

AOI22xp5_ASAP7_75t_L g14567 ( 
.A1(n_14523),
.A2(n_2717),
.B1(n_2715),
.B2(n_2716),
.Y(n_14567)
);

AOI221xp5_ASAP7_75t_L g14568 ( 
.A1(n_14514),
.A2(n_2717),
.B1(n_2715),
.B2(n_2716),
.C(n_2718),
.Y(n_14568)
);

AOI221xp5_ASAP7_75t_L g14569 ( 
.A1(n_14475),
.A2(n_2720),
.B1(n_2718),
.B2(n_2719),
.C(n_2721),
.Y(n_14569)
);

INVx1_ASAP7_75t_L g14570 ( 
.A(n_14482),
.Y(n_14570)
);

INVx1_ASAP7_75t_L g14571 ( 
.A(n_14477),
.Y(n_14571)
);

AOI22xp5_ASAP7_75t_L g14572 ( 
.A1(n_14528),
.A2(n_2721),
.B1(n_2719),
.B2(n_2720),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_14480),
.Y(n_14573)
);

INVx1_ASAP7_75t_L g14574 ( 
.A(n_14491),
.Y(n_14574)
);

INVx1_ASAP7_75t_L g14575 ( 
.A(n_14504),
.Y(n_14575)
);

INVx1_ASAP7_75t_L g14576 ( 
.A(n_14490),
.Y(n_14576)
);

INVx2_ASAP7_75t_L g14577 ( 
.A(n_14547),
.Y(n_14577)
);

INVx1_ASAP7_75t_SL g14578 ( 
.A(n_14502),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_14509),
.Y(n_14579)
);

AOI22xp5_ASAP7_75t_L g14580 ( 
.A1(n_14530),
.A2(n_2724),
.B1(n_2722),
.B2(n_2723),
.Y(n_14580)
);

INVxp67_ASAP7_75t_L g14581 ( 
.A(n_14510),
.Y(n_14581)
);

OAI22xp5_ASAP7_75t_L g14582 ( 
.A1(n_14513),
.A2(n_2724),
.B1(n_2722),
.B2(n_2723),
.Y(n_14582)
);

AOI22xp5_ASAP7_75t_L g14583 ( 
.A1(n_14521),
.A2(n_2727),
.B1(n_2725),
.B2(n_2726),
.Y(n_14583)
);

OAI22x1_ASAP7_75t_L g14584 ( 
.A1(n_14515),
.A2(n_2735),
.B1(n_2744),
.B2(n_2726),
.Y(n_14584)
);

CKINVDCx5p33_ASAP7_75t_R g14585 ( 
.A(n_14541),
.Y(n_14585)
);

HB1xp67_ASAP7_75t_L g14586 ( 
.A(n_14503),
.Y(n_14586)
);

A2O1A1Ixp33_ASAP7_75t_SL g14587 ( 
.A1(n_14487),
.A2(n_2730),
.B(n_2728),
.C(n_2729),
.Y(n_14587)
);

AOI31xp33_ASAP7_75t_L g14588 ( 
.A1(n_14549),
.A2(n_2732),
.A3(n_2729),
.B(n_2731),
.Y(n_14588)
);

O2A1O1Ixp33_ASAP7_75t_SL g14589 ( 
.A1(n_14501),
.A2(n_2733),
.B(n_2731),
.C(n_2732),
.Y(n_14589)
);

OAI22x1_ASAP7_75t_L g14590 ( 
.A1(n_14506),
.A2(n_2742),
.B1(n_2751),
.B2(n_2734),
.Y(n_14590)
);

INVx1_ASAP7_75t_L g14591 ( 
.A(n_14529),
.Y(n_14591)
);

OAI22xp5_ASAP7_75t_L g14592 ( 
.A1(n_14508),
.A2(n_2737),
.B1(n_2735),
.B2(n_2736),
.Y(n_14592)
);

AOI22xp5_ASAP7_75t_L g14593 ( 
.A1(n_14518),
.A2(n_2739),
.B1(n_2736),
.B2(n_2738),
.Y(n_14593)
);

AND4x1_ASAP7_75t_L g14594 ( 
.A(n_14469),
.B(n_2740),
.C(n_2738),
.D(n_2739),
.Y(n_14594)
);

AOI22x1_ASAP7_75t_SL g14595 ( 
.A1(n_14548),
.A2(n_2744),
.B1(n_2741),
.B2(n_2742),
.Y(n_14595)
);

OA22x2_ASAP7_75t_L g14596 ( 
.A1(n_14511),
.A2(n_2747),
.B1(n_2745),
.B2(n_2746),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_14544),
.Y(n_14597)
);

NAND2xp5_ASAP7_75t_L g14598 ( 
.A(n_14508),
.B(n_2745),
.Y(n_14598)
);

INVx1_ASAP7_75t_L g14599 ( 
.A(n_14520),
.Y(n_14599)
);

INVx1_ASAP7_75t_L g14600 ( 
.A(n_14546),
.Y(n_14600)
);

AOI31xp33_ASAP7_75t_L g14601 ( 
.A1(n_14499),
.A2(n_2749),
.A3(n_2746),
.B(n_2748),
.Y(n_14601)
);

INVx2_ASAP7_75t_L g14602 ( 
.A(n_14488),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_14512),
.Y(n_14603)
);

INVx2_ASAP7_75t_L g14604 ( 
.A(n_14493),
.Y(n_14604)
);

INVx1_ASAP7_75t_L g14605 ( 
.A(n_14524),
.Y(n_14605)
);

OAI22xp5_ASAP7_75t_L g14606 ( 
.A1(n_14533),
.A2(n_2750),
.B1(n_2748),
.B2(n_2749),
.Y(n_14606)
);

AOI22xp5_ASAP7_75t_L g14607 ( 
.A1(n_14542),
.A2(n_2753),
.B1(n_2750),
.B2(n_2752),
.Y(n_14607)
);

INVx2_ASAP7_75t_L g14608 ( 
.A(n_14496),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_14534),
.Y(n_14609)
);

INVx1_ASAP7_75t_L g14610 ( 
.A(n_14527),
.Y(n_14610)
);

INVx2_ASAP7_75t_L g14611 ( 
.A(n_14545),
.Y(n_14611)
);

INVxp67_ASAP7_75t_L g14612 ( 
.A(n_14537),
.Y(n_14612)
);

AOI22xp5_ASAP7_75t_L g14613 ( 
.A1(n_14539),
.A2(n_2755),
.B1(n_2752),
.B2(n_2754),
.Y(n_14613)
);

OAI211xp5_ASAP7_75t_SL g14614 ( 
.A1(n_14551),
.A2(n_14526),
.B(n_14531),
.C(n_14505),
.Y(n_14614)
);

AOI221xp5_ASAP7_75t_L g14615 ( 
.A1(n_14563),
.A2(n_14535),
.B1(n_14532),
.B2(n_14525),
.C(n_14538),
.Y(n_14615)
);

INVx1_ASAP7_75t_L g14616 ( 
.A(n_14598),
.Y(n_14616)
);

NOR3xp33_ASAP7_75t_L g14617 ( 
.A(n_14576),
.B(n_14536),
.C(n_14540),
.Y(n_14617)
);

AND2x2_ASAP7_75t_L g14618 ( 
.A(n_14586),
.B(n_14494),
.Y(n_14618)
);

AOI211x1_ASAP7_75t_SL g14619 ( 
.A1(n_14556),
.A2(n_14481),
.B(n_14483),
.C(n_14476),
.Y(n_14619)
);

NAND2xp5_ASAP7_75t_L g14620 ( 
.A(n_14558),
.B(n_14472),
.Y(n_14620)
);

INVx1_ASAP7_75t_L g14621 ( 
.A(n_14559),
.Y(n_14621)
);

AO22x2_ASAP7_75t_L g14622 ( 
.A1(n_14553),
.A2(n_14470),
.B1(n_14522),
.B2(n_2756),
.Y(n_14622)
);

AOI221xp5_ASAP7_75t_L g14623 ( 
.A1(n_14562),
.A2(n_2756),
.B1(n_2754),
.B2(n_2755),
.C(n_2757),
.Y(n_14623)
);

OAI211xp5_ASAP7_75t_SL g14624 ( 
.A1(n_14581),
.A2(n_2759),
.B(n_2757),
.C(n_2758),
.Y(n_14624)
);

AOI221xp5_ASAP7_75t_L g14625 ( 
.A1(n_14564),
.A2(n_2761),
.B1(n_2758),
.B2(n_2760),
.C(n_2762),
.Y(n_14625)
);

NAND2xp5_ASAP7_75t_L g14626 ( 
.A(n_14552),
.B(n_3360),
.Y(n_14626)
);

A2O1A1Ixp33_ASAP7_75t_L g14627 ( 
.A1(n_14560),
.A2(n_2764),
.B(n_2760),
.C(n_2763),
.Y(n_14627)
);

CKINVDCx5p33_ASAP7_75t_R g14628 ( 
.A(n_14585),
.Y(n_14628)
);

AOI221xp5_ASAP7_75t_L g14629 ( 
.A1(n_14597),
.A2(n_2766),
.B1(n_2763),
.B2(n_2765),
.C(n_2767),
.Y(n_14629)
);

NAND4xp25_ASAP7_75t_L g14630 ( 
.A(n_14603),
.B(n_2767),
.C(n_2765),
.D(n_2766),
.Y(n_14630)
);

NAND4xp25_ASAP7_75t_SL g14631 ( 
.A(n_14578),
.B(n_2770),
.C(n_2768),
.D(n_2769),
.Y(n_14631)
);

NAND5xp2_ASAP7_75t_L g14632 ( 
.A(n_14574),
.B(n_3353),
.C(n_3354),
.D(n_3352),
.E(n_3351),
.Y(n_14632)
);

AOI21xp33_ASAP7_75t_SL g14633 ( 
.A1(n_14596),
.A2(n_2768),
.B(n_2771),
.Y(n_14633)
);

AOI221xp5_ASAP7_75t_L g14634 ( 
.A1(n_14554),
.A2(n_2773),
.B1(n_2771),
.B2(n_2772),
.C(n_2774),
.Y(n_14634)
);

AOI222xp33_ASAP7_75t_L g14635 ( 
.A1(n_14612),
.A2(n_2796),
.B1(n_2780),
.B2(n_2804),
.C1(n_2788),
.C2(n_2772),
.Y(n_14635)
);

OAI21xp33_ASAP7_75t_SL g14636 ( 
.A1(n_14575),
.A2(n_2773),
.B(n_2774),
.Y(n_14636)
);

INVx2_ASAP7_75t_L g14637 ( 
.A(n_14590),
.Y(n_14637)
);

NOR4xp25_ASAP7_75t_L g14638 ( 
.A(n_14579),
.B(n_2777),
.C(n_2775),
.D(n_2776),
.Y(n_14638)
);

AOI211xp5_ASAP7_75t_L g14639 ( 
.A1(n_14610),
.A2(n_2777),
.B(n_2775),
.C(n_2776),
.Y(n_14639)
);

OAI211xp5_ASAP7_75t_SL g14640 ( 
.A1(n_14609),
.A2(n_2781),
.B(n_2778),
.C(n_2779),
.Y(n_14640)
);

AOI211xp5_ASAP7_75t_L g14641 ( 
.A1(n_14565),
.A2(n_2783),
.B(n_2779),
.C(n_2782),
.Y(n_14641)
);

AOI221xp5_ASAP7_75t_L g14642 ( 
.A1(n_14571),
.A2(n_2784),
.B1(n_2782),
.B2(n_2783),
.C(n_2785),
.Y(n_14642)
);

OAI321xp33_ASAP7_75t_L g14643 ( 
.A1(n_14573),
.A2(n_2787),
.A3(n_2790),
.B1(n_2784),
.B2(n_2786),
.C(n_2789),
.Y(n_14643)
);

AOI221xp5_ASAP7_75t_L g14644 ( 
.A1(n_14591),
.A2(n_2790),
.B1(n_2787),
.B2(n_2789),
.C(n_2791),
.Y(n_14644)
);

NAND4xp25_ASAP7_75t_L g14645 ( 
.A(n_14561),
.B(n_2794),
.C(n_2792),
.D(n_2793),
.Y(n_14645)
);

AOI222xp33_ASAP7_75t_L g14646 ( 
.A1(n_14570),
.A2(n_2820),
.B1(n_2802),
.B2(n_2828),
.C1(n_2811),
.C2(n_2792),
.Y(n_14646)
);

AOI211xp5_ASAP7_75t_L g14647 ( 
.A1(n_14587),
.A2(n_2797),
.B(n_2793),
.C(n_2795),
.Y(n_14647)
);

O2A1O1Ixp5_ASAP7_75t_L g14648 ( 
.A1(n_14550),
.A2(n_3375),
.B(n_3377),
.C(n_3373),
.Y(n_14648)
);

O2A1O1Ixp5_ASAP7_75t_SL g14649 ( 
.A1(n_14600),
.A2(n_2798),
.B(n_2795),
.C(n_2797),
.Y(n_14649)
);

AOI211xp5_ASAP7_75t_L g14650 ( 
.A1(n_14605),
.A2(n_2800),
.B(n_2798),
.C(n_2799),
.Y(n_14650)
);

OAI221xp5_ASAP7_75t_SL g14651 ( 
.A1(n_14577),
.A2(n_2801),
.B1(n_2803),
.B2(n_2800),
.C(n_2802),
.Y(n_14651)
);

AND2x2_ASAP7_75t_L g14652 ( 
.A(n_14602),
.B(n_2799),
.Y(n_14652)
);

OAI21xp5_ASAP7_75t_SL g14653 ( 
.A1(n_14599),
.A2(n_2804),
.B(n_2803),
.Y(n_14653)
);

NAND2xp5_ASAP7_75t_L g14654 ( 
.A(n_14594),
.B(n_3355),
.Y(n_14654)
);

NOR2xp33_ASAP7_75t_R g14655 ( 
.A(n_14611),
.B(n_2801),
.Y(n_14655)
);

AOI222xp33_ASAP7_75t_L g14656 ( 
.A1(n_14604),
.A2(n_2831),
.B1(n_2814),
.B2(n_2840),
.C1(n_2823),
.C2(n_2805),
.Y(n_14656)
);

INVx1_ASAP7_75t_L g14657 ( 
.A(n_14595),
.Y(n_14657)
);

OAI22xp33_ASAP7_75t_SL g14658 ( 
.A1(n_14608),
.A2(n_2808),
.B1(n_2806),
.B2(n_2807),
.Y(n_14658)
);

AOI22xp5_ASAP7_75t_L g14659 ( 
.A1(n_14569),
.A2(n_2808),
.B1(n_2806),
.B2(n_2807),
.Y(n_14659)
);

AOI322xp5_ASAP7_75t_L g14660 ( 
.A1(n_14567),
.A2(n_2815),
.A3(n_2814),
.B1(n_2812),
.B2(n_2809),
.C1(n_2811),
.C2(n_2813),
.Y(n_14660)
);

A2O1A1Ixp33_ASAP7_75t_L g14661 ( 
.A1(n_14568),
.A2(n_2815),
.B(n_2809),
.C(n_2813),
.Y(n_14661)
);

NOR2x1_ASAP7_75t_SL g14662 ( 
.A(n_14582),
.B(n_2817),
.Y(n_14662)
);

OAI222xp33_ASAP7_75t_L g14663 ( 
.A1(n_14566),
.A2(n_2818),
.B1(n_2821),
.B2(n_2816),
.C1(n_2817),
.C2(n_2820),
.Y(n_14663)
);

AOI221xp5_ASAP7_75t_L g14664 ( 
.A1(n_14589),
.A2(n_2822),
.B1(n_2816),
.B2(n_2818),
.C(n_2824),
.Y(n_14664)
);

AOI22xp33_ASAP7_75t_L g14665 ( 
.A1(n_14584),
.A2(n_2825),
.B1(n_2822),
.B2(n_2824),
.Y(n_14665)
);

INVx1_ASAP7_75t_L g14666 ( 
.A(n_14588),
.Y(n_14666)
);

NOR2xp67_ASAP7_75t_L g14667 ( 
.A(n_14593),
.B(n_2826),
.Y(n_14667)
);

AOI21xp5_ASAP7_75t_L g14668 ( 
.A1(n_14601),
.A2(n_14606),
.B(n_14592),
.Y(n_14668)
);

OAI22xp33_ASAP7_75t_L g14669 ( 
.A1(n_14607),
.A2(n_2829),
.B1(n_2827),
.B2(n_2828),
.Y(n_14669)
);

AOI211xp5_ASAP7_75t_L g14670 ( 
.A1(n_14580),
.A2(n_2831),
.B(n_2827),
.C(n_2830),
.Y(n_14670)
);

OAI221xp5_ASAP7_75t_L g14671 ( 
.A1(n_14555),
.A2(n_2833),
.B1(n_2830),
.B2(n_2832),
.C(n_2834),
.Y(n_14671)
);

NAND2xp5_ASAP7_75t_L g14672 ( 
.A(n_14557),
.B(n_3351),
.Y(n_14672)
);

NOR4xp25_ASAP7_75t_L g14673 ( 
.A(n_14613),
.B(n_2837),
.C(n_2835),
.D(n_2836),
.Y(n_14673)
);

NAND4xp75_ASAP7_75t_L g14674 ( 
.A(n_14572),
.B(n_2839),
.C(n_2836),
.D(n_2837),
.Y(n_14674)
);

OAI211xp5_ASAP7_75t_L g14675 ( 
.A1(n_14583),
.A2(n_2843),
.B(n_2841),
.C(n_2842),
.Y(n_14675)
);

AOI221xp5_ASAP7_75t_L g14676 ( 
.A1(n_14563),
.A2(n_2845),
.B1(n_2842),
.B2(n_2844),
.C(n_2846),
.Y(n_14676)
);

NOR4xp25_ASAP7_75t_SL g14677 ( 
.A(n_14585),
.B(n_2846),
.C(n_2844),
.D(n_2845),
.Y(n_14677)
);

OAI221xp5_ASAP7_75t_L g14678 ( 
.A1(n_14587),
.A2(n_2849),
.B1(n_2847),
.B2(n_2848),
.C(n_2850),
.Y(n_14678)
);

AOI222xp33_ASAP7_75t_L g14679 ( 
.A1(n_14576),
.A2(n_2873),
.B1(n_2856),
.B2(n_2881),
.C1(n_2864),
.C2(n_2847),
.Y(n_14679)
);

AOI21xp5_ASAP7_75t_L g14680 ( 
.A1(n_14563),
.A2(n_2849),
.B(n_2850),
.Y(n_14680)
);

INVx1_ASAP7_75t_L g14681 ( 
.A(n_14598),
.Y(n_14681)
);

OAI211xp5_ASAP7_75t_SL g14682 ( 
.A1(n_14551),
.A2(n_2853),
.B(n_2851),
.C(n_2852),
.Y(n_14682)
);

INVx1_ASAP7_75t_L g14683 ( 
.A(n_14622),
.Y(n_14683)
);

NOR3xp33_ASAP7_75t_L g14684 ( 
.A(n_14614),
.B(n_2854),
.C(n_2855),
.Y(n_14684)
);

NOR4xp25_ASAP7_75t_L g14685 ( 
.A(n_14615),
.B(n_3365),
.C(n_2857),
.D(n_2855),
.Y(n_14685)
);

NOR4xp75_ASAP7_75t_L g14686 ( 
.A(n_14620),
.B(n_2858),
.C(n_2856),
.D(n_2857),
.Y(n_14686)
);

NAND2xp5_ASAP7_75t_L g14687 ( 
.A(n_14676),
.B(n_2859),
.Y(n_14687)
);

AO21x1_ASAP7_75t_L g14688 ( 
.A1(n_14680),
.A2(n_2858),
.B(n_2859),
.Y(n_14688)
);

OAI221xp5_ASAP7_75t_L g14689 ( 
.A1(n_14636),
.A2(n_2862),
.B1(n_2860),
.B2(n_2861),
.C(n_2863),
.Y(n_14689)
);

NOR3x1_ASAP7_75t_L g14690 ( 
.A(n_14674),
.B(n_2860),
.C(n_2861),
.Y(n_14690)
);

INVx1_ASAP7_75t_L g14691 ( 
.A(n_14622),
.Y(n_14691)
);

INVx1_ASAP7_75t_L g14692 ( 
.A(n_14654),
.Y(n_14692)
);

O2A1O1Ixp5_ASAP7_75t_L g14693 ( 
.A1(n_14637),
.A2(n_2865),
.B(n_2862),
.C(n_2863),
.Y(n_14693)
);

OA211x2_ASAP7_75t_L g14694 ( 
.A1(n_14664),
.A2(n_2867),
.B(n_2865),
.C(n_2866),
.Y(n_14694)
);

AND4x1_ASAP7_75t_L g14695 ( 
.A(n_14619),
.B(n_2869),
.C(n_2866),
.D(n_2868),
.Y(n_14695)
);

NAND4xp25_ASAP7_75t_SL g14696 ( 
.A(n_14647),
.B(n_2870),
.C(n_2868),
.D(n_2869),
.Y(n_14696)
);

NOR2x1_ASAP7_75t_L g14697 ( 
.A(n_14631),
.B(n_14657),
.Y(n_14697)
);

OR2x2_ASAP7_75t_L g14698 ( 
.A(n_14638),
.B(n_2872),
.Y(n_14698)
);

AND4x2_ASAP7_75t_L g14699 ( 
.A(n_14668),
.B(n_2876),
.C(n_2874),
.D(n_2875),
.Y(n_14699)
);

NOR2xp67_ASAP7_75t_L g14700 ( 
.A(n_14632),
.B(n_2875),
.Y(n_14700)
);

OAI221xp5_ASAP7_75t_L g14701 ( 
.A1(n_14665),
.A2(n_2877),
.B1(n_2874),
.B2(n_2876),
.C(n_2878),
.Y(n_14701)
);

AOI221xp5_ASAP7_75t_L g14702 ( 
.A1(n_14633),
.A2(n_2879),
.B1(n_2877),
.B2(n_2878),
.C(n_2880),
.Y(n_14702)
);

AND4x1_ASAP7_75t_L g14703 ( 
.A(n_14617),
.B(n_2882),
.C(n_2879),
.D(n_2880),
.Y(n_14703)
);

NOR3xp33_ASAP7_75t_L g14704 ( 
.A(n_14618),
.B(n_2882),
.C(n_2883),
.Y(n_14704)
);

AOI211xp5_ASAP7_75t_L g14705 ( 
.A1(n_14669),
.A2(n_2885),
.B(n_2883),
.C(n_2884),
.Y(n_14705)
);

NAND2xp5_ASAP7_75t_SL g14706 ( 
.A(n_14628),
.B(n_2884),
.Y(n_14706)
);

NAND3xp33_ASAP7_75t_SL g14707 ( 
.A(n_14677),
.B(n_2885),
.C(n_2886),
.Y(n_14707)
);

NOR3xp33_ASAP7_75t_L g14708 ( 
.A(n_14666),
.B(n_2887),
.C(n_2888),
.Y(n_14708)
);

AOI211xp5_ASAP7_75t_L g14709 ( 
.A1(n_14663),
.A2(n_2890),
.B(n_2887),
.C(n_2889),
.Y(n_14709)
);

OAI321xp33_ASAP7_75t_L g14710 ( 
.A1(n_14621),
.A2(n_2893),
.A3(n_2896),
.B1(n_2891),
.B2(n_2892),
.C(n_2895),
.Y(n_14710)
);

NOR3xp33_ASAP7_75t_SL g14711 ( 
.A(n_14682),
.B(n_2891),
.C(n_2895),
.Y(n_14711)
);

AOI21xp5_ASAP7_75t_L g14712 ( 
.A1(n_14672),
.A2(n_14662),
.B(n_14626),
.Y(n_14712)
);

AOI21xp5_ASAP7_75t_L g14713 ( 
.A1(n_14667),
.A2(n_2896),
.B(n_2897),
.Y(n_14713)
);

NAND4xp25_ASAP7_75t_SL g14714 ( 
.A(n_14649),
.B(n_2899),
.C(n_2897),
.D(n_2898),
.Y(n_14714)
);

NOR2xp33_ASAP7_75t_L g14715 ( 
.A(n_14678),
.B(n_3348),
.Y(n_14715)
);

NAND5xp2_ASAP7_75t_L g14716 ( 
.A(n_14616),
.B(n_2901),
.C(n_2898),
.D(n_2900),
.E(n_2902),
.Y(n_14716)
);

NAND2xp5_ASAP7_75t_SL g14717 ( 
.A(n_14673),
.B(n_2900),
.Y(n_14717)
);

NAND5xp2_ASAP7_75t_L g14718 ( 
.A(n_14681),
.B(n_2903),
.C(n_2901),
.D(n_2902),
.E(n_2904),
.Y(n_14718)
);

OAI22xp5_ASAP7_75t_SL g14719 ( 
.A1(n_14671),
.A2(n_2905),
.B1(n_2903),
.B2(n_2904),
.Y(n_14719)
);

NAND2xp5_ASAP7_75t_SL g14720 ( 
.A(n_14670),
.B(n_2905),
.Y(n_14720)
);

NOR3xp33_ASAP7_75t_L g14721 ( 
.A(n_14675),
.B(n_2906),
.C(n_2907),
.Y(n_14721)
);

OAI211xp5_ASAP7_75t_L g14722 ( 
.A1(n_14653),
.A2(n_2910),
.B(n_2911),
.C(n_2909),
.Y(n_14722)
);

OAI21xp33_ASAP7_75t_L g14723 ( 
.A1(n_14659),
.A2(n_2908),
.B(n_2910),
.Y(n_14723)
);

INVx1_ASAP7_75t_L g14724 ( 
.A(n_14655),
.Y(n_14724)
);

OAI211xp5_ASAP7_75t_SL g14725 ( 
.A1(n_14661),
.A2(n_2912),
.B(n_2908),
.C(n_2911),
.Y(n_14725)
);

NOR3xp33_ASAP7_75t_L g14726 ( 
.A(n_14624),
.B(n_2912),
.C(n_2913),
.Y(n_14726)
);

NAND2xp5_ASAP7_75t_L g14727 ( 
.A(n_14650),
.B(n_2914),
.Y(n_14727)
);

AOI221xp5_ASAP7_75t_L g14728 ( 
.A1(n_14648),
.A2(n_2916),
.B1(n_2913),
.B2(n_2915),
.C(n_2917),
.Y(n_14728)
);

NAND4xp25_ASAP7_75t_L g14729 ( 
.A(n_14639),
.B(n_2918),
.C(n_2915),
.D(n_2916),
.Y(n_14729)
);

NOR3xp33_ASAP7_75t_L g14730 ( 
.A(n_14640),
.B(n_2918),
.C(n_2919),
.Y(n_14730)
);

NAND2xp5_ASAP7_75t_SL g14731 ( 
.A(n_14658),
.B(n_2919),
.Y(n_14731)
);

NAND3xp33_ASAP7_75t_SL g14732 ( 
.A(n_14641),
.B(n_2920),
.C(n_2921),
.Y(n_14732)
);

OR2x2_ASAP7_75t_L g14733 ( 
.A(n_14630),
.B(n_2920),
.Y(n_14733)
);

OAI221xp5_ASAP7_75t_L g14734 ( 
.A1(n_14629),
.A2(n_14634),
.B1(n_14644),
.B2(n_14625),
.C(n_14642),
.Y(n_14734)
);

AOI211xp5_ASAP7_75t_L g14735 ( 
.A1(n_14651),
.A2(n_14645),
.B(n_14643),
.C(n_14627),
.Y(n_14735)
);

OA21x2_ASAP7_75t_L g14736 ( 
.A1(n_14623),
.A2(n_2921),
.B(n_2922),
.Y(n_14736)
);

A2O1A1Ixp33_ASAP7_75t_L g14737 ( 
.A1(n_14660),
.A2(n_14652),
.B(n_14679),
.C(n_14656),
.Y(n_14737)
);

NOR2x1_ASAP7_75t_L g14738 ( 
.A(n_14635),
.B(n_2923),
.Y(n_14738)
);

NAND3xp33_ASAP7_75t_SL g14739 ( 
.A(n_14646),
.B(n_2922),
.C(n_2923),
.Y(n_14739)
);

INVx3_ASAP7_75t_SL g14740 ( 
.A(n_14628),
.Y(n_14740)
);

HB1xp67_ASAP7_75t_L g14741 ( 
.A(n_14655),
.Y(n_14741)
);

NAND4xp25_ASAP7_75t_L g14742 ( 
.A(n_14615),
.B(n_2926),
.C(n_2924),
.D(n_2925),
.Y(n_14742)
);

INVx3_ASAP7_75t_L g14743 ( 
.A(n_14674),
.Y(n_14743)
);

AOI21xp5_ASAP7_75t_L g14744 ( 
.A1(n_14654),
.A2(n_2924),
.B(n_2925),
.Y(n_14744)
);

NOR2x1_ASAP7_75t_L g14745 ( 
.A(n_14631),
.B(n_2927),
.Y(n_14745)
);

NAND3xp33_ASAP7_75t_SL g14746 ( 
.A(n_14628),
.B(n_2926),
.C(n_2927),
.Y(n_14746)
);

NAND4xp25_ASAP7_75t_L g14747 ( 
.A(n_14615),
.B(n_2931),
.C(n_2928),
.D(n_2929),
.Y(n_14747)
);

INVxp33_ASAP7_75t_SL g14748 ( 
.A(n_14628),
.Y(n_14748)
);

NAND4xp75_ASAP7_75t_L g14749 ( 
.A(n_14615),
.B(n_2932),
.C(n_2928),
.D(n_2929),
.Y(n_14749)
);

NOR3x1_ASAP7_75t_L g14750 ( 
.A(n_14674),
.B(n_2932),
.C(n_2933),
.Y(n_14750)
);

OAI211xp5_ASAP7_75t_L g14751 ( 
.A1(n_14676),
.A2(n_2935),
.B(n_2936),
.C(n_2934),
.Y(n_14751)
);

NAND2xp5_ASAP7_75t_SL g14752 ( 
.A(n_14676),
.B(n_2933),
.Y(n_14752)
);

NOR2x1_ASAP7_75t_L g14753 ( 
.A(n_14631),
.B(n_2936),
.Y(n_14753)
);

NAND2xp5_ASAP7_75t_L g14754 ( 
.A(n_14676),
.B(n_2937),
.Y(n_14754)
);

NAND2xp5_ASAP7_75t_L g14755 ( 
.A(n_14676),
.B(n_2937),
.Y(n_14755)
);

NAND5xp2_ASAP7_75t_L g14756 ( 
.A(n_14615),
.B(n_2939),
.C(n_2935),
.D(n_2938),
.E(n_2940),
.Y(n_14756)
);

AOI21xp5_ASAP7_75t_L g14757 ( 
.A1(n_14654),
.A2(n_2938),
.B(n_2939),
.Y(n_14757)
);

BUFx8_ASAP7_75t_SL g14758 ( 
.A(n_14743),
.Y(n_14758)
);

HB1xp67_ASAP7_75t_L g14759 ( 
.A(n_14686),
.Y(n_14759)
);

NAND2xp33_ASAP7_75t_L g14760 ( 
.A(n_14704),
.B(n_2940),
.Y(n_14760)
);

CKINVDCx20_ASAP7_75t_R g14761 ( 
.A(n_14740),
.Y(n_14761)
);

AOI22xp5_ASAP7_75t_L g14762 ( 
.A1(n_14748),
.A2(n_2943),
.B1(n_2941),
.B2(n_2942),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_14699),
.Y(n_14763)
);

AOI21xp5_ASAP7_75t_L g14764 ( 
.A1(n_14717),
.A2(n_2941),
.B(n_2942),
.Y(n_14764)
);

INVx1_ASAP7_75t_SL g14765 ( 
.A(n_14698),
.Y(n_14765)
);

NAND2xp33_ASAP7_75t_R g14766 ( 
.A(n_14743),
.B(n_2944),
.Y(n_14766)
);

OAI21x1_ASAP7_75t_SL g14767 ( 
.A1(n_14688),
.A2(n_3375),
.B(n_2943),
.Y(n_14767)
);

XOR2xp5_ASAP7_75t_L g14768 ( 
.A(n_14749),
.B(n_2944),
.Y(n_14768)
);

NOR2xp33_ASAP7_75t_SL g14769 ( 
.A(n_14742),
.B(n_2945),
.Y(n_14769)
);

NAND2xp5_ASAP7_75t_L g14770 ( 
.A(n_14685),
.B(n_2946),
.Y(n_14770)
);

AND2x2_ASAP7_75t_L g14771 ( 
.A(n_14684),
.B(n_2946),
.Y(n_14771)
);

INVx1_ASAP7_75t_L g14772 ( 
.A(n_14695),
.Y(n_14772)
);

AOI21xp5_ASAP7_75t_L g14773 ( 
.A1(n_14731),
.A2(n_2948),
.B(n_2949),
.Y(n_14773)
);

NOR2xp33_ASAP7_75t_R g14774 ( 
.A(n_14707),
.B(n_2950),
.Y(n_14774)
);

AND2x2_ASAP7_75t_L g14775 ( 
.A(n_14700),
.B(n_2948),
.Y(n_14775)
);

BUFx2_ASAP7_75t_L g14776 ( 
.A(n_14745),
.Y(n_14776)
);

INVx1_ASAP7_75t_L g14777 ( 
.A(n_14694),
.Y(n_14777)
);

OAI211xp5_ASAP7_75t_L g14778 ( 
.A1(n_14747),
.A2(n_2952),
.B(n_2953),
.C(n_2951),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14733),
.Y(n_14779)
);

INVx1_ASAP7_75t_L g14780 ( 
.A(n_14753),
.Y(n_14780)
);

BUFx6f_ASAP7_75t_L g14781 ( 
.A(n_14683),
.Y(n_14781)
);

AOI211xp5_ASAP7_75t_L g14782 ( 
.A1(n_14689),
.A2(n_2952),
.B(n_2950),
.C(n_2951),
.Y(n_14782)
);

XNOR2xp5_ASAP7_75t_L g14783 ( 
.A(n_14703),
.B(n_2953),
.Y(n_14783)
);

AOI21xp5_ASAP7_75t_L g14784 ( 
.A1(n_14691),
.A2(n_2954),
.B(n_2955),
.Y(n_14784)
);

AOI21x1_ASAP7_75t_L g14785 ( 
.A1(n_14697),
.A2(n_2959),
.B(n_2958),
.Y(n_14785)
);

NOR2xp33_ASAP7_75t_R g14786 ( 
.A(n_14696),
.B(n_2958),
.Y(n_14786)
);

OAI21xp5_ASAP7_75t_SL g14787 ( 
.A1(n_14722),
.A2(n_14702),
.B(n_14725),
.Y(n_14787)
);

AOI31xp33_ASAP7_75t_L g14788 ( 
.A1(n_14709),
.A2(n_2960),
.A3(n_2957),
.B(n_2959),
.Y(n_14788)
);

BUFx2_ASAP7_75t_L g14789 ( 
.A(n_14736),
.Y(n_14789)
);

INVx1_ASAP7_75t_L g14790 ( 
.A(n_14736),
.Y(n_14790)
);

NAND2xp5_ASAP7_75t_L g14791 ( 
.A(n_14708),
.B(n_2957),
.Y(n_14791)
);

NAND2xp33_ASAP7_75t_L g14792 ( 
.A(n_14721),
.B(n_2961),
.Y(n_14792)
);

NAND2xp5_ASAP7_75t_L g14793 ( 
.A(n_14728),
.B(n_2961),
.Y(n_14793)
);

INVx1_ASAP7_75t_L g14794 ( 
.A(n_14690),
.Y(n_14794)
);

NAND2xp5_ASAP7_75t_SL g14795 ( 
.A(n_14730),
.B(n_2962),
.Y(n_14795)
);

AOI21xp33_ASAP7_75t_L g14796 ( 
.A1(n_14715),
.A2(n_2962),
.B(n_2963),
.Y(n_14796)
);

XOR2xp5_ASAP7_75t_L g14797 ( 
.A(n_14732),
.B(n_2963),
.Y(n_14797)
);

AOI221xp5_ASAP7_75t_L g14798 ( 
.A1(n_14714),
.A2(n_14723),
.B1(n_14739),
.B2(n_14726),
.C(n_14751),
.Y(n_14798)
);

AND3x4_ASAP7_75t_L g14799 ( 
.A(n_14711),
.B(n_2964),
.C(n_2965),
.Y(n_14799)
);

HB1xp67_ASAP7_75t_L g14800 ( 
.A(n_14706),
.Y(n_14800)
);

HB1xp67_ASAP7_75t_L g14801 ( 
.A(n_14750),
.Y(n_14801)
);

XOR2xp5_ASAP7_75t_L g14802 ( 
.A(n_14729),
.B(n_2964),
.Y(n_14802)
);

OAI21xp33_ASAP7_75t_L g14803 ( 
.A1(n_14756),
.A2(n_2965),
.B(n_2966),
.Y(n_14803)
);

NAND2xp33_ASAP7_75t_R g14804 ( 
.A(n_14724),
.B(n_2968),
.Y(n_14804)
);

INVx2_ASAP7_75t_SL g14805 ( 
.A(n_14738),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14687),
.Y(n_14806)
);

AND2x2_ASAP7_75t_SL g14807 ( 
.A(n_14741),
.B(n_2967),
.Y(n_14807)
);

HB1xp67_ASAP7_75t_L g14808 ( 
.A(n_14746),
.Y(n_14808)
);

NOR2x1_ASAP7_75t_L g14809 ( 
.A(n_14716),
.B(n_3350),
.Y(n_14809)
);

NAND4xp25_ASAP7_75t_SL g14810 ( 
.A(n_14705),
.B(n_2969),
.C(n_2967),
.D(n_2968),
.Y(n_14810)
);

AOI211xp5_ASAP7_75t_L g14811 ( 
.A1(n_14701),
.A2(n_2972),
.B(n_2969),
.C(n_2971),
.Y(n_14811)
);

OAI21xp5_ASAP7_75t_SL g14812 ( 
.A1(n_14744),
.A2(n_2971),
.B(n_2972),
.Y(n_14812)
);

NAND4xp25_ASAP7_75t_L g14813 ( 
.A(n_14735),
.B(n_3357),
.C(n_2975),
.D(n_2973),
.Y(n_14813)
);

BUFx2_ASAP7_75t_L g14814 ( 
.A(n_14754),
.Y(n_14814)
);

NAND2xp5_ASAP7_75t_L g14815 ( 
.A(n_14757),
.B(n_2973),
.Y(n_14815)
);

XNOR2xp5_ASAP7_75t_L g14816 ( 
.A(n_14719),
.B(n_2974),
.Y(n_14816)
);

OAI211xp5_ASAP7_75t_L g14817 ( 
.A1(n_14713),
.A2(n_2976),
.B(n_2977),
.C(n_2975),
.Y(n_14817)
);

NAND5xp2_ASAP7_75t_L g14818 ( 
.A(n_14798),
.B(n_14712),
.C(n_14734),
.D(n_14737),
.E(n_14692),
.Y(n_14818)
);

NAND4xp25_ASAP7_75t_L g14819 ( 
.A(n_14796),
.B(n_14755),
.C(n_14727),
.D(n_14693),
.Y(n_14819)
);

NAND2xp5_ASAP7_75t_L g14820 ( 
.A(n_14807),
.B(n_14752),
.Y(n_14820)
);

OR2x2_ASAP7_75t_L g14821 ( 
.A(n_14770),
.B(n_14718),
.Y(n_14821)
);

NOR4xp25_ASAP7_75t_L g14822 ( 
.A(n_14790),
.B(n_14765),
.C(n_14780),
.D(n_14794),
.Y(n_14822)
);

NOR2x1_ASAP7_75t_L g14823 ( 
.A(n_14789),
.B(n_14720),
.Y(n_14823)
);

NAND2xp5_ASAP7_75t_L g14824 ( 
.A(n_14775),
.B(n_14710),
.Y(n_14824)
);

NOR2x1_ASAP7_75t_L g14825 ( 
.A(n_14777),
.B(n_2974),
.Y(n_14825)
);

BUFx2_ASAP7_75t_L g14826 ( 
.A(n_14774),
.Y(n_14826)
);

INVx3_ASAP7_75t_L g14827 ( 
.A(n_14785),
.Y(n_14827)
);

NAND3xp33_ASAP7_75t_L g14828 ( 
.A(n_14781),
.B(n_2985),
.C(n_2977),
.Y(n_14828)
);

NAND4xp25_ASAP7_75t_L g14829 ( 
.A(n_14782),
.B(n_2980),
.C(n_2978),
.D(n_2979),
.Y(n_14829)
);

NAND2xp5_ASAP7_75t_L g14830 ( 
.A(n_14784),
.B(n_2978),
.Y(n_14830)
);

AND2x2_ASAP7_75t_L g14831 ( 
.A(n_14809),
.B(n_14771),
.Y(n_14831)
);

XNOR2x1_ASAP7_75t_L g14832 ( 
.A(n_14799),
.B(n_14783),
.Y(n_14832)
);

NOR3xp33_ASAP7_75t_SL g14833 ( 
.A(n_14766),
.B(n_2980),
.C(n_2981),
.Y(n_14833)
);

INVx2_ASAP7_75t_L g14834 ( 
.A(n_14767),
.Y(n_14834)
);

NOR2x1_ASAP7_75t_L g14835 ( 
.A(n_14763),
.B(n_2981),
.Y(n_14835)
);

NAND5xp2_ASAP7_75t_L g14836 ( 
.A(n_14769),
.B(n_2984),
.C(n_2982),
.D(n_2983),
.E(n_2985),
.Y(n_14836)
);

NAND3xp33_ASAP7_75t_SL g14837 ( 
.A(n_14761),
.B(n_2983),
.C(n_2984),
.Y(n_14837)
);

NAND3xp33_ASAP7_75t_L g14838 ( 
.A(n_14781),
.B(n_14804),
.C(n_14772),
.Y(n_14838)
);

BUFx3_ASAP7_75t_L g14839 ( 
.A(n_14776),
.Y(n_14839)
);

INVxp67_ASAP7_75t_SL g14840 ( 
.A(n_14759),
.Y(n_14840)
);

OR2x6_ASAP7_75t_L g14841 ( 
.A(n_14805),
.B(n_2986),
.Y(n_14841)
);

NOR2x1_ASAP7_75t_L g14842 ( 
.A(n_14813),
.B(n_2986),
.Y(n_14842)
);

NAND3xp33_ASAP7_75t_SL g14843 ( 
.A(n_14786),
.B(n_2987),
.C(n_2988),
.Y(n_14843)
);

NAND4xp25_ASAP7_75t_SL g14844 ( 
.A(n_14811),
.B(n_2989),
.C(n_2987),
.D(n_2988),
.Y(n_14844)
);

INVx1_ASAP7_75t_L g14845 ( 
.A(n_14768),
.Y(n_14845)
);

NAND2xp5_ASAP7_75t_L g14846 ( 
.A(n_14788),
.B(n_2990),
.Y(n_14846)
);

NOR3xp33_ASAP7_75t_SL g14847 ( 
.A(n_14812),
.B(n_2991),
.C(n_2992),
.Y(n_14847)
);

AND3x2_ASAP7_75t_L g14848 ( 
.A(n_14801),
.B(n_2994),
.C(n_2993),
.Y(n_14848)
);

NOR2x1p5_ASAP7_75t_L g14849 ( 
.A(n_14815),
.B(n_2992),
.Y(n_14849)
);

NOR2xp33_ASAP7_75t_L g14850 ( 
.A(n_14803),
.B(n_2993),
.Y(n_14850)
);

AND2x2_ASAP7_75t_SL g14851 ( 
.A(n_14792),
.B(n_2995),
.Y(n_14851)
);

NOR2x1_ASAP7_75t_L g14852 ( 
.A(n_14817),
.B(n_2996),
.Y(n_14852)
);

NOR2x1_ASAP7_75t_L g14853 ( 
.A(n_14810),
.B(n_2996),
.Y(n_14853)
);

NAND3xp33_ASAP7_75t_SL g14854 ( 
.A(n_14764),
.B(n_2997),
.C(n_2998),
.Y(n_14854)
);

AO211x2_ASAP7_75t_L g14855 ( 
.A1(n_14773),
.A2(n_3000),
.B(n_2997),
.C(n_2999),
.Y(n_14855)
);

NAND3xp33_ASAP7_75t_SL g14856 ( 
.A(n_14778),
.B(n_3000),
.C(n_3001),
.Y(n_14856)
);

NAND5xp2_ASAP7_75t_L g14857 ( 
.A(n_14787),
.B(n_3003),
.C(n_3001),
.D(n_3002),
.E(n_3004),
.Y(n_14857)
);

NAND4xp25_ASAP7_75t_L g14858 ( 
.A(n_14791),
.B(n_3004),
.C(n_3002),
.D(n_3003),
.Y(n_14858)
);

O2A1O1Ixp5_ASAP7_75t_L g14859 ( 
.A1(n_14795),
.A2(n_3007),
.B(n_3005),
.C(n_3006),
.Y(n_14859)
);

AND2x2_ASAP7_75t_L g14860 ( 
.A(n_14808),
.B(n_3005),
.Y(n_14860)
);

NOR3xp33_ASAP7_75t_L g14861 ( 
.A(n_14800),
.B(n_14779),
.C(n_14806),
.Y(n_14861)
);

OAI21xp5_ASAP7_75t_L g14862 ( 
.A1(n_14802),
.A2(n_3008),
.B(n_3009),
.Y(n_14862)
);

NOR2x1_ASAP7_75t_L g14863 ( 
.A(n_14816),
.B(n_14797),
.Y(n_14863)
);

NAND4xp75_ASAP7_75t_L g14864 ( 
.A(n_14823),
.B(n_14793),
.C(n_14758),
.D(n_14762),
.Y(n_14864)
);

OR2x2_ASAP7_75t_L g14865 ( 
.A(n_14836),
.B(n_14781),
.Y(n_14865)
);

NAND4xp75_ASAP7_75t_L g14866 ( 
.A(n_14863),
.B(n_14814),
.C(n_14760),
.D(n_3010),
.Y(n_14866)
);

NOR3xp33_ASAP7_75t_L g14867 ( 
.A(n_14838),
.B(n_3008),
.C(n_3009),
.Y(n_14867)
);

NOR3xp33_ASAP7_75t_SL g14868 ( 
.A(n_14818),
.B(n_3019),
.C(n_3011),
.Y(n_14868)
);

A2O1A1Ixp33_ASAP7_75t_L g14869 ( 
.A1(n_14859),
.A2(n_3013),
.B(n_3011),
.C(n_3012),
.Y(n_14869)
);

NOR3xp33_ASAP7_75t_L g14870 ( 
.A(n_14840),
.B(n_3012),
.C(n_3013),
.Y(n_14870)
);

NAND4xp75_ASAP7_75t_L g14871 ( 
.A(n_14831),
.B(n_3016),
.C(n_3014),
.D(n_3015),
.Y(n_14871)
);

HB1xp67_ASAP7_75t_L g14872 ( 
.A(n_14825),
.Y(n_14872)
);

A2O1A1Ixp33_ASAP7_75t_L g14873 ( 
.A1(n_14850),
.A2(n_3016),
.B(n_3014),
.C(n_3015),
.Y(n_14873)
);

INVx2_ASAP7_75t_L g14874 ( 
.A(n_14841),
.Y(n_14874)
);

AND2x2_ASAP7_75t_L g14875 ( 
.A(n_14847),
.B(n_3017),
.Y(n_14875)
);

OR2x6_ASAP7_75t_L g14876 ( 
.A(n_14834),
.B(n_3017),
.Y(n_14876)
);

AOI22xp5_ASAP7_75t_L g14877 ( 
.A1(n_14844),
.A2(n_3020),
.B1(n_3021),
.B2(n_3019),
.Y(n_14877)
);

NAND4xp25_ASAP7_75t_L g14878 ( 
.A(n_14861),
.B(n_3022),
.C(n_3018),
.D(n_3020),
.Y(n_14878)
);

AND2x2_ASAP7_75t_L g14879 ( 
.A(n_14842),
.B(n_3018),
.Y(n_14879)
);

NAND5xp2_ASAP7_75t_L g14880 ( 
.A(n_14833),
.B(n_3024),
.C(n_3022),
.D(n_3023),
.E(n_3025),
.Y(n_14880)
);

NOR2x1p5_ASAP7_75t_L g14881 ( 
.A(n_14846),
.B(n_3023),
.Y(n_14881)
);

NAND4xp75_ASAP7_75t_L g14882 ( 
.A(n_14835),
.B(n_14853),
.C(n_14845),
.D(n_14852),
.Y(n_14882)
);

AOI211xp5_ASAP7_75t_L g14883 ( 
.A1(n_14843),
.A2(n_3026),
.B(n_3024),
.C(n_3025),
.Y(n_14883)
);

CKINVDCx5p33_ASAP7_75t_R g14884 ( 
.A(n_14839),
.Y(n_14884)
);

NOR2x1_ASAP7_75t_L g14885 ( 
.A(n_14827),
.B(n_3026),
.Y(n_14885)
);

NOR3xp33_ASAP7_75t_L g14886 ( 
.A(n_14826),
.B(n_3027),
.C(n_3028),
.Y(n_14886)
);

NOR2xp33_ASAP7_75t_L g14887 ( 
.A(n_14856),
.B(n_3027),
.Y(n_14887)
);

NOR3x1_ASAP7_75t_L g14888 ( 
.A(n_14862),
.B(n_3028),
.C(n_3029),
.Y(n_14888)
);

INVx3_ASAP7_75t_SL g14889 ( 
.A(n_14832),
.Y(n_14889)
);

NAND2xp5_ASAP7_75t_L g14890 ( 
.A(n_14848),
.B(n_3029),
.Y(n_14890)
);

OR2x2_ASAP7_75t_L g14891 ( 
.A(n_14857),
.B(n_3030),
.Y(n_14891)
);

NOR4xp75_ASAP7_75t_L g14892 ( 
.A(n_14820),
.B(n_3032),
.C(n_3030),
.D(n_3031),
.Y(n_14892)
);

NAND4xp25_ASAP7_75t_L g14893 ( 
.A(n_14824),
.B(n_3034),
.C(n_3031),
.D(n_3032),
.Y(n_14893)
);

NAND4xp75_ASAP7_75t_L g14894 ( 
.A(n_14851),
.B(n_3039),
.C(n_3035),
.D(n_3037),
.Y(n_14894)
);

OAI211xp5_ASAP7_75t_SL g14895 ( 
.A1(n_14821),
.A2(n_3040),
.B(n_3035),
.C(n_3039),
.Y(n_14895)
);

INVx1_ASAP7_75t_L g14896 ( 
.A(n_14849),
.Y(n_14896)
);

OAI22xp5_ASAP7_75t_L g14897 ( 
.A1(n_14830),
.A2(n_3042),
.B1(n_3040),
.B2(n_3041),
.Y(n_14897)
);

NAND2xp5_ASAP7_75t_L g14898 ( 
.A(n_14860),
.B(n_3042),
.Y(n_14898)
);

NAND3xp33_ASAP7_75t_L g14899 ( 
.A(n_14822),
.B(n_3044),
.C(n_3045),
.Y(n_14899)
);

AND3x4_ASAP7_75t_L g14900 ( 
.A(n_14855),
.B(n_3044),
.C(n_3046),
.Y(n_14900)
);

AOI211xp5_ASAP7_75t_L g14901 ( 
.A1(n_14854),
.A2(n_3048),
.B(n_3046),
.C(n_3047),
.Y(n_14901)
);

OAI22xp5_ASAP7_75t_L g14902 ( 
.A1(n_14828),
.A2(n_3049),
.B1(n_3047),
.B2(n_3048),
.Y(n_14902)
);

NOR2x1_ASAP7_75t_L g14903 ( 
.A(n_14837),
.B(n_3050),
.Y(n_14903)
);

OAI21xp5_ASAP7_75t_L g14904 ( 
.A1(n_14829),
.A2(n_3051),
.B(n_3052),
.Y(n_14904)
);

INVx1_ASAP7_75t_L g14905 ( 
.A(n_14841),
.Y(n_14905)
);

NAND2x1p5_ASAP7_75t_L g14906 ( 
.A(n_14819),
.B(n_3051),
.Y(n_14906)
);

NAND3xp33_ASAP7_75t_SL g14907 ( 
.A(n_14858),
.B(n_3052),
.C(n_3053),
.Y(n_14907)
);

NOR4xp25_ASAP7_75t_L g14908 ( 
.A(n_14838),
.B(n_3055),
.C(n_3053),
.D(n_3054),
.Y(n_14908)
);

XNOR2x1_ASAP7_75t_L g14909 ( 
.A(n_14884),
.B(n_3055),
.Y(n_14909)
);

XNOR2x1_ASAP7_75t_L g14910 ( 
.A(n_14900),
.B(n_3056),
.Y(n_14910)
);

INVx1_ASAP7_75t_L g14911 ( 
.A(n_14906),
.Y(n_14911)
);

INVx1_ASAP7_75t_L g14912 ( 
.A(n_14890),
.Y(n_14912)
);

OAI211xp5_ASAP7_75t_L g14913 ( 
.A1(n_14899),
.A2(n_3357),
.B(n_3358),
.C(n_3356),
.Y(n_14913)
);

AOI211xp5_ASAP7_75t_SL g14914 ( 
.A1(n_14865),
.A2(n_3058),
.B(n_3056),
.C(n_3057),
.Y(n_14914)
);

NAND2xp5_ASAP7_75t_L g14915 ( 
.A(n_14885),
.B(n_3058),
.Y(n_14915)
);

INVxp33_ASAP7_75t_L g14916 ( 
.A(n_14868),
.Y(n_14916)
);

INVx1_ASAP7_75t_L g14917 ( 
.A(n_14881),
.Y(n_14917)
);

INVx2_ASAP7_75t_L g14918 ( 
.A(n_14871),
.Y(n_14918)
);

INVx2_ASAP7_75t_L g14919 ( 
.A(n_14894),
.Y(n_14919)
);

NAND2xp5_ASAP7_75t_L g14920 ( 
.A(n_14877),
.B(n_3059),
.Y(n_14920)
);

OR2x2_ASAP7_75t_L g14921 ( 
.A(n_14880),
.B(n_3057),
.Y(n_14921)
);

INVx1_ASAP7_75t_SL g14922 ( 
.A(n_14879),
.Y(n_14922)
);

AOI22xp33_ASAP7_75t_L g14923 ( 
.A1(n_14907),
.A2(n_3061),
.B1(n_3059),
.B2(n_3060),
.Y(n_14923)
);

NAND2xp5_ASAP7_75t_L g14924 ( 
.A(n_14883),
.B(n_3062),
.Y(n_14924)
);

NAND2x1_ASAP7_75t_L g14925 ( 
.A(n_14903),
.B(n_3060),
.Y(n_14925)
);

NAND2xp5_ASAP7_75t_L g14926 ( 
.A(n_14901),
.B(n_3063),
.Y(n_14926)
);

OAI22xp5_ASAP7_75t_L g14927 ( 
.A1(n_14891),
.A2(n_3064),
.B1(n_3062),
.B2(n_3063),
.Y(n_14927)
);

AND2x2_ASAP7_75t_L g14928 ( 
.A(n_14875),
.B(n_3064),
.Y(n_14928)
);

OA22x2_ASAP7_75t_L g14929 ( 
.A1(n_14904),
.A2(n_14902),
.B1(n_14889),
.B2(n_14905),
.Y(n_14929)
);

OAI22xp5_ASAP7_75t_L g14930 ( 
.A1(n_14873),
.A2(n_3067),
.B1(n_3065),
.B2(n_3066),
.Y(n_14930)
);

AOI221xp5_ASAP7_75t_L g14931 ( 
.A1(n_14908),
.A2(n_3067),
.B1(n_3065),
.B2(n_3066),
.C(n_3068),
.Y(n_14931)
);

OAI22xp5_ASAP7_75t_L g14932 ( 
.A1(n_14869),
.A2(n_3072),
.B1(n_3069),
.B2(n_3071),
.Y(n_14932)
);

NAND2xp5_ASAP7_75t_L g14933 ( 
.A(n_14867),
.B(n_3072),
.Y(n_14933)
);

INVx1_ASAP7_75t_L g14934 ( 
.A(n_14888),
.Y(n_14934)
);

NAND2x1_ASAP7_75t_L g14935 ( 
.A(n_14874),
.B(n_3069),
.Y(n_14935)
);

XNOR2xp5_ASAP7_75t_L g14936 ( 
.A(n_14864),
.B(n_3073),
.Y(n_14936)
);

OA22x2_ASAP7_75t_L g14937 ( 
.A1(n_14872),
.A2(n_3082),
.B1(n_3090),
.B2(n_3073),
.Y(n_14937)
);

AND3x4_ASAP7_75t_L g14938 ( 
.A(n_14892),
.B(n_14870),
.C(n_14886),
.Y(n_14938)
);

AOI22xp5_ASAP7_75t_L g14939 ( 
.A1(n_14887),
.A2(n_14895),
.B1(n_14866),
.B2(n_14896),
.Y(n_14939)
);

NAND2x1_ASAP7_75t_L g14940 ( 
.A(n_14898),
.B(n_3074),
.Y(n_14940)
);

INVxp67_ASAP7_75t_SL g14941 ( 
.A(n_14897),
.Y(n_14941)
);

OAI22xp5_ASAP7_75t_L g14942 ( 
.A1(n_14882),
.A2(n_3078),
.B1(n_3076),
.B2(n_3077),
.Y(n_14942)
);

XNOR2xp5_ASAP7_75t_L g14943 ( 
.A(n_14878),
.B(n_3076),
.Y(n_14943)
);

INVx1_ASAP7_75t_L g14944 ( 
.A(n_14893),
.Y(n_14944)
);

BUFx2_ASAP7_75t_L g14945 ( 
.A(n_14876),
.Y(n_14945)
);

AND2x2_ASAP7_75t_L g14946 ( 
.A(n_14876),
.B(n_3077),
.Y(n_14946)
);

AND2x2_ASAP7_75t_L g14947 ( 
.A(n_14868),
.B(n_3078),
.Y(n_14947)
);

BUFx2_ASAP7_75t_L g14948 ( 
.A(n_14885),
.Y(n_14948)
);

NOR3xp33_ASAP7_75t_L g14949 ( 
.A(n_14864),
.B(n_3079),
.C(n_3080),
.Y(n_14949)
);

INVx1_ASAP7_75t_L g14950 ( 
.A(n_14906),
.Y(n_14950)
);

INVx1_ASAP7_75t_L g14951 ( 
.A(n_14928),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14936),
.Y(n_14952)
);

HB1xp67_ASAP7_75t_L g14953 ( 
.A(n_14935),
.Y(n_14953)
);

INVx1_ASAP7_75t_L g14954 ( 
.A(n_14915),
.Y(n_14954)
);

BUFx2_ASAP7_75t_L g14955 ( 
.A(n_14946),
.Y(n_14955)
);

INVx3_ASAP7_75t_L g14956 ( 
.A(n_14925),
.Y(n_14956)
);

INVx1_ASAP7_75t_L g14957 ( 
.A(n_14940),
.Y(n_14957)
);

INVx1_ASAP7_75t_L g14958 ( 
.A(n_14921),
.Y(n_14958)
);

INVx1_ASAP7_75t_L g14959 ( 
.A(n_14947),
.Y(n_14959)
);

INVx1_ASAP7_75t_L g14960 ( 
.A(n_14943),
.Y(n_14960)
);

NAND2x1_ASAP7_75t_L g14961 ( 
.A(n_14948),
.B(n_3079),
.Y(n_14961)
);

INVx1_ASAP7_75t_L g14962 ( 
.A(n_14920),
.Y(n_14962)
);

INVxp67_ASAP7_75t_L g14963 ( 
.A(n_14910),
.Y(n_14963)
);

INVx1_ASAP7_75t_L g14964 ( 
.A(n_14933),
.Y(n_14964)
);

INVx1_ASAP7_75t_SL g14965 ( 
.A(n_14909),
.Y(n_14965)
);

INVx2_ASAP7_75t_L g14966 ( 
.A(n_14937),
.Y(n_14966)
);

INVx1_ASAP7_75t_L g14967 ( 
.A(n_14924),
.Y(n_14967)
);

INVx1_ASAP7_75t_L g14968 ( 
.A(n_14926),
.Y(n_14968)
);

INVx1_ASAP7_75t_L g14969 ( 
.A(n_14913),
.Y(n_14969)
);

INVx2_ASAP7_75t_L g14970 ( 
.A(n_14938),
.Y(n_14970)
);

INVx1_ASAP7_75t_L g14971 ( 
.A(n_14932),
.Y(n_14971)
);

INVx1_ASAP7_75t_SL g14972 ( 
.A(n_14945),
.Y(n_14972)
);

OAI22xp33_ASAP7_75t_L g14973 ( 
.A1(n_14916),
.A2(n_3082),
.B1(n_3080),
.B2(n_3081),
.Y(n_14973)
);

AOI22xp5_ASAP7_75t_L g14974 ( 
.A1(n_14949),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.Y(n_14974)
);

INVx1_ASAP7_75t_L g14975 ( 
.A(n_14927),
.Y(n_14975)
);

AOI22xp5_ASAP7_75t_L g14976 ( 
.A1(n_14930),
.A2(n_3086),
.B1(n_3083),
.B2(n_3084),
.Y(n_14976)
);

CKINVDCx20_ASAP7_75t_R g14977 ( 
.A(n_14939),
.Y(n_14977)
);

INVx1_ASAP7_75t_L g14978 ( 
.A(n_14934),
.Y(n_14978)
);

INVx1_ASAP7_75t_L g14979 ( 
.A(n_14919),
.Y(n_14979)
);

INVx5_ASAP7_75t_L g14980 ( 
.A(n_14918),
.Y(n_14980)
);

INVxp67_ASAP7_75t_L g14981 ( 
.A(n_14911),
.Y(n_14981)
);

INVx1_ASAP7_75t_L g14982 ( 
.A(n_14923),
.Y(n_14982)
);

INVx1_ASAP7_75t_L g14983 ( 
.A(n_14917),
.Y(n_14983)
);

INVx1_ASAP7_75t_L g14984 ( 
.A(n_14950),
.Y(n_14984)
);

OAI22xp33_ASAP7_75t_L g14985 ( 
.A1(n_14914),
.A2(n_3088),
.B1(n_3086),
.B2(n_3087),
.Y(n_14985)
);

INVx2_ASAP7_75t_L g14986 ( 
.A(n_14942),
.Y(n_14986)
);

INVx2_ASAP7_75t_L g14987 ( 
.A(n_14944),
.Y(n_14987)
);

INVx1_ASAP7_75t_L g14988 ( 
.A(n_14929),
.Y(n_14988)
);

INVx1_ASAP7_75t_L g14989 ( 
.A(n_14912),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14941),
.Y(n_14990)
);

OR3x2_ASAP7_75t_L g14991 ( 
.A(n_14922),
.B(n_3087),
.C(n_3089),
.Y(n_14991)
);

HB1xp67_ASAP7_75t_L g14992 ( 
.A(n_14961),
.Y(n_14992)
);

OAI21xp5_ASAP7_75t_L g14993 ( 
.A1(n_14981),
.A2(n_14931),
.B(n_3089),
.Y(n_14993)
);

OR2x2_ASAP7_75t_L g14994 ( 
.A(n_14974),
.B(n_3090),
.Y(n_14994)
);

NAND2x1p5_ASAP7_75t_L g14995 ( 
.A(n_14956),
.B(n_3091),
.Y(n_14995)
);

NAND2xp5_ASAP7_75t_L g14996 ( 
.A(n_14985),
.B(n_3369),
.Y(n_14996)
);

NAND2xp5_ASAP7_75t_L g14997 ( 
.A(n_14976),
.B(n_3092),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14991),
.Y(n_14998)
);

INVx1_ASAP7_75t_L g14999 ( 
.A(n_14953),
.Y(n_14999)
);

HB1xp67_ASAP7_75t_L g15000 ( 
.A(n_14988),
.Y(n_15000)
);

OAI221xp5_ASAP7_75t_L g15001 ( 
.A1(n_14972),
.A2(n_3094),
.B1(n_3092),
.B2(n_3093),
.C(n_3095),
.Y(n_15001)
);

CKINVDCx5p33_ASAP7_75t_R g15002 ( 
.A(n_14977),
.Y(n_15002)
);

INVx1_ASAP7_75t_L g15003 ( 
.A(n_14955),
.Y(n_15003)
);

NOR2x1_ASAP7_75t_L g15004 ( 
.A(n_14957),
.B(n_3094),
.Y(n_15004)
);

HB1xp67_ASAP7_75t_L g15005 ( 
.A(n_14990),
.Y(n_15005)
);

OAI22xp5_ASAP7_75t_L g15006 ( 
.A1(n_14980),
.A2(n_3096),
.B1(n_3097),
.B2(n_3095),
.Y(n_15006)
);

HB1xp67_ASAP7_75t_L g15007 ( 
.A(n_14980),
.Y(n_15007)
);

INVx1_ASAP7_75t_SL g15008 ( 
.A(n_14965),
.Y(n_15008)
);

OR3x2_ASAP7_75t_L g15009 ( 
.A(n_14984),
.B(n_3093),
.C(n_3096),
.Y(n_15009)
);

AND2x4_ASAP7_75t_L g15010 ( 
.A(n_14966),
.B(n_3097),
.Y(n_15010)
);

OR2x2_ASAP7_75t_L g15011 ( 
.A(n_14978),
.B(n_3098),
.Y(n_15011)
);

BUFx2_ASAP7_75t_L g15012 ( 
.A(n_14969),
.Y(n_15012)
);

CKINVDCx20_ASAP7_75t_R g15013 ( 
.A(n_14970),
.Y(n_15013)
);

INVx1_ASAP7_75t_L g15014 ( 
.A(n_14951),
.Y(n_15014)
);

OR2x2_ASAP7_75t_L g15015 ( 
.A(n_14979),
.B(n_3098),
.Y(n_15015)
);

INVx1_ASAP7_75t_SL g15016 ( 
.A(n_14980),
.Y(n_15016)
);

CKINVDCx5p33_ASAP7_75t_R g15017 ( 
.A(n_14958),
.Y(n_15017)
);

INVx1_ASAP7_75t_L g15018 ( 
.A(n_14975),
.Y(n_15018)
);

AOI22xp5_ASAP7_75t_L g15019 ( 
.A1(n_15002),
.A2(n_14983),
.B1(n_14989),
.B2(n_14987),
.Y(n_15019)
);

AOI22xp5_ASAP7_75t_L g15020 ( 
.A1(n_15013),
.A2(n_14952),
.B1(n_14982),
.B2(n_14986),
.Y(n_15020)
);

INVx1_ASAP7_75t_L g15021 ( 
.A(n_14996),
.Y(n_15021)
);

INVx1_ASAP7_75t_L g15022 ( 
.A(n_14997),
.Y(n_15022)
);

INVx1_ASAP7_75t_L g15023 ( 
.A(n_14994),
.Y(n_15023)
);

INVx1_ASAP7_75t_SL g15024 ( 
.A(n_15016),
.Y(n_15024)
);

OA22x2_ASAP7_75t_L g15025 ( 
.A1(n_14993),
.A2(n_15007),
.B1(n_14999),
.B2(n_15000),
.Y(n_15025)
);

AOI22xp5_ASAP7_75t_L g15026 ( 
.A1(n_15003),
.A2(n_14963),
.B1(n_14959),
.B2(n_14954),
.Y(n_15026)
);

HB1xp67_ASAP7_75t_L g15027 ( 
.A(n_15004),
.Y(n_15027)
);

INVx1_ASAP7_75t_L g15028 ( 
.A(n_15005),
.Y(n_15028)
);

INVx1_ASAP7_75t_L g15029 ( 
.A(n_14992),
.Y(n_15029)
);

AOI22xp5_ASAP7_75t_L g15030 ( 
.A1(n_15014),
.A2(n_14960),
.B1(n_14962),
.B2(n_14964),
.Y(n_15030)
);

OAI22x1_ASAP7_75t_L g15031 ( 
.A1(n_15018),
.A2(n_14971),
.B1(n_14968),
.B2(n_14967),
.Y(n_15031)
);

AOI22xp5_ASAP7_75t_L g15032 ( 
.A1(n_15008),
.A2(n_14973),
.B1(n_3101),
.B2(n_3099),
.Y(n_15032)
);

A2O1A1Ixp33_ASAP7_75t_SL g15033 ( 
.A1(n_14998),
.A2(n_3104),
.B(n_3100),
.C(n_3103),
.Y(n_15033)
);

OAI22xp5_ASAP7_75t_L g15034 ( 
.A1(n_15009),
.A2(n_3104),
.B1(n_3100),
.B2(n_3103),
.Y(n_15034)
);

AO22x2_ASAP7_75t_L g15035 ( 
.A1(n_15012),
.A2(n_3107),
.B1(n_3105),
.B2(n_3106),
.Y(n_15035)
);

INVx1_ASAP7_75t_L g15036 ( 
.A(n_14995),
.Y(n_15036)
);

INVx1_ASAP7_75t_L g15037 ( 
.A(n_15017),
.Y(n_15037)
);

AOI22xp5_ASAP7_75t_L g15038 ( 
.A1(n_15001),
.A2(n_3107),
.B1(n_3105),
.B2(n_3106),
.Y(n_15038)
);

AOI22xp5_ASAP7_75t_L g15039 ( 
.A1(n_15024),
.A2(n_15006),
.B1(n_15010),
.B2(n_15015),
.Y(n_15039)
);

AND4x1_ASAP7_75t_L g15040 ( 
.A(n_15019),
.B(n_15010),
.C(n_15011),
.D(n_3110),
.Y(n_15040)
);

XNOR2xp5_ASAP7_75t_L g15041 ( 
.A(n_15020),
.B(n_3108),
.Y(n_15041)
);

NOR2x1p5_ASAP7_75t_L g15042 ( 
.A(n_15028),
.B(n_3109),
.Y(n_15042)
);

NOR3xp33_ASAP7_75t_L g15043 ( 
.A(n_15029),
.B(n_3108),
.C(n_3109),
.Y(n_15043)
);

NAND3xp33_ASAP7_75t_L g15044 ( 
.A(n_15026),
.B(n_3110),
.C(n_3111),
.Y(n_15044)
);

AOI221xp5_ASAP7_75t_SL g15045 ( 
.A1(n_15031),
.A2(n_3113),
.B1(n_3115),
.B2(n_3112),
.C(n_3114),
.Y(n_15045)
);

INVx1_ASAP7_75t_L g15046 ( 
.A(n_15032),
.Y(n_15046)
);

OAI221xp5_ASAP7_75t_L g15047 ( 
.A1(n_15038),
.A2(n_3114),
.B1(n_3111),
.B2(n_3113),
.C(n_3116),
.Y(n_15047)
);

AOI22xp5_ASAP7_75t_L g15048 ( 
.A1(n_15034),
.A2(n_3124),
.B1(n_3133),
.B2(n_3116),
.Y(n_15048)
);

NAND4xp25_ASAP7_75t_L g15049 ( 
.A(n_15030),
.B(n_3119),
.C(n_3117),
.D(n_3118),
.Y(n_15049)
);

OR5x1_ASAP7_75t_L g15050 ( 
.A(n_15025),
.B(n_3120),
.C(n_3117),
.D(n_3119),
.E(n_3121),
.Y(n_15050)
);

OAI221xp5_ASAP7_75t_L g15051 ( 
.A1(n_15033),
.A2(n_3124),
.B1(n_3122),
.B2(n_3123),
.C(n_3125),
.Y(n_15051)
);

AOI22xp33_ASAP7_75t_L g15052 ( 
.A1(n_15037),
.A2(n_3125),
.B1(n_3122),
.B2(n_3123),
.Y(n_15052)
);

OAI221xp5_ASAP7_75t_L g15053 ( 
.A1(n_15027),
.A2(n_3128),
.B1(n_3126),
.B2(n_3127),
.C(n_3129),
.Y(n_15053)
);

NAND2xp5_ASAP7_75t_L g15054 ( 
.A(n_15040),
.B(n_15036),
.Y(n_15054)
);

INVx2_ASAP7_75t_L g15055 ( 
.A(n_15042),
.Y(n_15055)
);

INVx1_ASAP7_75t_L g15056 ( 
.A(n_15039),
.Y(n_15056)
);

AOI21xp5_ASAP7_75t_L g15057 ( 
.A1(n_15046),
.A2(n_15023),
.B(n_15022),
.Y(n_15057)
);

OR2x6_ASAP7_75t_L g15058 ( 
.A(n_15044),
.B(n_15021),
.Y(n_15058)
);

AOI22xp5_ASAP7_75t_L g15059 ( 
.A1(n_15048),
.A2(n_15035),
.B1(n_3130),
.B2(n_3131),
.Y(n_15059)
);

INVx2_ASAP7_75t_L g15060 ( 
.A(n_15041),
.Y(n_15060)
);

INVx1_ASAP7_75t_L g15061 ( 
.A(n_15051),
.Y(n_15061)
);

AOI21xp5_ASAP7_75t_L g15062 ( 
.A1(n_15047),
.A2(n_15035),
.B(n_3126),
.Y(n_15062)
);

AO22x2_ASAP7_75t_L g15063 ( 
.A1(n_15043),
.A2(n_3131),
.B1(n_3127),
.B2(n_3130),
.Y(n_15063)
);

INVx4_ASAP7_75t_L g15064 ( 
.A(n_15050),
.Y(n_15064)
);

XNOR2xp5_ASAP7_75t_L g15065 ( 
.A(n_15049),
.B(n_3134),
.Y(n_15065)
);

NAND2xp5_ASAP7_75t_L g15066 ( 
.A(n_15045),
.B(n_3136),
.Y(n_15066)
);

AOI21xp33_ASAP7_75t_L g15067 ( 
.A1(n_15053),
.A2(n_3135),
.B(n_3136),
.Y(n_15067)
);

AOI21xp5_ASAP7_75t_L g15068 ( 
.A1(n_15052),
.A2(n_3135),
.B(n_3137),
.Y(n_15068)
);

OAI221xp5_ASAP7_75t_L g15069 ( 
.A1(n_15059),
.A2(n_3139),
.B1(n_3137),
.B2(n_3138),
.C(n_3140),
.Y(n_15069)
);

AND2x4_ASAP7_75t_L g15070 ( 
.A(n_15055),
.B(n_3138),
.Y(n_15070)
);

CKINVDCx20_ASAP7_75t_R g15071 ( 
.A(n_15056),
.Y(n_15071)
);

AOI22xp33_ASAP7_75t_L g15072 ( 
.A1(n_15067),
.A2(n_3142),
.B1(n_3139),
.B2(n_3141),
.Y(n_15072)
);

AOI22xp5_ASAP7_75t_L g15073 ( 
.A1(n_15066),
.A2(n_3143),
.B1(n_3141),
.B2(n_3142),
.Y(n_15073)
);

AOI22xp5_ASAP7_75t_L g15074 ( 
.A1(n_15061),
.A2(n_3145),
.B1(n_3143),
.B2(n_3144),
.Y(n_15074)
);

NOR2xp67_ASAP7_75t_L g15075 ( 
.A(n_15064),
.B(n_3144),
.Y(n_15075)
);

INVx1_ASAP7_75t_L g15076 ( 
.A(n_15065),
.Y(n_15076)
);

AOI22xp33_ASAP7_75t_L g15077 ( 
.A1(n_15060),
.A2(n_3147),
.B1(n_3145),
.B2(n_3146),
.Y(n_15077)
);

CKINVDCx20_ASAP7_75t_R g15078 ( 
.A(n_15054),
.Y(n_15078)
);

INVx1_ASAP7_75t_L g15079 ( 
.A(n_15058),
.Y(n_15079)
);

INVx2_ASAP7_75t_L g15080 ( 
.A(n_15063),
.Y(n_15080)
);

HB1xp67_ASAP7_75t_L g15081 ( 
.A(n_15079),
.Y(n_15081)
);

BUFx2_ASAP7_75t_L g15082 ( 
.A(n_15071),
.Y(n_15082)
);

INVx4_ASAP7_75t_L g15083 ( 
.A(n_15080),
.Y(n_15083)
);

INVx2_ASAP7_75t_L g15084 ( 
.A(n_15078),
.Y(n_15084)
);

BUFx2_ASAP7_75t_L g15085 ( 
.A(n_15076),
.Y(n_15085)
);

INVx1_ASAP7_75t_L g15086 ( 
.A(n_15075),
.Y(n_15086)
);

OAI22xp5_ASAP7_75t_L g15087 ( 
.A1(n_15072),
.A2(n_15058),
.B1(n_15057),
.B2(n_15062),
.Y(n_15087)
);

INVx1_ASAP7_75t_L g15088 ( 
.A(n_15081),
.Y(n_15088)
);

HB1xp67_ASAP7_75t_L g15089 ( 
.A(n_15082),
.Y(n_15089)
);

INVx1_ASAP7_75t_L g15090 ( 
.A(n_15084),
.Y(n_15090)
);

INVx1_ASAP7_75t_L g15091 ( 
.A(n_15086),
.Y(n_15091)
);

AOI22xp5_ASAP7_75t_L g15092 ( 
.A1(n_15088),
.A2(n_15083),
.B1(n_15085),
.B2(n_15087),
.Y(n_15092)
);

AOI22xp5_ASAP7_75t_L g15093 ( 
.A1(n_15089),
.A2(n_15068),
.B1(n_15069),
.B2(n_15073),
.Y(n_15093)
);

AOI22xp5_ASAP7_75t_L g15094 ( 
.A1(n_15092),
.A2(n_15090),
.B1(n_15091),
.B2(n_15074),
.Y(n_15094)
);

AOI22xp5_ASAP7_75t_L g15095 ( 
.A1(n_15093),
.A2(n_15077),
.B1(n_15070),
.B2(n_3148),
.Y(n_15095)
);

OAI21xp5_ASAP7_75t_L g15096 ( 
.A1(n_15094),
.A2(n_3146),
.B(n_3147),
.Y(n_15096)
);

NAND2xp33_ASAP7_75t_L g15097 ( 
.A(n_15095),
.B(n_3148),
.Y(n_15097)
);

AOI222xp33_ASAP7_75t_L g15098 ( 
.A1(n_15097),
.A2(n_3151),
.B1(n_3154),
.B2(n_3149),
.C1(n_3150),
.C2(n_3152),
.Y(n_15098)
);

AOI21xp5_ASAP7_75t_L g15099 ( 
.A1(n_15098),
.A2(n_15096),
.B(n_3151),
.Y(n_15099)
);

AOI22xp5_ASAP7_75t_L g15100 ( 
.A1(n_15099),
.A2(n_3154),
.B1(n_3149),
.B2(n_3150),
.Y(n_15100)
);

AOI31xp33_ASAP7_75t_L g15101 ( 
.A1(n_15099),
.A2(n_3157),
.A3(n_3155),
.B(n_3156),
.Y(n_15101)
);

AOI22xp33_ASAP7_75t_L g15102 ( 
.A1(n_15100),
.A2(n_3159),
.B1(n_3156),
.B2(n_3158),
.Y(n_15102)
);

AOI211xp5_ASAP7_75t_L g15103 ( 
.A1(n_15102),
.A2(n_15101),
.B(n_3160),
.C(n_3158),
.Y(n_15103)
);


endmodule