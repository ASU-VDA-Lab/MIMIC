module real_aes_681_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_0), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_1), .B(n_133), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_2), .A2(n_141), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_3), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_4), .B(n_133), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_5), .B(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_6), .B(n_160), .Y(n_491) );
INVx1_ASAP7_75t_L g129 ( .A(n_7), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_8), .B(n_160), .Y(n_540) );
CKINVDCx16_ASAP7_75t_R g786 ( .A(n_9), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_10), .A2(n_14), .B1(n_769), .B2(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_10), .Y(n_769) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_11), .B(n_158), .Y(n_532) );
AND2x2_ASAP7_75t_L g163 ( .A(n_12), .B(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g174 ( .A(n_13), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_14), .Y(n_770) );
INVx2_ASAP7_75t_L g120 ( .A(n_15), .Y(n_120) );
AOI221x1_ASAP7_75t_L g476 ( .A1(n_16), .A2(n_28), .B1(n_133), .B2(n_141), .C(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_17), .A2(n_767), .B1(n_772), .B2(n_773), .Y(n_766) );
INVx1_ASAP7_75t_L g772 ( .A(n_17), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_18), .B(n_160), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_19), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_19), .B(n_785), .C(n_787), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_20), .B(n_133), .Y(n_528) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_21), .A2(n_175), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_22), .B(n_118), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_23), .B(n_160), .Y(n_465) );
AO21x1_ASAP7_75t_L g486 ( .A1(n_24), .A2(n_133), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_25), .B(n_133), .Y(n_216) );
INVx1_ASAP7_75t_L g444 ( .A(n_26), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_27), .A2(n_92), .B1(n_124), .B2(n_133), .Y(n_123) );
NAND2x1_ASAP7_75t_L g507 ( .A(n_29), .B(n_160), .Y(n_507) );
NAND2x1_ASAP7_75t_L g539 ( .A(n_30), .B(n_158), .Y(n_539) );
OR2x2_ASAP7_75t_L g121 ( .A(n_31), .B(n_89), .Y(n_121) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_31), .A2(n_89), .B(n_120), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_32), .B(n_158), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_33), .B(n_160), .Y(n_531) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_34), .A2(n_164), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_35), .B(n_158), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_36), .A2(n_141), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_37), .B(n_160), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_38), .A2(n_141), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g131 ( .A(n_39), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g139 ( .A(n_39), .B(n_129), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_39), .Y(n_145) );
OR2x6_ASAP7_75t_L g442 ( .A(n_40), .B(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g787 ( .A(n_40), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_41), .B(n_133), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_42), .B(n_133), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_43), .B(n_160), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_44), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_45), .B(n_158), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_46), .B(n_133), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_47), .A2(n_141), .B(n_156), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_48), .A2(n_104), .B1(n_779), .B2(n_788), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_49), .A2(n_743), .B1(n_744), .B2(n_747), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_49), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_50), .A2(n_141), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_51), .B(n_158), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_52), .B(n_158), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_53), .B(n_133), .Y(n_197) );
INVx1_ASAP7_75t_L g127 ( .A(n_54), .Y(n_127) );
INVx1_ASAP7_75t_L g136 ( .A(n_54), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_55), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g206 ( .A(n_56), .B(n_118), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_57), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_58), .B(n_160), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_59), .B(n_158), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_60), .A2(n_141), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_61), .B(n_133), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_62), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_63), .B(n_133), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_64), .A2(n_141), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g222 ( .A(n_65), .B(n_119), .Y(n_222) );
AO21x1_ASAP7_75t_L g488 ( .A1(n_66), .A2(n_141), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_67), .B(n_133), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_68), .B(n_158), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_69), .B(n_133), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_70), .B(n_158), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_71), .A2(n_96), .B1(n_141), .B2(n_143), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_72), .B(n_160), .Y(n_219) );
AND2x2_ASAP7_75t_L g501 ( .A(n_73), .B(n_119), .Y(n_501) );
INVx1_ASAP7_75t_L g132 ( .A(n_74), .Y(n_132) );
INVx1_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
AND2x2_ASAP7_75t_L g542 ( .A(n_75), .B(n_164), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_76), .B(n_158), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_77), .A2(n_141), .B(n_210), .Y(n_209) );
AOI22xp5_ASAP7_75t_SL g744 ( .A1(n_78), .A2(n_83), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_78), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_79), .A2(n_141), .B(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_80), .A2(n_141), .B(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g232 ( .A(n_81), .B(n_119), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_82), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g745 ( .A(n_83), .Y(n_745) );
INVx1_ASAP7_75t_L g445 ( .A(n_84), .Y(n_445) );
AND2x2_ASAP7_75t_L g453 ( .A(n_85), .B(n_164), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_86), .B(n_133), .Y(n_467) );
AND2x2_ASAP7_75t_L g187 ( .A(n_87), .B(n_175), .Y(n_187) );
AND2x2_ASAP7_75t_L g487 ( .A(n_88), .B(n_202), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_90), .B(n_158), .Y(n_466) );
AND2x2_ASAP7_75t_L g510 ( .A(n_91), .B(n_164), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_93), .B(n_160), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_94), .A2(n_141), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_95), .B(n_158), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_97), .A2(n_141), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_98), .B(n_160), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_99), .B(n_160), .Y(n_458) );
BUFx2_ASAP7_75t_L g221 ( .A(n_100), .Y(n_221) );
BUFx2_ASAP7_75t_L g762 ( .A(n_101), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_102), .A2(n_141), .B(n_530), .Y(n_529) );
AO221x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_758), .B1(n_763), .B2(n_766), .C(n_774), .Y(n_104) );
OAI222xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_742), .B1(n_748), .B2(n_749), .C1(n_754), .C2(n_757), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_437), .B1(n_446), .B2(n_738), .Y(n_107) );
INVx3_ASAP7_75t_L g751 ( .A(n_108), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_108), .A2(n_751), .B1(n_768), .B2(n_771), .Y(n_767) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_362), .Y(n_108) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_298), .C(n_345), .Y(n_109) );
NAND4xp25_ASAP7_75t_SL g110 ( .A(n_111), .B(n_233), .C(n_251), .D(n_277), .Y(n_110) );
OAI21xp33_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_191), .B(n_192), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g112 ( .A(n_113), .B(n_176), .Y(n_112) );
INVx1_ASAP7_75t_L g413 ( .A(n_113), .Y(n_413) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_148), .Y(n_113) );
INVx2_ASAP7_75t_L g237 ( .A(n_114), .Y(n_237) );
AND2x2_ASAP7_75t_L g257 ( .A(n_114), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g359 ( .A(n_114), .B(n_178), .Y(n_359) );
AND2x2_ASAP7_75t_L g419 ( .A(n_114), .B(n_238), .Y(n_419) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_115), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g303 ( .A(n_116), .B(n_151), .Y(n_303) );
BUFx3_ASAP7_75t_L g313 ( .A(n_116), .Y(n_313) );
AND2x2_ASAP7_75t_L g376 ( .A(n_116), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_122), .Y(n_116) );
AND2x4_ASAP7_75t_L g190 ( .A(n_117), .B(n_122), .Y(n_190) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_118), .A2(n_123), .B(n_140), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_118), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_118), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_118), .A2(n_455), .B(n_456), .Y(n_454) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_118), .A2(n_476), .B(n_480), .Y(n_475) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_118), .A2(n_476), .B(n_480), .Y(n_546) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x4_ASAP7_75t_L g202 ( .A(n_120), .B(n_121), .Y(n_202) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_130), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g142 ( .A(n_127), .B(n_129), .Y(n_142) );
AND2x4_ASAP7_75t_L g160 ( .A(n_127), .B(n_137), .Y(n_160) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x6_ASAP7_75t_L g141 ( .A(n_131), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g147 ( .A(n_132), .Y(n_147) );
AND2x6_ASAP7_75t_L g158 ( .A(n_132), .B(n_135), .Y(n_158) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx5_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
AND2x4_ASAP7_75t_L g143 ( .A(n_142), .B(n_144), .Y(n_143) );
NOR2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g422 ( .A(n_149), .Y(n_422) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_165), .Y(n_149) );
AND2x2_ASAP7_75t_L g189 ( .A(n_150), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g377 ( .A(n_150), .Y(n_377) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g191 ( .A(n_151), .B(n_180), .Y(n_191) );
AND2x2_ASAP7_75t_L g254 ( .A(n_151), .B(n_165), .Y(n_254) );
INVx2_ASAP7_75t_L g259 ( .A(n_151), .Y(n_259) );
AND2x2_ASAP7_75t_L g261 ( .A(n_151), .B(n_166), .Y(n_261) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_163), .Y(n_151) );
INVx4_ASAP7_75t_L g164 ( .A(n_152), .Y(n_164) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_162), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_158), .B(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_161), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_161), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_161), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_161), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_161), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_161), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_161), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_161), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_161), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_161), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_161), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_161), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_539), .B(n_540), .Y(n_538) );
INVx3_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
INVx1_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
INVx2_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
AND2x4_ASAP7_75t_SL g274 ( .A(n_165), .B(n_180), .Y(n_274) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_165), .Y(n_306) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_174), .Y(n_166) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_167), .A2(n_536), .B(n_542), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_173), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_175), .A2(n_216), .B(n_217), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_189), .Y(n_176) );
AND2x2_ASAP7_75t_L g340 ( .A(n_177), .B(n_285), .Y(n_340) );
INVx2_ASAP7_75t_SL g428 ( .A(n_177), .Y(n_428) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_188), .Y(n_178) );
NAND2x1p5_ASAP7_75t_L g241 ( .A(n_179), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g348 ( .A(n_179), .B(n_261), .Y(n_348) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g236 ( .A(n_180), .Y(n_236) );
AND2x4_ASAP7_75t_L g238 ( .A(n_180), .B(n_239), .Y(n_238) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_180), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g331 ( .A(n_180), .Y(n_331) );
AND2x2_ASAP7_75t_L g350 ( .A(n_180), .B(n_289), .Y(n_350) );
AND2x2_ASAP7_75t_L g381 ( .A(n_180), .B(n_290), .Y(n_381) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_187), .Y(n_180) );
AND2x2_ASAP7_75t_L g320 ( .A(n_189), .B(n_274), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_189), .B(n_331), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_189), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
AND2x2_ASAP7_75t_L g433 ( .A(n_189), .B(n_240), .Y(n_433) );
INVx3_ASAP7_75t_L g286 ( .A(n_190), .Y(n_286) );
AND2x2_ASAP7_75t_L g289 ( .A(n_190), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_191), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g314 ( .A(n_191), .Y(n_314) );
AND2x4_ASAP7_75t_SL g192 ( .A(n_193), .B(n_203), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_193), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g365 ( .A(n_193), .B(n_366), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_193), .B(n_327), .C(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g435 ( .A(n_193), .B(n_329), .Y(n_435) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g250 ( .A(n_195), .B(n_214), .Y(n_250) );
INVx1_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
INVx2_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_195), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_195), .B(n_282), .Y(n_309) );
AND2x2_ASAP7_75t_L g388 ( .A(n_195), .B(n_205), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_202), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_202), .A2(n_208), .B(n_209), .Y(n_207) );
INVx1_ASAP7_75t_SL g461 ( .A(n_202), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_202), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_202), .A2(n_528), .B(n_529), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_203), .A2(n_252), .B1(n_255), .B2(n_262), .C(n_268), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_203), .A2(n_381), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
INVx2_ASAP7_75t_L g322 ( .A(n_204), .Y(n_322) );
AND2x2_ASAP7_75t_L g382 ( .A(n_204), .B(n_266), .Y(n_382) );
AND2x2_ASAP7_75t_L g392 ( .A(n_204), .B(n_278), .Y(n_392) );
OR2x2_ASAP7_75t_L g432 ( .A(n_204), .B(n_316), .Y(n_432) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_SL g249 ( .A(n_205), .B(n_250), .Y(n_249) );
NAND2x1_ASAP7_75t_L g265 ( .A(n_205), .B(n_214), .Y(n_265) );
INVx4_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
OR2x2_ASAP7_75t_L g336 ( .A(n_205), .B(n_223), .Y(n_336) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x2_ASAP7_75t_L g387 ( .A(n_213), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
INVx2_ASAP7_75t_SL g275 ( .A(n_214), .Y(n_275) );
NOR2x1_ASAP7_75t_SL g281 ( .A(n_214), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g296 ( .A(n_214), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g327 ( .A(n_214), .B(n_294), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_214), .B(n_280), .Y(n_334) );
BUFx2_ASAP7_75t_L g368 ( .A(n_214), .Y(n_368) );
AND2x2_ASAP7_75t_L g379 ( .A(n_214), .B(n_294), .Y(n_379) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_222), .Y(n_214) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_223), .Y(n_247) );
AND2x2_ASAP7_75t_L g266 ( .A(n_223), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g297 ( .A(n_223), .Y(n_297) );
AND2x2_ASAP7_75t_L g323 ( .A(n_223), .B(n_279), .Y(n_323) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
AO21x1_ASAP7_75t_SL g282 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_282) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_225), .A2(n_495), .B(n_501), .Y(n_494) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_225), .A2(n_504), .B(n_510), .Y(n_503) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_225), .A2(n_504), .B(n_510), .Y(n_516) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_225), .A2(n_495), .B(n_501), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
OAI31xp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_238), .A3(n_240), .B(n_244), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g342 ( .A(n_236), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_237), .A2(n_326), .A3(n_333), .B1(n_337), .B2(n_338), .C1(n_340), .C2(n_341), .Y(n_332) );
AND2x2_ASAP7_75t_L g404 ( .A(n_237), .B(n_381), .Y(n_404) );
AOI221xp5_ASAP7_75t_SL g317 ( .A1(n_238), .A2(n_318), .B1(n_320), .B2(n_321), .C(n_324), .Y(n_317) );
INVx2_ASAP7_75t_L g337 ( .A(n_238), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_240), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_240), .B(n_333), .Y(n_436) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g311 ( .A(n_241), .B(n_286), .Y(n_311) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g290 ( .A(n_243), .B(n_259), .Y(n_290) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g361 ( .A(n_247), .Y(n_361) );
O2A1O1Ixp5_ASAP7_75t_L g352 ( .A1(n_248), .A2(n_353), .B(n_355), .C(n_357), .Y(n_352) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_249), .A2(n_385), .B1(n_386), .B2(n_389), .Y(n_384) );
OR2x2_ASAP7_75t_L g339 ( .A(n_250), .B(n_336), .Y(n_339) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_256), .B(n_260), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g272 ( .A(n_259), .Y(n_272) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_261), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g315 ( .A(n_265), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_265), .B(n_266), .Y(n_358) );
OR2x2_ASAP7_75t_L g360 ( .A(n_265), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_265), .B(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
NOR4xp25_ASAP7_75t_L g268 ( .A(n_269), .B(n_273), .C(n_275), .D(n_276), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g396 ( .A(n_270), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g424 ( .A(n_270), .B(n_273), .Y(n_424) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g354 ( .A(n_272), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_273), .B(n_302), .Y(n_389) );
AOI321xp33_ASAP7_75t_L g391 ( .A1(n_273), .A2(n_392), .A3(n_393), .B1(n_394), .B2(n_396), .C(n_399), .Y(n_391) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_SL g353 ( .A(n_274), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_274), .B(n_313), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_275), .B(n_297), .Y(n_402) );
OR2x2_ASAP7_75t_L g429 ( .A(n_276), .B(n_313), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_283), .B(n_287), .Y(n_277) );
AND2x2_ASAP7_75t_L g318 ( .A(n_278), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g344 ( .A(n_280), .B(n_282), .Y(n_344) );
INVx2_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_284), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g385 ( .A(n_285), .B(n_337), .Y(n_385) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g343 ( .A(n_286), .B(n_344), .Y(n_343) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_286), .B(n_422), .Y(n_421) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g372 ( .A(n_290), .Y(n_372) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_294), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
BUFx2_ASAP7_75t_L g401 ( .A(n_294), .Y(n_401) );
INVxp67_ASAP7_75t_L g409 ( .A(n_297), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_317), .C(n_332), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_307), .B(n_310), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g330 ( .A(n_303), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g383 ( .A(n_304), .Y(n_383) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g398 ( .A(n_306), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_307), .A2(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g316 ( .A(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g378 ( .A(n_309), .B(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_315), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_311), .A2(n_358), .B1(n_359), .B2(n_360), .Y(n_357) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
OR2x2_ASAP7_75t_L g395 ( .A(n_316), .B(n_327), .Y(n_395) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_319), .B(n_368), .C(n_428), .D(n_429), .Y(n_427) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
OR2x2_ASAP7_75t_L g328 ( .A(n_322), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_322), .B(n_344), .Y(n_426) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_328), .B(n_330), .Y(n_324) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g415 ( .A(n_327), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g423 ( .A(n_329), .Y(n_423) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVxp67_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g367 ( .A(n_336), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g416 ( .A(n_344), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B(n_351), .C(n_352), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_390), .C(n_411), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_369), .B(n_373), .C(n_380), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g412 ( .A1(n_376), .A2(n_413), .B(n_414), .C(n_417), .Y(n_412) );
BUFx2_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .Y(n_390) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_400), .A2(n_406), .B1(n_407), .B2(n_410), .Y(n_405) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_412), .B(n_420), .C(n_430), .D(n_436), .Y(n_411) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_424), .B2(n_425), .C(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx6p67_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_439), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
AND2x6_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OR2x6_ASAP7_75t_SL g740 ( .A(n_441), .B(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g756 ( .A(n_441), .B(n_442), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_441), .B(n_741), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_442), .Y(n_741) );
INVx1_ASAP7_75t_L g783 ( .A(n_443), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx3_ASAP7_75t_SL g753 ( .A(n_446), .Y(n_753) );
NOR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_625), .Y(n_446) );
AO211x2_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_470), .B(n_520), .C(n_593), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AND3x2_ASAP7_75t_L g674 ( .A(n_450), .B(n_555), .C(n_571), .Y(n_674) );
AND2x4_ASAP7_75t_L g677 ( .A(n_450), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_451), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g586 ( .A(n_451), .Y(n_586) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_451), .B(n_580), .Y(n_671) );
AND2x2_ASAP7_75t_L g714 ( .A(n_451), .B(n_535), .Y(n_714) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g563 ( .A(n_452), .Y(n_563) );
AND2x2_ASAP7_75t_L g582 ( .A(n_452), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_452), .B(n_535), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_452), .B(n_534), .Y(n_660) );
NOR2x1_ASAP7_75t_SL g687 ( .A(n_452), .B(n_460), .Y(n_687) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_460), .B(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_468), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_461), .B(n_469), .Y(n_468) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_461), .A2(n_462), .B(n_468), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
AO21x1_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_502), .B(n_511), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_472), .A2(n_569), .B1(n_573), .B2(n_574), .Y(n_568) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
AND2x2_ASAP7_75t_L g629 ( .A(n_473), .B(n_517), .Y(n_629) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g562 ( .A(n_474), .B(n_545), .Y(n_562) );
AND2x2_ASAP7_75t_L g634 ( .A(n_474), .B(n_519), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_474), .B(n_619), .Y(n_653) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_475), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_481), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g613 ( .A(n_482), .B(n_514), .Y(n_613) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
AND2x2_ASAP7_75t_L g517 ( .A(n_483), .B(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g550 ( .A(n_483), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_483), .B(n_546), .Y(n_610) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g703 ( .A(n_484), .Y(n_703) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g545 ( .A(n_485), .Y(n_545) );
OAI21x1_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_488), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g493 ( .A(n_487), .Y(n_493) );
INVx2_ASAP7_75t_L g551 ( .A(n_494), .Y(n_551) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_494), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_500), .Y(n_495) );
INVx2_ASAP7_75t_L g547 ( .A(n_502), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_502), .B(n_679), .Y(n_705) );
AND2x2_ASAP7_75t_L g724 ( .A(n_502), .B(n_714), .Y(n_724) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_503), .B(n_551), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_512), .B(n_561), .Y(n_596) );
INVx1_ASAP7_75t_SL g723 ( .A(n_512), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_513), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
AND2x2_ASAP7_75t_L g735 ( .A(n_514), .B(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g611 ( .A(n_515), .B(n_518), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_515), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g665 ( .A(n_515), .B(n_519), .Y(n_665) );
AND2x2_ASAP7_75t_L g696 ( .A(n_515), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g561 ( .A(n_516), .B(n_519), .Y(n_561) );
INVxp67_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
BUFx3_ASAP7_75t_L g619 ( .A(n_516), .Y(n_619) );
AND2x2_ASAP7_75t_L g639 ( .A(n_517), .B(n_640), .Y(n_639) );
NAND2xp33_ASAP7_75t_L g652 ( .A(n_517), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_518), .B(n_545), .Y(n_608) );
AND2x2_ASAP7_75t_L g697 ( .A(n_518), .B(n_546), .Y(n_697) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g624 ( .A(n_519), .B(n_546), .Y(n_624) );
OR3x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_568), .C(n_583), .Y(n_520) );
OAI321xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_533), .A3(n_543), .B1(n_548), .B2(n_552), .C(n_560), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_525), .Y(n_599) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_525), .Y(n_617) );
OR2x2_ASAP7_75t_L g621 ( .A(n_525), .B(n_533), .Y(n_621) );
BUFx3_ASAP7_75t_L g555 ( .A(n_526), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_558), .Y(n_572) );
INVx1_ASAP7_75t_L g589 ( .A(n_526), .Y(n_589) );
INVx2_ASAP7_75t_L g605 ( .A(n_526), .Y(n_605) );
OR2x2_ASAP7_75t_L g644 ( .A(n_526), .B(n_534), .Y(n_644) );
INVx2_ASAP7_75t_L g632 ( .A(n_533), .Y(n_632) );
AND2x2_ASAP7_75t_L g556 ( .A(n_534), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g571 ( .A(n_534), .Y(n_571) );
AND2x4_ASAP7_75t_L g580 ( .A(n_534), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_534), .B(n_557), .Y(n_603) );
AND2x2_ASAP7_75t_L g710 ( .A(n_534), .B(n_605), .Y(n_710) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_535), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g597 ( .A(n_543), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_547), .Y(n_543) );
AND2x2_ASAP7_75t_L g684 ( .A(n_544), .B(n_611), .Y(n_684) );
INVx1_ASAP7_75t_SL g701 ( .A(n_544), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_544), .B(n_677), .Y(n_730) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OR2x2_ASAP7_75t_L g573 ( .A(n_545), .B(n_546), .Y(n_573) );
AND2x2_ASAP7_75t_L g666 ( .A(n_547), .B(n_562), .Y(n_666) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_551), .B(n_562), .Y(n_689) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_553), .A2(n_702), .B1(n_707), .B2(n_709), .Y(n_706) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g631 ( .A(n_554), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g726 ( .A(n_554), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g682 ( .A(n_555), .B(n_600), .Y(n_682) );
AND2x4_ASAP7_75t_L g636 ( .A(n_556), .B(n_582), .Y(n_636) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_558), .Y(n_734) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g567 ( .A(n_559), .Y(n_567) );
INVx1_ASAP7_75t_L g581 ( .A(n_559), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .D(n_564), .Y(n_560) );
AND2x2_ASAP7_75t_L g718 ( .A(n_561), .B(n_703), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_561), .B(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_562), .B(n_638), .Y(n_637) );
OAI322xp33_ASAP7_75t_L g645 ( .A1(n_562), .A2(n_646), .A3(n_650), .B1(n_652), .B2(n_654), .C1(n_656), .C2(n_661), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_562), .B(n_611), .Y(n_661) );
INVx1_ASAP7_75t_L g729 ( .A(n_562), .Y(n_729) );
INVx2_ASAP7_75t_L g575 ( .A(n_563), .Y(n_575) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_566), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_567), .B(n_586), .Y(n_643) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_570), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g616 ( .A(n_571), .Y(n_616) );
AND2x2_ASAP7_75t_L g688 ( .A(n_571), .B(n_599), .Y(n_688) );
AOI31xp33_ASAP7_75t_L g574 ( .A1(n_572), .A2(n_575), .A3(n_576), .B(n_579), .Y(n_574) );
AND2x2_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g713 ( .A(n_572), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_572), .B(n_600), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_572), .Y(n_721) );
INVx1_ASAP7_75t_SL g679 ( .A(n_573), .Y(n_679) );
NAND3xp33_ASAP7_75t_SL g707 ( .A(n_573), .B(n_701), .C(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g607 ( .A(n_578), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g588 ( .A(n_580), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g649 ( .A(n_580), .Y(n_649) );
AOI322xp5_ASAP7_75t_L g731 ( .A1(n_580), .A2(n_610), .A3(n_613), .B1(n_732), .B2(n_733), .C1(n_735), .C2(n_737), .Y(n_731) );
AND2x2_ASAP7_75t_L g737 ( .A(n_580), .B(n_586), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B(n_590), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_586), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g732 ( .A(n_586), .B(n_619), .Y(n_732) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
AND2x2_ASAP7_75t_L g686 ( .A(n_589), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g733 ( .A(n_589), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g638 ( .A(n_592), .Y(n_638) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
O2A1O1Ixp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_598), .C(n_601), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g655 ( .A(n_600), .B(n_605), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .B(n_612), .C(n_614), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_602), .A2(n_628), .B1(n_630), .B2(n_633), .C(n_635), .Y(n_627) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g647 ( .A(n_604), .Y(n_647) );
OR2x2_ASAP7_75t_L g667 ( .A(n_604), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g712 ( .A(n_607), .Y(n_712) );
INVx1_ASAP7_75t_L g736 ( .A(n_608), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_610), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_610), .B(n_680), .Y(n_692) );
INVx1_ASAP7_75t_L g672 ( .A(n_611), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B1(n_620), .B2(n_622), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_SL g680 ( .A(n_619), .Y(n_680) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND4xp75_ASAP7_75t_L g625 ( .A(n_626), .B(n_662), .C(n_690), .D(n_715), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_627), .B(n_645), .Y(n_626) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_634), .B(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_639), .B2(n_641), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_638), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
OR2x2_ASAP7_75t_L g693 ( .A(n_644), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g708 ( .A(n_653), .Y(n_708) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g699 ( .A1(n_655), .A2(n_700), .B(n_702), .Y(n_699) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_675), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_667), .B1(n_670), .B2(n_672), .C(n_673), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g711 ( .A1(n_665), .A2(n_712), .B(n_713), .Y(n_711) );
INVx3_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .A3(n_680), .B1(n_681), .B2(n_683), .C1(n_685), .C2(n_689), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g698 ( .A(n_686), .Y(n_698) );
INVx1_ASAP7_75t_L g694 ( .A(n_687), .Y(n_694) );
AND2x2_ASAP7_75t_L g709 ( .A(n_687), .B(n_710), .Y(n_709) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_704), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_698), .C(n_699), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_698), .A2(n_705), .B(n_706), .C(n_711), .Y(n_704) );
INVx2_ASAP7_75t_SL g727 ( .A(n_714), .Y(n_727) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_725), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_721), .B2(n_722), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_728), .B(n_730), .C(n_731), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g752 ( .A(n_739), .Y(n_752) );
CKINVDCx11_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
CKINVDCx12_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
BUFx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2x1_ASAP7_75t_R g763 ( .A(n_762), .B(n_764), .Y(n_763) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_R g778 ( .A(n_765), .Y(n_778) );
INVx1_ASAP7_75t_L g773 ( .A(n_767), .Y(n_773) );
INVx1_ASAP7_75t_L g771 ( .A(n_768), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVxp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g789 ( .A(n_781), .Y(n_789) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_SL g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
endmodule