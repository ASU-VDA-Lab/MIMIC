module fake_jpeg_29362_n_361 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_361);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_51),
.B(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_23),
.B(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_24),
.B1(n_29),
.B2(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_43),
.B1(n_17),
.B2(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx3_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_67),
.Y(n_125)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_12),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_12),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_74),
.Y(n_126)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_78),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_11),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_81),
.Y(n_133)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_82),
.Y(n_122)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_85),
.B1(n_32),
.B2(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_97),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_42),
.B1(n_18),
.B2(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_89),
.A2(n_91),
.B1(n_95),
.B2(n_100),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_42),
.B1(n_18),
.B2(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_114),
.B1(n_120),
.B2(n_124),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_31),
.B1(n_38),
.B2(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_22),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_22),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_101),
.B(n_103),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_37),
.B1(n_34),
.B2(n_26),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_109),
.A2(n_111),
.B1(n_121),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_28),
.B1(n_30),
.B2(n_39),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_16),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_127),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_44),
.B1(n_39),
.B2(n_20),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_59),
.B(n_44),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_0),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_85),
.B1(n_68),
.B2(n_78),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_28),
.B1(n_22),
.B2(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_22),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_40),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_0),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_40),
.B1(n_11),
.B2(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_54),
.A2(n_40),
.B1(n_9),
.B2(n_21),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_75),
.B1(n_66),
.B2(n_81),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_151),
.B1(n_153),
.B2(n_130),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_59),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g201 ( 
.A(n_143),
.B(n_117),
.C(n_94),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_150),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_40),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_0),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_5),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_175),
.B1(n_130),
.B2(n_94),
.Y(n_187)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_7),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_173),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_7),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_8),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_8),
.B(n_97),
.C(n_87),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_87),
.B(n_8),
.Y(n_176)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_102),
.B1(n_92),
.B2(n_90),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_180),
.B1(n_194),
.B2(n_209),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_102),
.B1(n_92),
.B2(n_90),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_130),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_183),
.B(n_185),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_88),
.CI(n_129),
.CON(n_185),
.SN(n_185)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_192),
.B1(n_205),
.B2(n_175),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_87),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_197),
.C(n_144),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_140),
.A2(n_170),
.B1(n_157),
.B2(n_138),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_136),
.B1(n_99),
.B2(n_112),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_113),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_189),
.B(n_204),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_138),
.B(n_170),
.CI(n_140),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_8),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_157),
.B1(n_160),
.B2(n_149),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_150),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_153),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_221),
.C(n_206),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_167),
.B1(n_175),
.B2(n_142),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_223),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_175),
.B1(n_171),
.B2(n_155),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_204),
.B1(n_210),
.B2(n_199),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_205),
.B1(n_207),
.B2(n_201),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_226),
.B(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_163),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_127),
.C(n_103),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_165),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_223),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_175),
.B1(n_171),
.B2(n_141),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_232),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_228),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_94),
.B1(n_105),
.B2(n_145),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_105),
.B(n_110),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_234),
.B(n_188),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_230),
.Y(n_262)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_231),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_177),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_236),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_139),
.B(n_166),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_152),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_182),
.B(n_110),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_259),
.B1(n_223),
.B2(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_260),
.C(n_261),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_216),
.B1(n_234),
.B2(n_240),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_256),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_237),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_182),
.B(n_181),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_199),
.B1(n_184),
.B2(n_190),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_184),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_196),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_190),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_234),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_193),
.C(n_115),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_229),
.C(n_232),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_164),
.C(n_196),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_219),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_245),
.B1(n_247),
.B2(n_234),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_246),
.B(n_220),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_269),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_273),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_271),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_212),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_228),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_278),
.C(n_273),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_227),
.C(n_225),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_259),
.B1(n_241),
.B2(n_249),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_283),
.B1(n_285),
.B2(n_262),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_262),
.B1(n_230),
.B2(n_258),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_231),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_236),
.Y(n_300)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_256),
.Y(n_286)
);

OAI322xp33_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_257),
.A3(n_250),
.B1(n_251),
.B2(n_265),
.C1(n_253),
.C2(n_261),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_298),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_250),
.B(n_284),
.C(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_255),
.C(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_299),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_244),
.C(n_264),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_304),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_254),
.C(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_282),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_230),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_243),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_272),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_208),
.C(n_235),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_286),
.B(n_269),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_306),
.B(n_316),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_266),
.B(n_279),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_272),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_288),
.B(n_281),
.CI(n_280),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_314),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_270),
.B(n_282),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_317),
.A2(n_300),
.B1(n_200),
.B2(n_191),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_154),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_292),
.C(n_296),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_289),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_323),
.C(n_324),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_316),
.B1(n_306),
.B2(n_293),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_313),
.B1(n_311),
.B2(n_310),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_298),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_287),
.B1(n_291),
.B2(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_331),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_191),
.B1(n_115),
.B2(n_193),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_330),
.A2(n_318),
.B(n_317),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_340),
.B(n_334),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_324),
.B1(n_320),
.B2(n_321),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_328),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_323),
.A2(n_313),
.B(n_319),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_99),
.C(n_136),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_320),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_347),
.Y(n_352)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_339),
.A2(n_333),
.B(n_336),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_345),
.A2(n_166),
.B(n_137),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_346),
.B(n_348),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_341),
.B(n_332),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_336),
.A2(n_159),
.B1(n_147),
.B2(n_137),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_112),
.C(n_117),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_350),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_355),
.Y(n_358)
);

AOI322xp5_ASAP7_75t_L g355 ( 
.A1(n_349),
.A2(n_345),
.A3(n_352),
.B1(n_342),
.B2(n_147),
.C1(n_159),
.C2(n_116),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_349),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_357),
.Y(n_361)
);


endmodule