module fake_netlist_6_1010_n_104 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_104);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_104;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_17),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_R g40 ( 
.A(n_24),
.B(n_14),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_R g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_26),
.C(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_19),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_20),
.B(n_23),
.C(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_20),
.Y(n_51)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_27),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_27),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_39),
.B(n_38),
.C(n_26),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_37),
.B1(n_42),
.B2(n_31),
.Y(n_56)
);

AO32x2_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_43),
.A3(n_40),
.B1(n_19),
.B2(n_30),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_31),
.C(n_30),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI21x1_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_50),
.B(n_52),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_47),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_52),
.B(n_39),
.Y(n_63)
);

AO32x2_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_45),
.A3(n_53),
.B1(n_3),
.B2(n_5),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AOI211xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_38),
.B(n_53),
.C(n_58),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

AOI31xp33_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_64),
.A3(n_53),
.B(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_63),
.Y(n_78)
);

OR2x6_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_64),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_71),
.Y(n_84)
);

NOR2xp67_ASAP7_75t_SL g85 ( 
.A(n_83),
.B(n_72),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_78),
.B(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_70),
.B1(n_45),
.B2(n_64),
.Y(n_87)
);

AOI211xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_81),
.B(n_79),
.C(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_81),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_84),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_79),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_91),
.B1(n_87),
.B2(n_45),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_82),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_95),
.Y(n_100)
);

AO211x2_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_94),
.B(n_2),
.C(n_6),
.Y(n_101)
);

OAI211xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_99),
.B(n_101),
.C(n_9),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_0),
.B1(n_7),
.B2(n_9),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_7),
.B(n_11),
.Y(n_104)
);


endmodule