module fake_jpeg_15805_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_16),
.C(n_35),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_0),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_19),
.A2(n_29),
.B1(n_36),
.B2(n_34),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_33),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_7),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_73),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_29),
.B1(n_19),
.B2(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_67),
.A2(n_72),
.B1(n_78),
.B2(n_90),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_68),
.A2(n_71),
.B1(n_92),
.B2(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_36),
.B1(n_31),
.B2(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_0),
.B1(n_6),
.B2(n_8),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_20),
.B1(n_31),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_14),
.B1(n_92),
.B2(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_84),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_86),
.B(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_0),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_23),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_33),
.C(n_3),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_44),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_18),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_32),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_10),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_108),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_0),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_6),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_11),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_11),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_95),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_76),
.B1(n_66),
.B2(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_14),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_130),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_14),
.B(n_84),
.C(n_80),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_87),
.C(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_85),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_85),
.B(n_96),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_154),
.B(n_111),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_74),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_112),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_66),
.B(n_77),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_115),
.B(n_116),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_95),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_82),
.B1(n_83),
.B2(n_123),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_110),
.B1(n_107),
.B2(n_102),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_82),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_115),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_128),
.B1(n_122),
.B2(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_172),
.B1(n_178),
.B2(n_173),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_120),
.B(n_104),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_122),
.B1(n_104),
.B2(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_143),
.B(n_118),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_154),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_141),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_144),
.B1(n_134),
.B2(n_132),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_143),
.B(n_147),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_146),
.B1(n_152),
.B2(n_155),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_184),
.B1(n_198),
.B2(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_193),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_136),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_140),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_177),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_203),
.A2(n_189),
.B1(n_181),
.B2(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_211),
.B1(n_201),
.B2(n_179),
.Y(n_214)
);

OAI321xp33_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_196),
.A3(n_186),
.B1(n_170),
.B2(n_159),
.C(n_177),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_200),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_184),
.B1(n_160),
.B2(n_183),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_204),
.B(n_202),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_207),
.B1(n_209),
.B2(n_206),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_182),
.A3(n_214),
.B1(n_188),
.B2(n_212),
.C1(n_201),
.C2(n_185),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_R g217 ( 
.A(n_216),
.B(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_172),
.Y(n_219)
);


endmodule