module real_aes_12168_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1584;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_0), .A2(n_143), .B1(n_366), .B2(n_823), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_0), .A2(n_143), .B1(n_503), .B2(n_809), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_1), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_1), .A2(n_11), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_2), .A2(n_79), .B1(n_634), .B2(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g970 ( .A(n_2), .Y(n_970) );
INVx1_ASAP7_75t_L g681 ( .A(n_3), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_4), .A2(n_302), .B1(n_1269), .B2(n_1277), .Y(n_1295) );
INVx1_ASAP7_75t_L g1182 ( .A(n_5), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_6), .A2(n_205), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_6), .A2(n_205), .B1(n_469), .B2(n_471), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_7), .A2(n_17), .B1(n_997), .B2(n_998), .Y(n_996) );
INVxp67_ASAP7_75t_SL g1027 ( .A(n_7), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_8), .A2(n_153), .B1(n_471), .B2(n_482), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1538 ( .A1(n_8), .A2(n_153), .B1(n_660), .B2(n_666), .Y(n_1538) );
INVx1_ASAP7_75t_L g358 ( .A(n_9), .Y(n_358) );
INVx1_ASAP7_75t_L g942 ( .A(n_10), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_10), .A2(n_228), .B1(n_455), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g380 ( .A(n_11), .Y(n_380) );
INVxp33_ASAP7_75t_SL g989 ( .A(n_12), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_12), .A2(n_278), .B1(n_695), .B2(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g891 ( .A(n_13), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_13), .A2(n_66), .B1(n_401), .B2(n_815), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g1242 ( .A1(n_14), .A2(n_262), .B1(n_482), .B2(n_1243), .Y(n_1242) );
INVxp67_ASAP7_75t_L g1252 ( .A(n_14), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g985 ( .A(n_15), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_15), .A2(n_193), .B1(n_414), .B2(n_800), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1565 ( .A(n_16), .Y(n_1565) );
INVxp67_ASAP7_75t_SL g1028 ( .A(n_17), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_18), .A2(n_68), .B1(n_1610), .B2(n_1614), .C(n_1617), .Y(n_1609) );
INVx1_ASAP7_75t_L g1625 ( .A(n_18), .Y(n_1625) );
INVx1_ASAP7_75t_L g346 ( .A(n_19), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_19), .A2(n_60), .B1(n_401), .B2(n_444), .Y(n_458) );
INVx1_ASAP7_75t_L g617 ( .A(n_20), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_20), .A2(n_282), .B1(n_645), .B2(n_647), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_21), .A2(n_256), .B1(n_1285), .B2(n_1291), .Y(n_1296) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_22), .A2(n_306), .B1(n_366), .B2(n_823), .Y(n_960) );
INVx1_ASAP7_75t_L g966 ( .A(n_22), .Y(n_966) );
XOR2x2_ASAP7_75t_L g976 ( .A(n_23), .B(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_24), .A2(n_73), .B1(n_533), .B2(n_536), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_24), .A2(n_73), .B1(n_567), .B2(n_570), .Y(n_566) );
CKINVDCx16_ASAP7_75t_R g1322 ( .A(n_25), .Y(n_1322) );
INVxp67_ASAP7_75t_SL g1195 ( .A(n_26), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_26), .A2(n_190), .B1(n_775), .B2(n_998), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_27), .A2(n_225), .B1(n_441), .B2(n_442), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_27), .A2(n_225), .B1(n_634), .B2(n_843), .Y(n_911) );
OAI211xp5_ASAP7_75t_L g1135 ( .A1(n_28), .A2(n_654), .B(n_1136), .C(n_1137), .Y(n_1135) );
INVx1_ASAP7_75t_L g1155 ( .A(n_28), .Y(n_1155) );
INVx1_ASAP7_75t_L g504 ( .A(n_29), .Y(n_504) );
INVx1_ASAP7_75t_L g1229 ( .A(n_30), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_30), .A2(n_33), .B1(n_411), .B2(n_968), .Y(n_1249) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_31), .A2(n_84), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_31), .A2(n_84), .B1(n_775), .B2(n_1122), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_32), .Y(n_1162) );
INVx1_ASAP7_75t_L g1230 ( .A(n_33), .Y(n_1230) );
INVx1_ASAP7_75t_L g880 ( .A(n_34), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_34), .A2(n_141), .B1(n_482), .B2(n_483), .Y(n_915) );
INVx1_ASAP7_75t_L g317 ( .A(n_35), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g1517 ( .A1(n_36), .A2(n_209), .B1(n_1052), .B2(n_1105), .C(n_1518), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_36), .A2(n_209), .B1(n_482), .B2(n_483), .Y(n_1528) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_37), .A2(n_58), .B1(n_326), .B2(n_430), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_37), .A2(n_297), .B1(n_645), .B2(n_647), .Y(n_868) );
XNOR2xp5_ASAP7_75t_L g673 ( .A(n_38), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_38), .A2(n_139), .B1(n_1269), .B2(n_1277), .Y(n_1268) );
INVxp67_ASAP7_75t_L g749 ( .A(n_39), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_39), .A2(n_243), .B1(n_775), .B2(n_776), .Y(n_774) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_40), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_40), .A2(n_170), .B1(n_455), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1232 ( .A(n_41), .Y(n_1232) );
INVxp67_ASAP7_75t_SL g740 ( .A(n_42), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_42), .A2(n_311), .B1(n_411), .B2(n_414), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_43), .A2(n_184), .B1(n_1281), .B2(n_1310), .Y(n_1309) );
INVxp33_ASAP7_75t_L g1101 ( .A(n_44), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_44), .A2(n_251), .B1(n_478), .B2(n_1120), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_45), .A2(n_294), .B1(n_645), .B2(n_656), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_45), .A2(n_216), .B1(n_550), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_46), .A2(n_269), .B1(n_441), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_46), .A2(n_269), .B1(n_642), .B2(n_843), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_47), .A2(n_112), .B1(n_1269), .B2(n_1277), .Y(n_1289) );
AO221x2_ASAP7_75t_L g1297 ( .A1(n_48), .A2(n_219), .B1(n_1285), .B2(n_1291), .C(n_1298), .Y(n_1297) );
CKINVDCx16_ASAP7_75t_R g1323 ( .A(n_49), .Y(n_1323) );
AOI22xp5_ASAP7_75t_SL g1327 ( .A1(n_50), .A2(n_204), .B1(n_1281), .B2(n_1285), .Y(n_1327) );
INVxp33_ASAP7_75t_SL g1183 ( .A(n_51), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_51), .A2(n_173), .B1(n_455), .B2(n_812), .Y(n_1200) );
INVxp33_ASAP7_75t_SL g1197 ( .A(n_52), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_52), .A2(n_70), .B1(n_523), .B2(n_1212), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_53), .A2(n_77), .B1(n_660), .B2(n_666), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_53), .A2(n_77), .B1(n_642), .B2(n_770), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_54), .A2(n_56), .B1(n_756), .B2(n_758), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_54), .A2(n_56), .B1(n_699), .B2(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_55), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_55), .A2(n_69), .B1(n_483), .B2(n_580), .Y(n_579) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_57), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_57), .A2(n_188), .B1(n_550), .B2(n_1052), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_58), .A2(n_160), .B1(n_564), .B2(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1530 ( .A(n_59), .Y(n_1530) );
INVx1_ASAP7_75t_L g369 ( .A(n_60), .Y(n_369) );
INVx1_ASAP7_75t_L g399 ( .A(n_61), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_61), .A2(n_220), .B1(n_478), .B2(n_479), .Y(n_477) );
OAI211xp5_ASAP7_75t_L g1510 ( .A1(n_62), .A2(n_654), .B(n_1511), .C(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g1524 ( .A(n_62), .Y(n_1524) );
CKINVDCx14_ASAP7_75t_R g1371 ( .A(n_63), .Y(n_1371) );
INVx1_ASAP7_75t_L g883 ( .A(n_64), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_64), .A2(n_155), .B1(n_466), .B2(n_914), .Y(n_913) );
OAI211xp5_ASAP7_75t_L g920 ( .A1(n_64), .A2(n_511), .B(n_921), .C(n_924), .Y(n_920) );
XNOR2xp5_ASAP7_75t_L g934 ( .A(n_65), .B(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g896 ( .A(n_66), .Y(n_896) );
OAI211xp5_ASAP7_75t_L g928 ( .A1(n_66), .A2(n_654), .B(n_929), .C(n_931), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g1580 ( .A1(n_67), .A2(n_276), .B1(n_1581), .B2(n_1583), .Y(n_1580) );
INVx1_ASAP7_75t_L g1618 ( .A(n_67), .Y(n_1618) );
INVx1_ASAP7_75t_L g1627 ( .A(n_68), .Y(n_1627) );
INVxp67_ASAP7_75t_SL g510 ( .A(n_69), .Y(n_510) );
INVxp67_ASAP7_75t_SL g1191 ( .A(n_70), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_71), .A2(n_126), .B1(n_695), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_71), .A2(n_126), .B1(n_769), .B2(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g893 ( .A(n_72), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_72), .A2(n_285), .B1(n_455), .B2(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g857 ( .A(n_74), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_75), .A2(n_179), .B1(n_1269), .B2(n_1308), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_76), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_78), .A2(n_230), .B1(n_753), .B2(n_1159), .C(n_1160), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_78), .A2(n_230), .B1(n_483), .B2(n_569), .Y(n_1168) );
INVx1_ASAP7_75t_L g971 ( .A(n_79), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_80), .A2(n_90), .B1(n_816), .B2(n_1208), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_80), .A2(n_90), .B1(n_523), .B2(n_1212), .Y(n_1211) );
CKINVDCx14_ASAP7_75t_R g1299 ( .A(n_81), .Y(n_1299) );
AOI22xp33_ASAP7_75t_SL g1542 ( .A1(n_81), .A2(n_1543), .B1(n_1546), .B2(n_1630), .Y(n_1542) );
AO22x2_ASAP7_75t_L g1548 ( .A1(n_81), .A2(n_1299), .B1(n_1549), .B2(n_1629), .Y(n_1548) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_82), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_83), .A2(n_215), .B1(n_660), .B2(n_666), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_83), .A2(n_215), .B1(n_471), .B2(n_569), .Y(n_1172) );
BUFx2_ASAP7_75t_L g396 ( .A(n_85), .Y(n_396) );
BUFx2_ASAP7_75t_L g437 ( .A(n_85), .Y(n_437) );
INVx1_ASAP7_75t_L g559 ( .A(n_85), .Y(n_559) );
OR2x2_ASAP7_75t_L g1584 ( .A(n_85), .B(n_1585), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_86), .A2(n_218), .B1(n_766), .B2(n_993), .Y(n_992) );
INVxp67_ASAP7_75t_SL g1022 ( .A(n_86), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_87), .A2(n_211), .B1(n_541), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_87), .A2(n_211), .B1(n_699), .B2(n_701), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_88), .A2(n_299), .B1(n_775), .B2(n_776), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_88), .A2(n_299), .B1(n_1009), .B2(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1185 ( .A(n_89), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_89), .A2(n_103), .B1(n_444), .B2(n_544), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_91), .A2(n_280), .B1(n_544), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_91), .A2(n_280), .B1(n_366), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_92), .A2(n_244), .B1(n_766), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_92), .A2(n_244), .B1(n_502), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_93), .A2(n_242), .B1(n_455), .B2(n_1204), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_93), .A2(n_242), .B1(n_847), .B2(n_1214), .Y(n_1213) );
XNOR2xp5_ASAP7_75t_L g781 ( .A(n_94), .B(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_95), .A2(n_270), .B1(n_541), .B2(n_544), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_95), .A2(n_270), .B1(n_562), .B2(n_564), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_96), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_97), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_98), .A2(n_303), .B1(n_564), .B2(n_841), .Y(n_1241) );
INVxp33_ASAP7_75t_L g1254 ( .A(n_98), .Y(n_1254) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_99), .A2(n_217), .B1(n_656), .B2(n_657), .Y(n_1515) );
AOI221xp5_ASAP7_75t_L g1521 ( .A1(n_99), .A2(n_217), .B1(n_533), .B2(n_551), .C(n_1522), .Y(n_1521) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_100), .A2(n_1505), .B1(n_1506), .B2(n_1507), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1505 ( .A(n_100), .Y(n_1505) );
INVx1_ASAP7_75t_L g869 ( .A(n_101), .Y(n_869) );
INVx1_ASAP7_75t_L g1519 ( .A(n_102), .Y(n_1519) );
INVxp33_ASAP7_75t_SL g1179 ( .A(n_103), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_104), .A2(n_134), .B1(n_448), .B2(n_809), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_104), .A2(n_134), .B1(n_478), .B2(n_479), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g1161 ( .A(n_105), .Y(n_1161) );
AO22x2_ASAP7_75t_L g1219 ( .A1(n_106), .A2(n_1220), .B1(n_1255), .B2(n_1256), .Y(n_1219) );
INVx1_ASAP7_75t_L g1255 ( .A(n_106), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_107), .A2(n_202), .B1(n_714), .B2(n_716), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_107), .A2(n_202), .B1(n_660), .B2(n_666), .Y(n_726) );
INVx1_ASAP7_75t_L g1514 ( .A(n_108), .Y(n_1514) );
INVxp33_ASAP7_75t_SL g1098 ( .A(n_109), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_109), .A2(n_191), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_110), .A2(n_223), .B1(n_562), .B2(n_766), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g1068 ( .A(n_110), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_111), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_111), .A2(n_260), .B1(n_478), .B2(n_766), .Y(n_773) );
XOR2xp5_ASAP7_75t_L g590 ( .A(n_112), .B(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_113), .A2(n_266), .B1(n_483), .B2(n_569), .Y(n_1236) );
AOI22xp33_ASAP7_75t_SL g1244 ( .A1(n_113), .A2(n_266), .B1(n_441), .B2(n_442), .Y(n_1244) );
INVx1_ASAP7_75t_L g941 ( .A(n_114), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_114), .A2(n_231), .B1(n_544), .B2(n_815), .Y(n_954) );
INVx1_ASAP7_75t_L g1042 ( .A(n_115), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_115), .A2(n_263), .B1(n_411), .B2(n_968), .Y(n_1069) );
INVxp33_ASAP7_75t_L g516 ( .A(n_116), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_116), .A2(n_163), .B1(n_541), .B2(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_117), .A2(n_216), .B1(n_647), .B2(n_657), .Y(n_677) );
INVxp33_ASAP7_75t_SL g725 ( .A(n_117), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g1107 ( .A1(n_118), .A2(n_258), .B1(n_1108), .B2(n_1110), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_118), .A2(n_258), .B1(n_993), .B2(n_1120), .Y(n_1119) );
INVxp33_ASAP7_75t_SL g1085 ( .A(n_119), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_119), .A2(n_295), .B1(n_1113), .B2(n_1115), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_120), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_120), .A2(n_187), .B1(n_503), .B2(n_833), .Y(n_1239) );
XNOR2xp5_ASAP7_75t_L g727 ( .A(n_121), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g494 ( .A(n_122), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g1563 ( .A(n_123), .Y(n_1563) );
INVx1_ASAP7_75t_L g614 ( .A(n_124), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_124), .A2(n_252), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI22xp5_ASAP7_75t_SL g1326 ( .A1(n_125), .A2(n_146), .B1(n_1269), .B2(n_1277), .Y(n_1326) );
INVxp33_ASAP7_75t_SL g1224 ( .A(n_127), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1238 ( .A1(n_127), .A2(n_275), .B1(n_441), .B2(n_442), .Y(n_1238) );
INVx1_ASAP7_75t_L g1273 ( .A(n_128), .Y(n_1273) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_129), .A2(n_511), .B(n_662), .C(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_129), .A2(n_227), .B1(n_819), .B2(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1558 ( .A(n_130), .Y(n_1558) );
AOI22xp33_ASAP7_75t_SL g1606 ( .A1(n_130), .A2(n_272), .B1(n_471), .B2(n_849), .Y(n_1606) );
INVxp33_ASAP7_75t_SL g1034 ( .A(n_131), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_131), .A2(n_167), .B1(n_541), .B2(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_132), .A2(n_214), .B1(n_444), .B2(n_448), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_132), .A2(n_214), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_133), .A2(n_203), .B1(n_805), .B2(n_806), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_133), .A2(n_203), .B1(n_642), .B2(n_770), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_135), .Y(n_497) );
INVx1_ASAP7_75t_L g1091 ( .A(n_136), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_136), .A2(n_247), .B1(n_506), .B2(n_968), .Y(n_1096) );
AO22x2_ASAP7_75t_SL g1029 ( .A1(n_137), .A2(n_1030), .B1(n_1031), .B2(n_1075), .Y(n_1029) );
CKINVDCx16_ASAP7_75t_R g1030 ( .A(n_137), .Y(n_1030) );
INVx1_ASAP7_75t_L g637 ( .A(n_138), .Y(n_637) );
OAI22xp33_ASAP7_75t_SL g665 ( .A1(n_138), .A2(n_152), .B1(n_326), .B2(n_666), .Y(n_665) );
INVxp33_ASAP7_75t_SL g980 ( .A(n_140), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_140), .A2(n_150), .B1(n_502), .B2(n_542), .Y(n_1010) );
INVx1_ASAP7_75t_L g881 ( .A(n_141), .Y(n_881) );
INVx1_ASAP7_75t_L g1274 ( .A(n_142), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_142), .B(n_1272), .Y(n_1279) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_144), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_145), .A2(n_197), .B1(n_503), .B2(n_809), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_145), .A2(n_197), .B1(n_366), .B2(n_823), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_147), .A2(n_157), .B1(n_645), .B2(n_656), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_147), .A2(n_264), .B1(n_533), .B2(n_1049), .C(n_1151), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_148), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_148), .A2(n_194), .B1(n_753), .B2(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g329 ( .A(n_149), .Y(n_329) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_150), .Y(n_983) );
INVxp33_ASAP7_75t_L g1084 ( .A(n_151), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_151), .A2(n_288), .B1(n_503), .B2(n_756), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_152), .A2(n_246), .B1(n_471), .B2(n_642), .Y(n_641) );
BUFx3_ASAP7_75t_L g355 ( .A(n_154), .Y(n_355) );
INVx1_ASAP7_75t_L g388 ( .A(n_154), .Y(n_388) );
INVx1_ASAP7_75t_L g887 ( .A(n_155), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_156), .A2(n_158), .B1(n_701), .B2(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g724 ( .A(n_156), .Y(n_724) );
INVx1_ASAP7_75t_L g1152 ( .A(n_157), .Y(n_1152) );
INVx1_ASAP7_75t_L g721 ( .A(n_158), .Y(n_721) );
INVxp33_ASAP7_75t_L g508 ( .A(n_159), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_159), .A2(n_212), .B1(n_562), .B2(n_583), .Y(n_582) );
OAI211xp5_ASAP7_75t_SL g852 ( .A1(n_160), .A2(n_511), .B(n_853), .C(n_856), .Y(n_852) );
INVx1_ASAP7_75t_L g1552 ( .A(n_161), .Y(n_1552) );
AOI21xp33_ASAP7_75t_L g1607 ( .A1(n_161), .A2(n_569), .B(n_1608), .Y(n_1607) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_162), .A2(n_207), .B1(n_533), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_162), .A2(n_207), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_L g521 ( .A(n_163), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_164), .A2(n_281), .B1(n_550), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_164), .A2(n_281), .B1(n_703), .B2(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_165), .A2(n_304), .B1(n_541), .B2(n_1047), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_165), .A2(n_304), .B1(n_523), .B2(n_699), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_166), .A2(n_297), .B1(n_544), .B2(n_809), .Y(n_837) );
INVx1_ASAP7_75t_L g863 ( .A(n_166), .Y(n_863) );
INVx1_ASAP7_75t_L g1040 ( .A(n_167), .Y(n_1040) );
INVx1_ASAP7_75t_L g737 ( .A(n_168), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_168), .A2(n_172), .B1(n_688), .B2(n_756), .Y(n_763) );
INVx1_ASAP7_75t_L g790 ( .A(n_169), .Y(n_790) );
INVx1_ASAP7_75t_L g793 ( .A(n_170), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g1130 ( .A(n_171), .B(n_1131), .Y(n_1130) );
INVxp33_ASAP7_75t_SL g731 ( .A(n_172), .Y(n_731) );
INVxp33_ASAP7_75t_SL g1180 ( .A(n_173), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_174), .A2(n_248), .B1(n_645), .B2(n_647), .Y(n_1509) );
INVx1_ASAP7_75t_L g1537 ( .A(n_174), .Y(n_1537) );
INVx1_ASAP7_75t_L g394 ( .A(n_175), .Y(n_394) );
INVx1_ASAP7_75t_L g1591 ( .A(n_175), .Y(n_1591) );
INVx1_ASAP7_75t_L g858 ( .A(n_176), .Y(n_858) );
INVxp67_ASAP7_75t_L g435 ( .A(n_177), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_177), .A2(n_253), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g946 ( .A(n_178), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_178), .A2(n_283), .B1(n_506), .B2(n_968), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g1369 ( .A(n_180), .Y(n_1369) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_181), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_181), .A2(n_287), .B1(n_471), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_182), .A2(n_301), .B1(n_441), .B2(n_442), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_182), .A2(n_301), .B1(n_847), .B2(n_958), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g1562 ( .A(n_183), .Y(n_1562) );
CKINVDCx14_ASAP7_75t_R g1301 ( .A(n_185), .Y(n_1301) );
INVx1_ASAP7_75t_L g1513 ( .A(n_186), .Y(n_1513) );
INVxp33_ASAP7_75t_SL g1223 ( .A(n_187), .Y(n_1223) );
INVxp33_ASAP7_75t_SL g1035 ( .A(n_188), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_189), .A2(n_261), .B1(n_634), .B2(n_847), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_189), .A2(n_261), .B1(n_660), .B2(n_666), .Y(n_851) );
INVxp33_ASAP7_75t_L g1194 ( .A(n_190), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g1099 ( .A(n_191), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_192), .A2(n_264), .B1(n_647), .B2(n_657), .Y(n_1134) );
INVx1_ASAP7_75t_L g1147 ( .A(n_192), .Y(n_1147) );
INVxp67_ASAP7_75t_SL g986 ( .A(n_193), .Y(n_986) );
INVxp33_ASAP7_75t_SL g732 ( .A(n_194), .Y(n_732) );
INVx1_ASAP7_75t_L g1037 ( .A(n_195), .Y(n_1037) );
INVx1_ASAP7_75t_L g602 ( .A(n_196), .Y(n_602) );
INVx1_ASAP7_75t_L g988 ( .A(n_198), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1575 ( .A1(n_199), .A2(n_206), .B1(n_1576), .B2(n_1578), .Y(n_1575) );
INVx1_ASAP7_75t_L g1599 ( .A(n_199), .Y(n_1599) );
OA332x1_ASAP7_75t_L g1550 ( .A1(n_200), .A2(n_594), .A3(n_1551), .B1(n_1557), .B2(n_1561), .B3(n_1564), .C1(n_1569), .C2(n_1570), .Y(n_1550) );
AOI21xp5_ASAP7_75t_L g1603 ( .A1(n_200), .A2(n_823), .B(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g789 ( .A(n_201), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g1602 ( .A1(n_206), .A2(n_276), .B1(n_471), .B2(n_569), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_208), .A2(n_235), .B1(n_544), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_208), .A2(n_235), .B1(n_478), .B2(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g1520 ( .A(n_210), .Y(n_1520) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_212), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_213), .A2(n_239), .B1(n_441), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g867 ( .A(n_213), .Y(n_867) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_218), .Y(n_1025) );
INVxp33_ASAP7_75t_L g419 ( .A(n_220), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_221), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g1317 ( .A(n_222), .Y(n_1317) );
INVxp33_ASAP7_75t_L g1074 ( .A(n_223), .Y(n_1074) );
BUFx3_ASAP7_75t_L g357 ( .A(n_224), .Y(n_357) );
INVx1_ASAP7_75t_L g383 ( .A(n_224), .Y(n_383) );
INVx1_ASAP7_75t_L g1531 ( .A(n_226), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_227), .A2(n_284), .B1(n_326), .B2(n_430), .Y(n_801) );
INVx1_ASAP7_75t_L g939 ( .A(n_228), .Y(n_939) );
AO221x2_ASAP7_75t_L g1366 ( .A1(n_229), .A2(n_286), .B1(n_1310), .B2(n_1367), .C(n_1368), .Y(n_1366) );
INVx1_ASAP7_75t_L g944 ( .A(n_231), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1290 ( .A1(n_232), .A2(n_233), .B1(n_1285), .B2(n_1291), .Y(n_1290) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_234), .Y(n_325) );
INVx1_ASAP7_75t_L g462 ( .A(n_234), .Y(n_462) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_234), .B(n_409), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_234), .B(n_292), .Y(n_1585) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_236), .Y(n_653) );
INVx1_ASAP7_75t_L g342 ( .A(n_237), .Y(n_342) );
INVx2_ASAP7_75t_L g350 ( .A(n_238), .Y(n_350) );
OR2x2_ASAP7_75t_L g1590 ( .A(n_238), .B(n_1591), .Y(n_1590) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_239), .Y(n_866) );
INVx1_ASAP7_75t_L g1087 ( .A(n_240), .Y(n_1087) );
INVx1_ASAP7_75t_L g1187 ( .A(n_241), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_241), .A2(n_273), .B1(n_411), .B2(n_414), .Y(n_1192) );
INVxp67_ASAP7_75t_L g748 ( .A(n_243), .Y(n_748) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_245), .A2(n_638), .B(n_654), .C(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_245), .A2(n_294), .B1(n_542), .B2(n_688), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_246), .A2(n_282), .B1(n_430), .B2(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1092 ( .A(n_247), .Y(n_1092) );
INVx1_ASAP7_75t_L g1523 ( .A(n_248), .Y(n_1523) );
AOI22xp5_ASAP7_75t_SL g1280 ( .A1(n_249), .A2(n_254), .B1(n_1281), .B2(n_1285), .Y(n_1280) );
INVx1_ASAP7_75t_L g734 ( .A(n_250), .Y(n_734) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_251), .Y(n_1095) );
INVx1_ASAP7_75t_L g612 ( .A(n_252), .Y(n_612) );
INVx1_ASAP7_75t_L g427 ( .A(n_253), .Y(n_427) );
AO22x2_ASAP7_75t_L g876 ( .A1(n_255), .A2(n_877), .B1(n_916), .B2(n_917), .Y(n_876) );
INVxp67_ASAP7_75t_L g916 ( .A(n_255), .Y(n_916) );
INVx1_ASAP7_75t_L g640 ( .A(n_257), .Y(n_640) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_257), .A2(n_511), .B(n_662), .C(n_664), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_259), .A2(n_290), .B1(n_371), .B2(n_376), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_259), .A2(n_290), .B1(n_411), .B2(n_414), .Y(n_410) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_260), .Y(n_745) );
INVxp33_ASAP7_75t_L g1251 ( .A(n_262), .Y(n_1251) );
INVx1_ASAP7_75t_L g1043 ( .A(n_263), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_265), .Y(n_888) );
INVx1_ASAP7_75t_L g489 ( .A(n_267), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g1568 ( .A(n_268), .Y(n_1568) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_271), .A2(n_284), .B1(n_645), .B2(n_647), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_271), .A2(n_296), .B1(n_815), .B2(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g1554 ( .A(n_272), .Y(n_1554) );
INVx1_ASAP7_75t_L g1186 ( .A(n_273), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_274), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_274), .A2(n_293), .B1(n_550), .B2(n_551), .Y(n_549) );
INVxp33_ASAP7_75t_SL g1233 ( .A(n_275), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_277), .B(n_317), .Y(n_1276) );
AND3x2_ASAP7_75t_L g1284 ( .A(n_277), .B(n_317), .C(n_1273), .Y(n_1284) );
INVxp33_ASAP7_75t_SL g981 ( .A(n_278), .Y(n_981) );
INVx2_ASAP7_75t_L g330 ( .A(n_279), .Y(n_330) );
INVx1_ASAP7_75t_L g945 ( .A(n_283), .Y(n_945) );
INVx1_ASAP7_75t_L g898 ( .A(n_285), .Y(n_898) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_287), .Y(n_604) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_288), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_289), .Y(n_1138) );
INVx1_ASAP7_75t_L g598 ( .A(n_291), .Y(n_598) );
INVx1_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
INVx2_ASAP7_75t_L g409 ( .A(n_292), .Y(n_409) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_293), .Y(n_519) );
INVxp33_ASAP7_75t_L g1088 ( .A(n_295), .Y(n_1088) );
INVx1_ASAP7_75t_L g786 ( .A(n_296), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g1139 ( .A(n_298), .Y(n_1139) );
INVx1_ASAP7_75t_L g680 ( .A(n_300), .Y(n_680) );
XOR2x2_ASAP7_75t_L g1175 ( .A(n_302), .B(n_1176), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_303), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1559 ( .A(n_305), .Y(n_1559) );
INVx1_ASAP7_75t_L g973 ( .A(n_306), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_307), .A2(n_309), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
INVxp33_ASAP7_75t_L g1071 ( .A(n_307), .Y(n_1071) );
INVx1_ASAP7_75t_L g620 ( .A(n_308), .Y(n_620) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_309), .Y(n_1072) );
AO22x1_ASAP7_75t_L g1079 ( .A1(n_310), .A2(n_1080), .B1(n_1081), .B2(n_1129), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_310), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_311), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_333), .B(n_1261), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
AND2x4_ASAP7_75t_L g1545 ( .A(n_315), .B(n_321), .Y(n_1545) );
NOR2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_SL g1541 ( .A(n_316), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_316), .B(n_318), .Y(n_1632) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_318), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g436 ( .A(n_323), .B(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_L g513 ( .A(n_323), .B(n_437), .Y(n_513) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g452 ( .A(n_324), .B(n_332), .Y(n_452) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g595 ( .A(n_325), .B(n_422), .Y(n_595) );
INVx8_ASAP7_75t_L g418 ( .A(n_326), .Y(n_418) );
OR2x6_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
OR2x6_ASAP7_75t_L g430 ( .A(n_327), .B(n_421), .Y(n_430) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_327), .Y(n_597) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_327), .Y(n_616) );
INVx2_ASAP7_75t_SL g1154 ( .A(n_327), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_327), .B(n_1584), .Y(n_1583) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g403 ( .A(n_329), .Y(n_403) );
INVx1_ASAP7_75t_L g416 ( .A(n_329), .Y(n_416) );
INVx2_ASAP7_75t_L g424 ( .A(n_329), .Y(n_424) );
AND2x4_ASAP7_75t_L g434 ( .A(n_329), .B(n_404), .Y(n_434) );
AND2x2_ASAP7_75t_L g447 ( .A(n_329), .B(n_330), .Y(n_447) );
INVx2_ASAP7_75t_L g404 ( .A(n_330), .Y(n_404) );
INVx1_ASAP7_75t_L g413 ( .A(n_330), .Y(n_413) );
INVx1_ASAP7_75t_L g426 ( .A(n_330), .Y(n_426) );
INVx1_ASAP7_75t_L g601 ( .A(n_330), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_330), .B(n_424), .Y(n_607) );
AND2x4_ASAP7_75t_L g412 ( .A(n_331), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g414 ( .A(n_332), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g968 ( .A(n_332), .B(n_415), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_871), .B2(n_872), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_670), .B1(n_671), .B2(n_870), .Y(n_335) );
INVx1_ASAP7_75t_L g870 ( .A(n_336), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_586), .B2(n_669), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_487), .B2(n_585), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
XNOR2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_392), .B(n_397), .C(n_438), .Y(n_343) );
NAND4xp25_ASAP7_75t_L g344 ( .A(n_345), .B(n_362), .C(n_379), .D(n_389), .Y(n_344) );
AOI22xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B1(n_358), .B2(n_359), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_347), .A2(n_381), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_347), .A2(n_381), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_347), .A2(n_381), .B1(n_941), .B2(n_942), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_347), .A2(n_381), .B1(n_390), .B2(n_980), .C(n_981), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_347), .A2(n_381), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_347), .A2(n_381), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_347), .A2(n_381), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
AND2x6_ASAP7_75t_L g385 ( .A(n_348), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g892 ( .A(n_348), .B(n_351), .Y(n_892) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_350), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
AND2x2_ASAP7_75t_L g475 ( .A(n_350), .B(n_394), .Y(n_475) );
INVx2_ASAP7_75t_L g486 ( .A(n_350), .Y(n_486) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g465 ( .A(n_352), .Y(n_465) );
INVx2_ASAP7_75t_L g563 ( .A(n_352), .Y(n_563) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_352), .Y(n_700) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_352), .Y(n_712) );
INVx1_ASAP7_75t_L g849 ( .A(n_352), .Y(n_849) );
INVx2_ASAP7_75t_SL g995 ( .A(n_352), .Y(n_995) );
INVx6_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g359 ( .A(n_353), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g478 ( .A(n_353), .Y(n_478) );
INVx2_ASAP7_75t_L g824 ( .A(n_353), .Y(n_824) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_353), .B(n_1595), .Y(n_1619) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g368 ( .A(n_355), .B(n_357), .Y(n_368) );
AND2x4_ASAP7_75t_L g382 ( .A(n_355), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g387 ( .A(n_357), .B(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_358), .A2(n_429), .B1(n_431), .B2(n_435), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_359), .A2(n_385), .B1(n_494), .B2(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g647 ( .A(n_359), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_359), .A2(n_385), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_359), .A2(n_385), .B1(n_888), .B2(n_898), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_359), .A2(n_385), .B1(n_938), .B2(n_939), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_359), .A2(n_385), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_359), .A2(n_385), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_359), .A2(n_385), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_359), .A2(n_385), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_359), .A2(n_385), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
AND2x4_ASAP7_75t_L g525 ( .A(n_360), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_360), .B(n_526), .Y(n_739) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_369), .B(n_370), .Y(n_362) );
INVx1_ASAP7_75t_L g1511 ( .A(n_363), .Y(n_1511) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
AND2x6_ASAP7_75t_L g381 ( .A(n_364), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
INVx1_ASAP7_75t_L g646 ( .A(n_364), .Y(n_646) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x6_ASAP7_75t_L g377 ( .A(n_365), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_366), .Y(n_895) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_366), .Y(n_1041) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g390 ( .A(n_367), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g467 ( .A(n_367), .Y(n_467) );
INVx2_ASAP7_75t_L g565 ( .A(n_367), .Y(n_565) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_367), .Y(n_767) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_368), .Y(n_480) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_372), .A2(n_377), .B1(n_620), .B2(n_650), .C1(n_652), .C2(n_653), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_372), .A2(n_377), .B1(n_857), .B2(n_858), .C1(n_863), .C2(n_864), .Y(n_862) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g526 ( .A(n_374), .Y(n_526) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g1613 ( .A(n_375), .Y(n_1613) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_377), .A2(n_497), .B1(n_504), .B2(n_521), .C1(n_522), .C2(n_524), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_377), .A2(n_525), .B1(n_680), .B2(n_681), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g736 ( .A1(n_377), .A2(n_583), .B1(n_737), .B2(n_738), .C1(n_739), .C2(n_740), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g785 ( .A1(n_377), .A2(n_739), .B1(n_786), .B2(n_787), .C1(n_789), .C2(n_790), .Y(n_785) );
AOI222xp33_ASAP7_75t_L g894 ( .A1(n_377), .A2(n_524), .B1(n_884), .B2(n_885), .C1(n_895), .C2(n_896), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_377), .A2(n_525), .B1(n_884), .B2(n_885), .Y(n_931) );
AOI222xp33_ASAP7_75t_L g943 ( .A1(n_377), .A2(n_701), .B1(n_739), .B2(n_944), .C1(n_945), .C2(n_946), .Y(n_943) );
AOI222xp33_ASAP7_75t_L g982 ( .A1(n_377), .A2(n_739), .B1(n_983), .B2(n_984), .C1(n_985), .C2(n_986), .Y(n_982) );
AOI222xp33_ASAP7_75t_L g1039 ( .A1(n_377), .A2(n_524), .B1(n_1040), .B2(n_1041), .C1(n_1042), .C2(n_1043), .Y(n_1039) );
AOI222xp33_ASAP7_75t_L g1089 ( .A1(n_377), .A2(n_479), .B1(n_739), .B2(n_1090), .C1(n_1091), .C2(n_1092), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_377), .A2(n_525), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
AOI222xp33_ASAP7_75t_L g1184 ( .A1(n_377), .A2(n_739), .B1(n_766), .B2(n_1185), .C1(n_1186), .C2(n_1187), .Y(n_1184) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_377), .A2(n_739), .B1(n_1226), .B2(n_1227), .C1(n_1229), .C2(n_1230), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_377), .A2(n_525), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
BUFx3_ASAP7_75t_L g1616 ( .A(n_378), .Y(n_1616) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_384), .B2(n_385), .Y(n_379) );
CKINVDCx6p67_ASAP7_75t_R g656 ( .A(n_381), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_381), .A2(n_385), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_381), .A2(n_385), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp5_ASAP7_75t_SL g890 ( .A1(n_381), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_381), .A2(n_892), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
INVx2_ASAP7_75t_SL g470 ( .A(n_382), .Y(n_470) );
BUFx3_ASAP7_75t_L g482 ( .A(n_382), .Y(n_482) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_382), .Y(n_569) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_382), .Y(n_634) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_382), .Y(n_642) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_382), .Y(n_769) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_382), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_382), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_382), .Y(n_1214) );
INVx1_ASAP7_75t_L g628 ( .A(n_383), .Y(n_628) );
INVx4_ASAP7_75t_L g657 ( .A(n_385), .Y(n_657) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_386), .Y(n_483) );
INVx1_ASAP7_75t_L g777 ( .A(n_386), .Y(n_777) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_386), .Y(n_847) );
INVx1_ASAP7_75t_L g963 ( .A(n_386), .Y(n_963) );
INVx1_ASAP7_75t_L g1123 ( .A(n_386), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_387), .Y(n_471) );
INVx1_ASAP7_75t_L g571 ( .A(n_387), .Y(n_571) );
INVx1_ASAP7_75t_L g844 ( .A(n_387), .Y(n_844) );
INVx2_ASAP7_75t_L g1001 ( .A(n_387), .Y(n_1001) );
INVx1_ASAP7_75t_L g627 ( .A(n_388), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_389), .B(n_515), .C(n_518), .D(n_520), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g889 ( .A(n_389), .B(n_890), .C(n_894), .D(n_897), .Y(n_889) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_389), .B(n_937), .C(n_940), .D(n_943), .Y(n_936) );
NAND4xp25_ASAP7_75t_SL g1032 ( .A(n_389), .B(n_1033), .C(n_1036), .D(n_1039), .Y(n_1032) );
NAND4xp25_ASAP7_75t_SL g1082 ( .A(n_389), .B(n_1083), .C(n_1086), .D(n_1089), .Y(n_1082) );
INVx5_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
CKINVDCx8_ASAP7_75t_R g654 ( .A(n_390), .Y(n_654) );
OAI31xp33_ASAP7_75t_SL g643 ( .A1(n_392), .A2(n_644), .A3(n_648), .B(n_655), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g675 ( .A1(n_392), .A2(n_676), .A3(n_677), .B(n_678), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_392), .A2(n_784), .B(n_794), .Y(n_783) );
OAI21xp5_ASAP7_75t_SL g860 ( .A1(n_392), .A2(n_861), .B(n_868), .Y(n_860) );
AOI211xp5_ASAP7_75t_L g935 ( .A1(n_392), .A2(n_936), .B(n_947), .C(n_964), .Y(n_935) );
OAI31xp33_ASAP7_75t_SL g1132 ( .A1(n_392), .A2(n_1133), .A3(n_1134), .B(n_1135), .Y(n_1132) );
AOI211x1_ASAP7_75t_L g1220 ( .A1(n_392), .A2(n_1221), .B(n_1234), .C(n_1246), .Y(n_1220) );
OAI31xp33_ASAP7_75t_L g1508 ( .A1(n_392), .A2(n_1509), .A3(n_1510), .B(n_1515), .Y(n_1508) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x4_ASAP7_75t_L g529 ( .A(n_393), .B(n_395), .Y(n_529) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g485 ( .A(n_394), .B(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g1620 ( .A(n_395), .Y(n_1620) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
OR2x6_ASAP7_75t_L g594 ( .A(n_396), .B(n_595), .Y(n_594) );
AOI31xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_417), .A3(n_428), .B(n_436), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_405), .C(n_410), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g1535 ( .A1(n_400), .A2(n_412), .B1(n_498), .B2(n_1513), .C1(n_1514), .C2(n_1531), .Y(n_1535) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g405 ( .A(n_402), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g449 ( .A(n_402), .Y(n_449) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_402), .Y(n_503) );
BUFx3_ASAP7_75t_L g545 ( .A(n_402), .Y(n_545) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_402), .Y(n_690) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_402), .Y(n_1056) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
CKINVDCx11_ASAP7_75t_R g511 ( .A(n_405), .Y(n_511) );
AOI211xp5_ASAP7_75t_L g744 ( .A1(n_405), .A2(n_448), .B(n_745), .C(n_746), .Y(n_744) );
AOI211xp5_ASAP7_75t_L g965 ( .A1(n_405), .A2(n_502), .B(n_966), .C(n_967), .Y(n_965) );
AOI211xp5_ASAP7_75t_L g1021 ( .A1(n_405), .A2(n_544), .B(n_1022), .C(n_1023), .Y(n_1021) );
AOI211xp5_ASAP7_75t_L g1067 ( .A1(n_405), .A2(n_544), .B(n_1068), .C(n_1069), .Y(n_1067) );
AOI211xp5_ASAP7_75t_L g1094 ( .A1(n_405), .A2(n_502), .B(n_1095), .C(n_1096), .Y(n_1094) );
AOI211xp5_ASAP7_75t_L g1189 ( .A1(n_405), .A2(n_1190), .B(n_1191), .C(n_1192), .Y(n_1189) );
AOI211xp5_ASAP7_75t_L g1247 ( .A1(n_405), .A2(n_502), .B(n_1248), .C(n_1249), .Y(n_1247) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g500 ( .A(n_407), .Y(n_500) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_408), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g422 ( .A(n_409), .Y(n_422) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g506 ( .A(n_412), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_412), .A2(n_498), .B1(n_652), .B2(n_653), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_412), .A2(n_680), .B1(n_681), .B2(n_690), .C1(n_721), .C2(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g800 ( .A(n_412), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_412), .A2(n_498), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI222xp33_ASAP7_75t_SL g1142 ( .A1(n_412), .A2(n_722), .B1(n_1138), .B2(n_1139), .C1(n_1143), .C2(n_1144), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1623 ( .A(n_413), .Y(n_1623) );
INVx1_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_416), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g619 ( .A(n_416), .B(n_601), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_427), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_418), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_418), .A2(n_493), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_418), .A2(n_429), .B1(n_734), .B2(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_418), .A2(n_493), .B1(n_887), .B2(n_888), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_418), .A2(n_493), .B1(n_938), .B2(n_973), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_418), .A2(n_493), .B1(n_988), .B2(n_1025), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_418), .A2(n_429), .B1(n_1037), .B2(n_1074), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g1100 ( .A1(n_418), .A2(n_429), .B1(n_1087), .B2(n_1101), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_418), .A2(n_493), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_418), .A2(n_429), .B1(n_1182), .B2(n_1197), .Y(n_1196) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_418), .A2(n_429), .B1(n_1232), .B2(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_418), .A2(n_493), .B1(n_1530), .B2(n_1537), .Y(n_1536) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_420), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
AOI22xp5_ASAP7_75t_SL g747 ( .A1(n_420), .A2(n_431), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_420), .A2(n_431), .B1(n_880), .B2(n_881), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_420), .A2(n_509), .B1(n_970), .B2(n_971), .Y(n_969) );
AOI22xp5_ASAP7_75t_SL g1026 ( .A1(n_420), .A2(n_509), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_420), .A2(n_431), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_420), .A2(n_509), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_420), .A2(n_509), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
AOI22xp33_ASAP7_75t_SL g1250 ( .A1(n_420), .A2(n_509), .B1(n_1251), .B2(n_1252), .Y(n_1250) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x4_ASAP7_75t_L g431 ( .A(n_421), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g509 ( .A(n_421), .B(n_432), .Y(n_509) );
INVx1_ASAP7_75t_L g667 ( .A(n_421), .Y(n_667) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_423), .Y(n_441) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_423), .Y(n_535) );
BUFx2_ASAP7_75t_L g550 ( .A(n_423), .Y(n_550) );
INVx1_ASAP7_75t_L g754 ( .A(n_423), .Y(n_754) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_423), .Y(n_1105) );
INVx1_ASAP7_75t_L g1114 ( .A(n_423), .Y(n_1114) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx5_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g493 ( .A(n_430), .Y(n_493) );
INVx5_ASAP7_75t_SL g660 ( .A(n_431), .Y(n_660) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_433), .Y(n_457) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_434), .Y(n_442) );
INVx3_ASAP7_75t_L g539 ( .A(n_434), .Y(n_539) );
INVx1_ASAP7_75t_L g1016 ( .A(n_434), .Y(n_1016) );
AOI31xp33_ASAP7_75t_L g1246 ( .A1(n_436), .A2(n_1247), .A3(n_1250), .B(n_1253), .Y(n_1246) );
AND2x4_ASAP7_75t_L g484 ( .A(n_437), .B(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g578 ( .A(n_437), .B(n_485), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_453), .C(n_463), .D(n_476), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .C(n_450), .Y(n_439) );
INVx2_ASAP7_75t_SL g552 ( .A(n_442), .Y(n_552) );
INVx4_ASAP7_75t_L g686 ( .A(n_442), .Y(n_686) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_442), .Y(n_1050) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_442), .Y(n_1052) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_SL g809 ( .A(n_445), .Y(n_809) );
INVx2_ASAP7_75t_L g833 ( .A(n_445), .Y(n_833) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g815 ( .A(n_446), .Y(n_815) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g543 ( .A(n_447), .Y(n_543) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g547 ( .A(n_450), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_450), .B(n_752), .C(n_755), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_450), .B(n_804), .C(n_808), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_450), .B(n_830), .C(n_832), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_450), .B(n_903), .C(n_904), .Y(n_902) );
NAND3xp33_ASAP7_75t_L g948 ( .A(n_450), .B(n_949), .C(n_950), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_450), .B(n_1104), .C(n_1107), .Y(n_1103) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_450), .Y(n_1163) );
NAND3xp33_ASAP7_75t_L g1202 ( .A(n_450), .B(n_1203), .C(n_1207), .Y(n_1202) );
AOI33xp33_ASAP7_75t_L g1240 ( .A1(n_450), .A2(n_484), .A3(n_1241), .B1(n_1242), .B2(n_1244), .B3(n_1245), .Y(n_1240) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AND2x2_ASAP7_75t_L g459 ( .A(n_451), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g473 ( .A(n_451), .B(n_474), .Y(n_473) );
OR2x6_ASAP7_75t_L g573 ( .A(n_451), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g692 ( .A(n_451), .B(n_452), .Y(n_692) );
OR2x2_ASAP7_75t_L g708 ( .A(n_451), .B(n_574), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_458), .C(n_459), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g621 ( .A(n_459), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_459), .B(n_906), .C(n_908), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_459), .B(n_952), .C(n_954), .Y(n_951) );
AOI33xp33_ASAP7_75t_L g1235 ( .A1(n_459), .A2(n_472), .A3(n_1236), .B1(n_1237), .B2(n_1238), .B3(n_1239), .Y(n_1235) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x6_ASAP7_75t_L g557 ( .A(n_461), .B(n_558), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .C(n_472), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g958 ( .A(n_470), .Y(n_958) );
INVx1_ASAP7_75t_L g706 ( .A(n_471), .Y(n_706) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_471), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_472), .B(n_818), .C(n_820), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_472), .B(n_840), .C(n_842), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_472), .B(n_910), .C(n_911), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_472), .B(n_956), .C(n_957), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g1118 ( .A(n_472), .B(n_1119), .C(n_1121), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1210 ( .A(n_472), .B(n_1211), .C(n_1213), .Y(n_1210) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g622 ( .A1(n_473), .A2(n_577), .B1(n_623), .B2(n_635), .Y(n_622) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g574 ( .A(n_475), .Y(n_574) );
INVx1_ASAP7_75t_L g1608 ( .A(n_475), .Y(n_1608) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .C(n_484), .Y(n_476) );
INVx1_ASAP7_75t_L g584 ( .A(n_479), .Y(n_584) );
BUFx2_ASAP7_75t_SL g984 ( .A(n_479), .Y(n_984) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_480), .Y(n_523) );
INVx2_ASAP7_75t_SL g651 ( .A(n_480), .Y(n_651) );
BUFx3_ASAP7_75t_L g701 ( .A(n_480), .Y(n_701) );
INVx1_ASAP7_75t_L g788 ( .A(n_480), .Y(n_788) );
INVx1_ASAP7_75t_L g1228 ( .A(n_480), .Y(n_1228) );
AND2x4_ASAP7_75t_L g1593 ( .A(n_480), .B(n_1594), .Y(n_1593) );
INVx2_ASAP7_75t_SL g581 ( .A(n_482), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_483), .A2(n_563), .B1(n_1562), .B2(n_1568), .Y(n_1588) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_484), .B(n_822), .C(n_825), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_484), .B(n_846), .C(n_848), .Y(n_845) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_484), .B(n_913), .C(n_915), .Y(n_912) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_484), .B(n_960), .C(n_961), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g1124 ( .A(n_484), .B(n_1125), .C(n_1126), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_484), .B(n_1216), .C(n_1217), .Y(n_1215) );
INVx2_ASAP7_75t_SL g1604 ( .A(n_485), .Y(n_1604) );
AND2x4_ASAP7_75t_L g1595 ( .A(n_486), .B(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g585 ( .A(n_487), .Y(n_585) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
XNOR2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_512), .B1(n_514), .B2(n_527), .C(n_530), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .C(n_507), .D(n_511), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_501), .B2(n_502), .C1(n_504), .C2(n_505), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_498), .A2(n_789), .B1(n_790), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_498), .A2(n_799), .B1(n_884), .B2(n_885), .Y(n_924) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x4_ASAP7_75t_L g722 ( .A(n_499), .B(n_500), .Y(n_722) );
AND2x4_ASAP7_75t_L g1626 ( .A(n_499), .B(n_1624), .Y(n_1626) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g555 ( .A(n_503), .Y(n_555) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_503), .B(n_1572), .Y(n_1579) );
AOI222xp33_ASAP7_75t_L g882 ( .A1(n_505), .A2(n_544), .B1(n_722), .B2(n_883), .C1(n_884), .C2(n_885), .Y(n_882) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_511), .B(n_720), .C(n_723), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g878 ( .A(n_511), .B(n_879), .C(n_882), .D(n_886), .Y(n_878) );
NAND3xp33_ASAP7_75t_SL g1141 ( .A(n_511), .B(n_1142), .C(n_1145), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1534 ( .A(n_511), .B(n_1535), .C(n_1536), .Y(n_1534) );
OAI31xp33_ASAP7_75t_SL g658 ( .A1(n_512), .A2(n_659), .A3(n_661), .B(n_665), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_512), .A2(n_719), .B(n_726), .Y(n_718) );
OAI31xp33_ASAP7_75t_L g795 ( .A1(n_512), .A2(n_796), .A3(n_797), .B(n_801), .Y(n_795) );
OAI31xp33_ASAP7_75t_SL g850 ( .A1(n_512), .A2(n_851), .A3(n_852), .B(n_859), .Y(n_850) );
AOI221x1_ASAP7_75t_L g877 ( .A1(n_512), .A2(n_878), .B1(n_889), .B2(n_899), .C(n_900), .Y(n_877) );
OAI31xp33_ASAP7_75t_L g918 ( .A1(n_512), .A2(n_919), .A3(n_920), .B(n_925), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g1140 ( .A1(n_512), .A2(n_1141), .B(n_1148), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_512), .A2(n_529), .B1(n_1177), .B2(n_1188), .C(n_1198), .Y(n_1176) );
OAI21xp5_ASAP7_75t_L g1533 ( .A1(n_512), .A2(n_1534), .B(n_1538), .Y(n_1533) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
AOI31xp33_ASAP7_75t_L g741 ( .A1(n_513), .A2(n_742), .A3(n_744), .B(n_747), .Y(n_741) );
AOI31xp33_ASAP7_75t_L g964 ( .A1(n_513), .A2(n_965), .A3(n_969), .B(n_972), .Y(n_964) );
AOI31xp33_ASAP7_75t_SL g1020 ( .A1(n_513), .A2(n_1021), .A3(n_1024), .B(n_1026), .Y(n_1020) );
AOI31xp33_ASAP7_75t_L g1066 ( .A1(n_513), .A2(n_1067), .A3(n_1070), .B(n_1073), .Y(n_1066) );
AOI31xp33_ASAP7_75t_L g1093 ( .A1(n_513), .A2(n_1094), .A3(n_1097), .B(n_1100), .Y(n_1093) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_523), .A2(n_958), .B1(n_1563), .B2(n_1565), .Y(n_1589) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI31xp33_ASAP7_75t_L g978 ( .A1(n_528), .A2(n_979), .A3(n_982), .B(n_987), .Y(n_978) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AO211x2_ASAP7_75t_L g728 ( .A1(n_529), .A2(n_729), .B(n_741), .C(n_750), .Y(n_728) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_529), .Y(n_899) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_531), .B(n_548), .C(n_560), .D(n_575), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_540), .C(n_546), .Y(n_531) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_535), .B(n_1572), .Y(n_1577) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
BUFx3_ASAP7_75t_L g695 ( .A(n_538), .Y(n_695) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g610 ( .A(n_539), .Y(n_610) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_539), .Y(n_813) );
BUFx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_SL g757 ( .A(n_543), .Y(n_757) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_543), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_544), .Y(n_1190) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI33xp33_ASAP7_75t_L g1045 ( .A1(n_546), .A2(n_838), .A3(n_1046), .B1(n_1048), .B2(n_1051), .B3(n_1053), .Y(n_1045) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .C(n_556), .Y(n_548) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_555), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_556), .B(n_694), .C(n_696), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_556), .B(n_760), .C(n_763), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_556), .B(n_811), .C(n_814), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g1007 ( .A(n_556), .B(n_1008), .C(n_1010), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1111 ( .A(n_556), .B(n_1112), .C(n_1117), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_556), .B(n_1200), .C(n_1201), .Y(n_1199) );
INVx5_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx6_ASAP7_75t_L g838 ( .A(n_557), .Y(n_838) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_559), .B(n_1573), .Y(n_1572) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_566), .C(n_572), .Y(n_560) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g1120 ( .A(n_565), .Y(n_1120) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g716 ( .A(n_571), .Y(n_716) );
INVx1_ASAP7_75t_L g1060 ( .A(n_571), .Y(n_1060) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g771 ( .A(n_573), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_573), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .C(n_582), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_SL g1164 ( .A1(n_577), .A2(n_708), .B1(n_1165), .B2(n_1169), .Y(n_1164) );
OAI22xp5_ASAP7_75t_SL g1525 ( .A1(n_577), .A2(n_708), .B1(n_1526), .B2(n_1529), .Y(n_1525) );
INVx4_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx4f_ASAP7_75t_L g717 ( .A(n_578), .Y(n_717) );
BUFx4f_ASAP7_75t_L g778 ( .A(n_578), .Y(n_778) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g669 ( .A(n_586), .Y(n_669) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_643), .C(n_658), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_622), .Y(n_592) );
OAI33xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .A3(n_603), .B1(n_611), .B2(n_615), .B3(n_621), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_597), .A2(n_923), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g1561 ( .A1(n_597), .A2(n_599), .B1(n_1562), .B2(n_1563), .Y(n_1561) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_602), .B1(n_624), .B2(n_629), .C(n_633), .Y(n_623) );
INVx2_ASAP7_75t_L g1157 ( .A(n_599), .Y(n_1157) );
BUFx3_ASAP7_75t_L g1560 ( .A(n_599), .Y(n_1560) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_605), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g1567 ( .A(n_606), .Y(n_1567) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g668 ( .A(n_607), .Y(n_668) );
INVx1_ASAP7_75t_L g1159 ( .A(n_609), .Y(n_1159) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g762 ( .A(n_610), .Y(n_762) );
INVx2_ASAP7_75t_L g807 ( .A(n_610), .Y(n_807) );
INVx2_ASAP7_75t_L g1116 ( .A(n_610), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1556 ( .A(n_610), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_610), .B(n_1572), .Y(n_1582) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_620), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g1518 ( .A1(n_616), .A2(n_923), .B1(n_1519), .B2(n_1520), .Y(n_1518) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g663 ( .A(n_619), .Y(n_663) );
INVx2_ASAP7_75t_L g855 ( .A(n_619), .Y(n_855) );
INVx3_ASAP7_75t_L g923 ( .A(n_619), .Y(n_923) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g636 ( .A(n_625), .Y(n_636) );
INVx2_ASAP7_75t_L g1527 ( .A(n_625), .Y(n_1527) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g645 ( .A(n_626), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g632 ( .A(n_627), .B(n_628), .Y(n_632) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g639 ( .A(n_632), .Y(n_639) );
INVx1_ASAP7_75t_L g930 ( .A(n_632), .Y(n_930) );
INVx2_ASAP7_75t_L g1167 ( .A(n_632), .Y(n_1167) );
BUFx4f_ASAP7_75t_L g1171 ( .A(n_632), .Y(n_1171) );
INVx2_ASAP7_75t_L g704 ( .A(n_634), .Y(n_704) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_634), .Y(n_1064) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_640), .C(n_641), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_636), .A2(n_1161), .B1(n_1162), .B2(n_1166), .C(n_1168), .Y(n_1165) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_636), .A2(n_1143), .B1(n_1146), .B2(n_1170), .C(n_1172), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_638), .Y(n_1136) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g715 ( .A(n_642), .Y(n_715) );
BUFx3_ASAP7_75t_L g997 ( .A(n_642), .Y(n_997) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_654), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g819 ( .A(n_651), .Y(n_819) );
NAND4xp25_ASAP7_75t_SL g729 ( .A(n_654), .B(n_730), .C(n_733), .D(n_736), .Y(n_729) );
NAND3xp33_ASAP7_75t_SL g784 ( .A(n_654), .B(n_785), .C(n_791), .Y(n_784) );
NAND3xp33_ASAP7_75t_SL g861 ( .A(n_654), .B(n_862), .C(n_865), .Y(n_861) );
NAND4xp25_ASAP7_75t_L g1177 ( .A(n_654), .B(n_1178), .C(n_1181), .D(n_1184), .Y(n_1177) );
NAND4xp25_ASAP7_75t_L g1221 ( .A(n_654), .B(n_1222), .C(n_1225), .D(n_1231), .Y(n_1221) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
BUFx2_ASAP7_75t_L g1553 ( .A(n_668), .Y(n_1553) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_779), .Y(n_671) );
XOR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_727), .Y(n_672) );
NAND3x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_682), .C(n_718), .Y(n_674) );
AND4x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_693), .C(n_697), .D(n_709), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .C(n_691), .Y(n_683) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g816 ( .A(n_689), .Y(n_816) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_L g758 ( .A(n_690), .Y(n_758) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_690), .Y(n_1110) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g1011 ( .A(n_692), .B(n_1012), .C(n_1017), .Y(n_1011) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .C(n_707), .Y(n_697) );
INVx4_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g914 ( .A(n_700), .Y(n_914) );
INVx2_ASAP7_75t_L g1212 ( .A(n_700), .Y(n_1212) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g1004 ( .A(n_712), .Y(n_1004) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
AOI33xp33_ASAP7_75t_L g1057 ( .A1(n_717), .A2(n_1006), .A3(n_1058), .B1(n_1061), .B2(n_1062), .B3(n_1063), .Y(n_1057) );
NAND4xp25_ASAP7_75t_L g750 ( .A(n_751), .B(n_759), .C(n_764), .D(n_772), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g805 ( .A(n_754), .Y(n_805) );
INVx1_ASAP7_75t_L g1009 ( .A(n_754), .Y(n_1009) );
BUFx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g1019 ( .A(n_757), .Y(n_1019) );
INVx1_ASAP7_75t_L g1209 ( .A(n_757), .Y(n_1209) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_762), .Y(n_1106) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_768), .C(n_771), .Y(n_764) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
BUFx4f_ASAP7_75t_L g775 ( .A(n_769), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .C(n_778), .Y(n_772) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_778), .B(n_992), .C(n_996), .Y(n_991) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
XOR2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_826), .Y(n_780) );
NAND3x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_795), .C(n_802), .Y(n_782) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g864 ( .A(n_788), .Y(n_864) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AND4x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_810), .C(n_817), .D(n_821), .Y(n_802) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g831 ( .A(n_813), .Y(n_831) );
INVx2_ASAP7_75t_L g836 ( .A(n_813), .Y(n_836) );
INVx3_ASAP7_75t_L g907 ( .A(n_813), .Y(n_907) );
INVx2_ASAP7_75t_SL g953 ( .A(n_813), .Y(n_953) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_SL g841 ( .A(n_824), .Y(n_841) );
XOR2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_869), .Y(n_826) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_850), .C(n_860), .Y(n_827) );
AND4x1_ASAP7_75t_L g828 ( .A(n_829), .B(n_834), .C(n_839), .D(n_845), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_837), .C(n_838), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_838), .A2(n_1150), .B1(n_1158), .B2(n_1163), .C(n_1164), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1516 ( .A1(n_838), .A2(n_1163), .B1(n_1517), .B2(n_1521), .C(n_1525), .Y(n_1516) );
INVx1_ASAP7_75t_L g1569 ( .A(n_838), .Y(n_1569) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AO22x2_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_1077), .B1(n_1259), .B2(n_1260), .Y(n_872) );
INVx1_ASAP7_75t_L g1259 ( .A(n_873), .Y(n_1259) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_974), .Y(n_873) );
AO22x2_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B1(n_933), .B2(n_934), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g925 ( .A(n_879), .Y(n_925) );
INVx1_ASAP7_75t_L g919 ( .A(n_886), .Y(n_919) );
INVxp67_ASAP7_75t_L g927 ( .A(n_890), .Y(n_927) );
INVxp67_ASAP7_75t_L g932 ( .A(n_897), .Y(n_932) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_899), .A2(n_927), .A3(n_928), .B(n_932), .Y(n_926) );
AOI211x1_ASAP7_75t_SL g1031 ( .A1(n_899), .A2(n_1032), .B(n_1044), .C(n_1066), .Y(n_1031) );
AOI211xp5_ASAP7_75t_L g1081 ( .A1(n_899), .A2(n_1082), .B(n_1093), .C(n_1102), .Y(n_1081) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_901), .B(n_918), .C(n_926), .Y(n_917) );
AND4x1_ASAP7_75t_L g901 ( .A(n_902), .B(n_905), .C(n_909), .D(n_912), .Y(n_901) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI22xp33_ASAP7_75t_SL g1522 ( .A1(n_923), .A2(n_1153), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1601 ( .A(n_930), .Y(n_1601) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
NAND4xp25_ASAP7_75t_L g947 ( .A(n_948), .B(n_951), .C(n_955), .D(n_959), .Y(n_947) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_976), .B1(n_1029), .B2(n_1076), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
NOR3xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_990), .C(n_1020), .Y(n_977) );
NAND4xp25_ASAP7_75t_L g990 ( .A(n_991), .B(n_1002), .C(n_1007), .D(n_1011), .Y(n_990) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx2_ASAP7_75t_SL g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1128 ( .A(n_999), .Y(n_1128) );
INVx2_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
BUFx2_ASAP7_75t_L g1243 ( .A(n_1000), .Y(n_1243) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1001), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1005), .C(n_1006), .Y(n_1002) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1016), .Y(n_1206) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1029), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_1030), .A2(n_1316), .B1(n_1317), .B2(n_1318), .Y(n_1315) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1031), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1057), .Y(n_1044) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_1050), .A2(n_1565), .B1(n_1566), .B2(n_1568), .Y(n_1564) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1055), .Y(n_1144) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
AND2x4_ASAP7_75t_L g1628 ( .A(n_1056), .B(n_1624), .Y(n_1628) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1077), .Y(n_1260) );
AO22x2_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1173), .B1(n_1174), .B2(n_1258), .Y(n_1077) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1078), .Y(n_1258) );
XNOR2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1130), .Y(n_1078) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1081), .Y(n_1129) );
NAND4xp25_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1111), .C(n_1118), .D(n_1124), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1109), .B(n_1572), .Y(n_1571) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
NAND3x1_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1140), .C(n_1149), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_1152), .A2(n_1153), .B1(n_1155), .B2(n_1156), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1557 ( .A1(n_1153), .A2(n_1558), .B1(n_1559), .B2(n_1560), .Y(n_1557) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
OAI221xp5_ASAP7_75t_L g1526 ( .A1(n_1166), .A2(n_1519), .B1(n_1520), .B2(n_1527), .C(n_1528), .Y(n_1526) );
OAI221xp5_ASAP7_75t_L g1529 ( .A1(n_1166), .A2(n_1527), .B1(n_1530), .B2(n_1531), .C(n_1532), .Y(n_1529) );
BUFx3_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
OAI211xp5_ASAP7_75t_L g1605 ( .A1(n_1170), .A2(n_1559), .B(n_1606), .C(n_1607), .Y(n_1605) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_1174), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1218), .B1(n_1219), .B2(n_1257), .Y(n_1174) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1175), .Y(n_1257) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1193), .C(n_1196), .Y(n_1188) );
NAND4xp25_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1202), .C(n_1210), .D(n_1215), .Y(n_1198) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1220), .Y(n_1256) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1240), .Y(n_1234) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1502), .B1(n_1504), .B2(n_1539), .C(n_1542), .Y(n_1261) );
AOI21xp5_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1407), .B(n_1451), .Y(n_1262) );
NAND5xp2_ASAP7_75t_SL g1263 ( .A(n_1264), .B(n_1346), .C(n_1375), .D(n_1398), .E(n_1402), .Y(n_1263) );
AOI21xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1303), .B(n_1324), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1286), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1266), .B(n_1313), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1266), .B(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1266), .B(n_1335), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1266), .B(n_1313), .Y(n_1436) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1267), .B(n_1333), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1267), .B(n_1313), .Y(n_1345) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1267), .Y(n_1352) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1267), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1267), .B(n_1286), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1434 ( .A(n_1267), .B(n_1343), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1267), .B(n_1335), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1280), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1275), .Y(n_1269) );
OAI21xp33_ASAP7_75t_SL g1631 ( .A1(n_1270), .A2(n_1541), .B(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1271), .B(n_1276), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1274), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1274), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1275), .B(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1276), .B(n_1279), .Y(n_1302) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_1277), .Y(n_1308) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1281), .Y(n_1321) );
BUFx3_ASAP7_75t_L g1367 ( .A(n_1281), .Y(n_1367) );
AND2x4_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1284), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1282), .B(n_1284), .Y(n_1291) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_1283), .B(n_1284), .Y(n_1285) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1285), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1292), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1287), .B(n_1339), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1287), .B(n_1330), .Y(n_1395) );
A2O1A1Ixp33_ASAP7_75t_L g1468 ( .A1(n_1287), .A2(n_1469), .B(n_1472), .C(n_1473), .Y(n_1468) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
BUFx2_ASAP7_75t_L g1333 ( .A(n_1288), .Y(n_1333) );
BUFx3_ASAP7_75t_L g1343 ( .A(n_1288), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1288), .B(n_1330), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1290), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1292), .B(n_1333), .Y(n_1364) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1292), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1297), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1293), .B(n_1343), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1293), .B(n_1333), .Y(n_1414) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1294), .B(n_1297), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1294), .B(n_1340), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1294), .B(n_1343), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1294), .B(n_1297), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1386 ( .A(n_1294), .B(n_1343), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1296), .Y(n_1294) );
INVx2_ASAP7_75t_SL g1340 ( .A(n_1297), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1297), .B(n_1343), .Y(n_1360) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1301), .B2(n_1302), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g1316 ( .A(n_1300), .Y(n_1316) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1302), .Y(n_1319) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1303), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1312), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1304), .B(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1304), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1304), .B(n_1405), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1304), .B(n_1313), .Y(n_1440) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1305), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1305), .B(n_1325), .Y(n_1488) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1306), .B(n_1325), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1306), .B(n_1336), .Y(n_1383) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1306), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1309), .Y(n_1306) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_1311), .A2(n_1321), .B1(n_1322), .B2(n_1323), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1312), .B(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1312), .Y(n_1450) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1313), .B(n_1325), .Y(n_1353) );
INVx2_ASAP7_75t_SL g1389 ( .A(n_1313), .Y(n_1389) );
AND2x4_ASAP7_75t_L g1405 ( .A(n_1313), .B(n_1336), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g1442 ( .A(n_1313), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g1313 ( .A(n_1314), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1314), .B(n_1336), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1314), .B(n_1325), .Y(n_1397) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1320), .Y(n_1314) );
BUFx3_ASAP7_75t_L g1370 ( .A(n_1316), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_1318), .Y(n_1372) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
OAI211xp5_ASAP7_75t_SL g1324 ( .A1(n_1325), .A2(n_1328), .B(n_1334), .C(n_1341), .Y(n_1324) );
INVx3_ASAP7_75t_L g1336 ( .A(n_1325), .Y(n_1336) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1325), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1327), .Y(n_1325) );
OAI321xp33_ASAP7_75t_L g1433 ( .A1(n_1328), .A2(n_1348), .A3(n_1379), .B1(n_1427), .B2(n_1434), .C(n_1435), .Y(n_1433) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1329), .B(n_1389), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1329), .B(n_1480), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1332), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1330), .B(n_1359), .Y(n_1444) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_1331), .B(n_1434), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1332), .B(n_1379), .Y(n_1465) );
NOR2x1_ASAP7_75t_L g1432 ( .A(n_1333), .B(n_1340), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1333), .B(n_1379), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1337), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_1335), .A2(n_1409), .B1(n_1411), .B2(n_1417), .C(n_1418), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1336), .B(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1336), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1336), .B(n_1463), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_1336), .A2(n_1380), .B1(n_1478), .B2(n_1481), .C(n_1484), .Y(n_1477) );
O2A1O1Ixp33_ASAP7_75t_L g1421 ( .A1(n_1337), .A2(n_1404), .B(n_1422), .C(n_1424), .Y(n_1421) );
AOI222xp33_ASAP7_75t_L g1458 ( .A1(n_1337), .A2(n_1383), .B1(n_1459), .B2(n_1461), .C1(n_1464), .C2(n_1466), .Y(n_1458) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1338), .B(n_1351), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1339), .B(n_1343), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1339), .B(n_1352), .Y(n_1419) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1339), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1340), .B(n_1343), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1344), .Y(n_1341) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1342), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1342), .B(n_1359), .Y(n_1499) );
OR2x2_ASAP7_75t_L g1377 ( .A(n_1343), .B(n_1378), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1343), .B(n_1392), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1343), .B(n_1444), .Y(n_1472) );
O2A1O1Ixp33_ASAP7_75t_L g1484 ( .A1(n_1345), .A2(n_1485), .B(n_1486), .C(n_1487), .Y(n_1484) );
A2O1A1Ixp33_ASAP7_75t_L g1346 ( .A1(n_1347), .A2(n_1349), .B(n_1354), .C(n_1373), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1348), .B(n_1377), .Y(n_1376) );
O2A1O1Ixp33_ASAP7_75t_L g1418 ( .A1(n_1348), .A2(n_1352), .B(n_1419), .C(n_1420), .Y(n_1418) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1348), .B(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1353), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1351), .B(n_1386), .Y(n_1423) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1351), .B(n_1432), .Y(n_1431) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
AOI321xp33_ASAP7_75t_L g1375 ( .A1(n_1352), .A2(n_1376), .A3(n_1380), .B1(n_1382), .B2(n_1384), .C(n_1393), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1352), .B(n_1397), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1352), .B(n_1414), .Y(n_1413) );
NAND2xp5_ASAP7_75t_SL g1448 ( .A(n_1352), .B(n_1386), .Y(n_1448) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1353), .Y(n_1416) );
OAI211xp5_ASAP7_75t_SL g1354 ( .A1(n_1355), .A2(n_1357), .B(n_1361), .C(n_1365), .Y(n_1354) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_1355), .A2(n_1412), .B1(n_1415), .B2(n_1416), .Y(n_1411) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
A2O1A1Ixp33_ASAP7_75t_L g1446 ( .A1(n_1356), .A2(n_1447), .B(n_1449), .C(n_1450), .Y(n_1446) );
AOI31xp33_ASAP7_75t_L g1497 ( .A1(n_1357), .A2(n_1394), .A3(n_1498), .B(n_1500), .Y(n_1497) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1360), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1359), .B(n_1379), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1359), .B(n_1389), .Y(n_1494) );
INVxp67_ASAP7_75t_L g1415 ( .A(n_1360), .Y(n_1415) );
INVxp67_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .Y(n_1362) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1365), .Y(n_1445) );
INVx3_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx3_ASAP7_75t_L g1374 ( .A(n_1366), .Y(n_1374) );
OAI22xp33_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .B1(n_1371), .B2(n_1372), .Y(n_1368) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1370), .Y(n_1503) );
AOI21xp5_ASAP7_75t_L g1393 ( .A1(n_1378), .A2(n_1394), .B(n_1396), .Y(n_1393) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1380), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1381), .B(n_1389), .Y(n_1388) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1387), .B1(n_1390), .B2(n_1391), .Y(n_1384) );
INVxp33_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1389), .B(n_1430), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1456 ( .A(n_1389), .B(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1389), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1389), .B(n_1483), .Y(n_1482) );
NOR2xp33_ASAP7_75t_L g1501 ( .A(n_1389), .B(n_1462), .Y(n_1501) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1390), .Y(n_1417) );
A2O1A1Ixp33_ASAP7_75t_L g1426 ( .A1(n_1390), .A2(n_1427), .B(n_1428), .C(n_1433), .Y(n_1426) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_1395), .B(n_1401), .Y(n_1496) );
AOI221xp5_ASAP7_75t_L g1437 ( .A1(n_1397), .A2(n_1406), .B1(n_1438), .B2(n_1439), .C(n_1441), .Y(n_1437) );
CKINVDCx5p33_ASAP7_75t_R g1476 ( .A(n_1397), .Y(n_1476) );
INVxp67_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVxp67_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1406), .Y(n_1403) );
NAND5xp2_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1421), .C(n_1426), .D(n_1437), .E(n_1446), .Y(n_1407) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1452 ( .A1(n_1417), .A2(n_1453), .B1(n_1455), .B2(n_1456), .Y(n_1452) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1425), .Y(n_1490) );
INVxp67_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1438), .Y(n_1486) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
OAI21xp33_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1443), .B(n_1445), .Y(n_1441) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_1442), .B(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
NAND5xp2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1458), .C(n_1468), .D(n_1477), .E(n_1489), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1454), .Y(n_1475) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1454), .Y(n_1493) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1471), .Y(n_1469) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1476), .Y(n_1474) );
INVxp67_ASAP7_75t_SL g1478 ( .A(n_1479), .Y(n_1478) );
INVxp67_ASAP7_75t_SL g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
O2A1O1Ixp33_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1491), .B(n_1495), .C(n_1497), .Y(n_1489) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVxp67_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
NAND3x1_ASAP7_75t_SL g1507 ( .A(n_1508), .B(n_1516), .C(n_1533), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_1540), .Y(n_1539) );
BUFx3_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
BUFx2_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_SL g1629 ( .A(n_1549), .Y(n_1629) );
NAND4xp75_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1574), .C(n_1586), .D(n_1621), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1553), .B1(n_1554), .B2(n_1555), .Y(n_1551) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
BUFx2_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
NOR2x1_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1580), .Y(n_1574) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVxp67_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx2_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx3_ASAP7_75t_L g1624 ( .A(n_1584), .Y(n_1624) );
OAI31xp33_ASAP7_75t_L g1586 ( .A1(n_1587), .A2(n_1597), .A3(n_1609), .B(n_1620), .Y(n_1586) );
A2O1A1Ixp33_ASAP7_75t_L g1587 ( .A1(n_1588), .A2(n_1589), .B(n_1590), .C(n_1592), .Y(n_1587) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1591), .Y(n_1596) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
BUFx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND2x4_ASAP7_75t_L g1611 ( .A(n_1595), .B(n_1612), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1595), .B(n_1616), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1605), .Y(n_1597) );
OAI211xp5_ASAP7_75t_L g1598 ( .A1(n_1599), .A2(n_1600), .B(n_1602), .C(n_1603), .Y(n_1598) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1611), .Y(n_1610) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx3_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1619), .Y(n_1617) );
AOI221xp5_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1625), .B1(n_1626), .B2(n_1627), .C(n_1628), .Y(n_1621) );
AND2x4_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
HB1xp67_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
endmodule