module fake_netlist_6_4760_n_1843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1843;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_110),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_17),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_39),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_73),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_106),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_33),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_105),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_100),
.Y(n_205)
);

INVx4_ASAP7_75t_R g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_37),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_71),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_86),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_57),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_60),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_98),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_39),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_42),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_163),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_58),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_84),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_6),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_38),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_162),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_40),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_47),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_135),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_180),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_114),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_129),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_109),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_7),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_95),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_53),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_61),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_68),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_115),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_155),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_42),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_107),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_64),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_141),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_57),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_87),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_19),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_19),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_22),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_32),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_148),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_158),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_45),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_165),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_149),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_92),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_131),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_173),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_34),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_67),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_96),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_31),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_63),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_82),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_10),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_125),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_28),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_120),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_123),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_74),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_36),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_181),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_38),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_33),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_26),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_21),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_1),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_124),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_36),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_34),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_136),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_182),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_116),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_8),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_20),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_49),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_46),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_14),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_79),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_147),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_145),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_127),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_5),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_8),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_44),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_66),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_70),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_15),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_30),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_81),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_49),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_146),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_16),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_43),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_2),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_6),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_169),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_59),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_101),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_43),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_133),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_29),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_137),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_99),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_121),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_83),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_11),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_3),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_164),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_12),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_91),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_185),
.B(n_0),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_240),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_R g371 ( 
.A(n_248),
.B(n_113),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_0),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_240),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_212),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_212),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_212),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_283),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_230),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_238),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_237),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_285),
.B(n_3),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_339),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_301),
.B(n_4),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_4),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_252),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_212),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_253),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_255),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_241),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_239),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_210),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_188),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_239),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_256),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_273),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_239),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_271),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_239),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_261),
.B(n_239),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_301),
.B(n_5),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_264),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_188),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_219),
.B(n_7),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_264),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_288),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_244),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_197),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_288),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_219),
.B(n_12),
.Y(n_412)
);

BUFx2_ASAP7_75t_SL g413 ( 
.A(n_323),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_202),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_228),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_231),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_245),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_233),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_275),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_282),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_309),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_232),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_336),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_208),
.B(n_14),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_246),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_242),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_208),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_243),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_249),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_268),
.B(n_15),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_298),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_359),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_284),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_261),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_257),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_258),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_287),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_259),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_265),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_260),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_267),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_193),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_266),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_270),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_278),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_193),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_286),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_302),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_314),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_324),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_292),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_268),
.B(n_16),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_326),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_272),
.B(n_72),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_375),
.A2(n_377),
.B(n_376),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_377),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_336),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_413),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_372),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_425),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_431),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_432),
.Y(n_481)
);

XNOR2x2_ASAP7_75t_L g482 ( 
.A(n_383),
.B(n_236),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_194),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_441),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_381),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_443),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_382),
.B(n_200),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_448),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_449),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_391),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_382),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_408),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_387),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_393),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_397),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_387),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_440),
.B(n_261),
.Y(n_504)
);

BUFx8_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_389),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_389),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_421),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_414),
.B(n_201),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_390),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_454),
.B(n_334),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_390),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_R g515 ( 
.A(n_396),
.B(n_274),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_396),
.B(n_213),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_380),
.B(n_207),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_399),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_422),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_422),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_384),
.B(n_217),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_373),
.B(n_404),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_419),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_370),
.B(n_335),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_222),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_423),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_430),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_439),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_439),
.B(n_186),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_445),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_515),
.B(n_489),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_472),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_513),
.A2(n_402),
.B1(n_385),
.B2(n_367),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_510),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_476),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_469),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_482),
.A2(n_412),
.B1(n_460),
.B2(n_434),
.Y(n_546)
);

BUFx6f_ASAP7_75t_SL g547 ( 
.A(n_469),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_502),
.B(n_405),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_519),
.A2(n_401),
.B1(n_386),
.B2(n_369),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_513),
.B(n_450),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_463),
.B(n_445),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_524),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_498),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_531),
.B(n_459),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_470),
.B(n_363),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_530),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_470),
.B(n_363),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_502),
.B(n_360),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_532),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_503),
.B(n_360),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_363),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_529),
.B(n_524),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_528),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_528),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_360),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_466),
.B(n_459),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_536),
.B(n_374),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_471),
.B(n_360),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_468),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_472),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_494),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_497),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_466),
.B(n_371),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_517),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_487),
.B(n_403),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_478),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_471),
.B(n_360),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_480),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_471),
.B(n_360),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_472),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_464),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_482),
.A2(n_427),
.B1(n_342),
.B2(n_341),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_493),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_500),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_493),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_516),
.B(n_406),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_474),
.B(n_300),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_474),
.B(n_407),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_475),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_523),
.A2(n_357),
.B1(n_364),
.B2(n_458),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_474),
.B(n_410),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_476),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_499),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_411),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_464),
.B(n_415),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_465),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_501),
.Y(n_616)
);

AND3x1_ASAP7_75t_L g617 ( 
.A(n_483),
.B(n_451),
.C(n_447),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_534),
.A2(n_456),
.B1(n_453),
.B2(n_458),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_534),
.B(n_363),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_505),
.A2(n_457),
.B1(n_456),
.B2(n_455),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_514),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_505),
.B(n_229),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_504),
.B(n_409),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_473),
.B(n_462),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_505),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_501),
.B(n_452),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_473),
.B(n_234),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_506),
.B(n_461),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_506),
.B(n_247),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_507),
.B(n_512),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_507),
.B(n_453),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_520),
.B(n_186),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_520),
.B(n_250),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_537),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_521),
.B(n_251),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_477),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_521),
.B(n_198),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_522),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_522),
.B(n_204),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_533),
.B(n_254),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_533),
.Y(n_645)
);

NAND2x1p5_ASAP7_75t_L g646 ( 
.A(n_508),
.B(n_220),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_535),
.B(n_187),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_535),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_537),
.B(n_262),
.Y(n_649)
);

BUFx8_ASAP7_75t_SL g650 ( 
.A(n_492),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_363),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_508),
.B(n_455),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_495),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_479),
.Y(n_655)
);

AND2x2_ASAP7_75t_SL g656 ( 
.A(n_479),
.B(n_263),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_481),
.B(n_457),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_481),
.B(n_269),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_484),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_484),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_291),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_488),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_490),
.B(n_295),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_490),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_491),
.B(n_430),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_491),
.B(n_433),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_509),
.B(n_294),
.C(n_293),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_510),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_515),
.B(n_187),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_472),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_469),
.B(n_433),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_469),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_482),
.A2(n_303),
.B1(n_297),
.B2(n_306),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_510),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_487),
.B(n_435),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_487),
.B(n_435),
.Y(n_677)
);

BUFx8_ASAP7_75t_SL g678 ( 
.A(n_475),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_513),
.B(n_436),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_519),
.B(n_189),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_524),
.A2(n_322),
.B1(n_308),
.B2(n_318),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_515),
.B(n_189),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_307),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_472),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_500),
.B(n_289),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_541),
.A2(n_332),
.B1(n_296),
.B2(n_367),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_601),
.A2(n_312),
.B(n_328),
.C(n_366),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_561),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_593),
.A2(n_313),
.B(n_362),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_610),
.B(n_355),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_671),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_610),
.B(n_356),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_569),
.B(n_190),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_653),
.B(n_276),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_593),
.B(n_361),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_671),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_552),
.B(n_213),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_650),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_548),
.B(n_235),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_330),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_542),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_558),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_546),
.A2(n_203),
.B1(n_368),
.B2(n_225),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_612),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_557),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_612),
.A2(n_304),
.B(n_277),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_549),
.B(n_279),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_546),
.B(n_316),
.C(n_305),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_571),
.B(n_280),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_578),
.B(n_281),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_588),
.B(n_290),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_633),
.B(n_436),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_559),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_545),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_678),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_550),
.B(n_191),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_590),
.B(n_299),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_561),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_627),
.B(n_215),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_564),
.Y(n_723)
);

BUFx8_ASAP7_75t_L g724 ( 
.A(n_555),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_R g725 ( 
.A(n_544),
.B(n_191),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_622),
.B(n_192),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_600),
.B(n_311),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_622),
.B(n_315),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_665),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_560),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_565),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_609),
.B(n_321),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_613),
.B(n_192),
.Y(n_733)
);

AND2x6_ASAP7_75t_SL g734 ( 
.A(n_632),
.B(n_437),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_613),
.B(n_195),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_631),
.B(n_195),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_541),
.B(n_203),
.C(n_368),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_564),
.Y(n_738)
);

AND3x1_ASAP7_75t_L g739 ( 
.A(n_673),
.B(n_444),
.C(n_438),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_631),
.B(n_196),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_673),
.A2(n_345),
.B1(n_216),
.B2(n_226),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_566),
.B(n_196),
.Y(n_742)
);

INVx8_ASAP7_75t_L g743 ( 
.A(n_653),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_668),
.B(n_199),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_554),
.A2(n_199),
.B1(n_209),
.B2(n_358),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_545),
.B(n_437),
.Y(n_746)
);

O2A1O1Ixp5_ASAP7_75t_L g747 ( 
.A1(n_602),
.A2(n_683),
.B(n_607),
.C(n_603),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_674),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_205),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_602),
.B(n_209),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_211),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_557),
.B(n_211),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_628),
.A2(n_630),
.B1(n_663),
.B2(n_658),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_636),
.B(n_214),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_657),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_557),
.B(n_214),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_557),
.B(n_218),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_603),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_545),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_657),
.B(n_444),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_611),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_615),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_595),
.A2(n_348),
.B1(n_365),
.B2(n_215),
.Y(n_763)
);

BUFx8_ASAP7_75t_L g764 ( 
.A(n_637),
.Y(n_764)
);

INVx6_ASAP7_75t_L g765 ( 
.A(n_653),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_557),
.B(n_221),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_562),
.B(n_221),
.Y(n_767)
);

O2A1O1Ixp5_ASAP7_75t_L g768 ( 
.A1(n_683),
.A2(n_438),
.B(n_206),
.C(n_358),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_605),
.B(n_642),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_562),
.B(n_224),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_572),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_640),
.B(n_319),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_338),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_643),
.A2(n_338),
.B(n_354),
.C(n_224),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_636),
.B(n_225),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_562),
.B(n_227),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_554),
.B(n_227),
.Y(n_777)
);

O2A1O1Ixp5_ASAP7_75t_L g778 ( 
.A1(n_577),
.A2(n_343),
.B(n_354),
.C(n_344),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_585),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_562),
.B(n_327),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_629),
.B(n_327),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_586),
.B(n_343),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_639),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_585),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_672),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_586),
.B(n_329),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_638),
.B(n_329),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_638),
.B(n_344),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_587),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_658),
.A2(n_337),
.B1(n_349),
.B2(n_320),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_644),
.B(n_337),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_644),
.B(n_349),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_585),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_672),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_666),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_649),
.B(n_365),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_592),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_649),
.A2(n_352),
.B(n_351),
.C(n_350),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_677),
.B(n_352),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_577),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_543),
.B(n_351),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_543),
.B(n_350),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_589),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_666),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_625),
.B(n_348),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_573),
.B(n_346),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_679),
.B(n_635),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_658),
.A2(n_346),
.B1(n_345),
.B2(n_340),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_619),
.B(n_340),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_658),
.A2(n_333),
.B1(n_331),
.B2(n_325),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_573),
.B(n_333),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_647),
.B(n_331),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_672),
.B(n_325),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_539),
.B(n_226),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_656),
.B(n_216),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_582),
.B(n_77),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_553),
.B(n_21),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_580),
.B(n_23),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_582),
.B(n_538),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_592),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_540),
.B(n_78),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_589),
.Y(n_824)
);

INVx8_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_591),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_591),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_663),
.A2(n_85),
.B1(n_177),
.B2(n_167),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_592),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_563),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_556),
.B(n_575),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_608),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_579),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_581),
.B(n_25),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_680),
.B(n_25),
.C(n_27),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_596),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_563),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_583),
.B(n_27),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_599),
.B(n_69),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_667),
.B(n_28),
.C(n_29),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_656),
.B(n_93),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_604),
.B(n_90),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_623),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_632),
.B(n_30),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_670),
.A2(n_684),
.B(n_567),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_568),
.B(n_626),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_SL g848 ( 
.A(n_708),
.B(n_641),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_761),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_707),
.B(n_663),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_831),
.A2(n_663),
.B1(n_648),
.B2(n_584),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_821),
.A2(n_570),
.B(n_597),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_802),
.A2(n_570),
.B(n_597),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_753),
.B(n_637),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_805),
.A2(n_826),
.B(n_824),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_762),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_832),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_717),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_755),
.B(n_645),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_827),
.A2(n_570),
.B(n_597),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_841),
.A2(n_574),
.B(n_624),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_723),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_704),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_693),
.B(n_637),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_797),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_830),
.A2(n_570),
.B(n_594),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_837),
.A2(n_597),
.B(n_594),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_784),
.B(n_655),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_747),
.A2(n_778),
.B(n_735),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_703),
.B(n_685),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_729),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_735),
.A2(n_595),
.B(n_682),
.C(n_669),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_807),
.B(n_654),
.C(n_659),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_758),
.B(n_651),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_797),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_845),
.A2(n_624),
.B(n_620),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_709),
.A2(n_594),
.B(n_618),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_698),
.A2(n_594),
.B(n_618),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_807),
.B(n_817),
.C(n_686),
.Y(n_879)
);

BUFx8_ASAP7_75t_L g880 ( 
.A(n_701),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_846),
.A2(n_617),
.B(n_681),
.Y(n_881)
);

OR2x6_ASAP7_75t_SL g882 ( 
.A(n_718),
.B(n_664),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_747),
.A2(n_568),
.B(n_606),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_736),
.B(n_651),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_790),
.B(n_736),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_733),
.A2(n_627),
.B(n_652),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_702),
.A2(n_652),
.B(n_606),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_710),
.A2(n_738),
.B(n_723),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_836),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_740),
.B(n_651),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_738),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_831),
.B(n_634),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_740),
.B(n_660),
.C(n_662),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_754),
.B(n_651),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_688),
.A2(n_661),
.B(n_568),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_651),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_841),
.A2(n_568),
.B1(n_661),
.B2(n_547),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_790),
.B(n_662),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_689),
.A2(n_661),
.B(n_568),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_806),
.B(n_616),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_717),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_690),
.A2(n_655),
.B(n_646),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_721),
.A2(n_646),
.B(n_621),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_823),
.A2(n_621),
.B(n_547),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_809),
.A2(n_775),
.B1(n_772),
.B2(n_779),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_750),
.A2(n_621),
.B(n_117),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_775),
.B(n_634),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_746),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_819),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_760),
.B(n_616),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_717),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_801),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_782),
.B(n_715),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_809),
.A2(n_614),
.B1(n_598),
.B2(n_621),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_818),
.A2(n_621),
.B(n_102),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_792),
.B(n_614),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_843),
.B(n_700),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_771),
.A2(n_94),
.B(n_179),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_746),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_737),
.A2(n_598),
.B1(n_35),
.B2(n_37),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_833),
.Y(n_921)
);

O2A1O1Ixp5_ASAP7_75t_L g922 ( 
.A1(n_768),
.A2(n_150),
.B(n_139),
.C(n_134),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_793),
.B(n_692),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_778),
.A2(n_126),
.B(n_119),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_817),
.B(n_31),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_695),
.B(n_35),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_814),
.B(n_41),
.C(n_46),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_800),
.A2(n_41),
.B(n_47),
.C(n_50),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_705),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_751),
.B(n_788),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_686),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_814),
.B(n_51),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_693),
.B(n_104),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_716),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_787),
.B(n_118),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_717),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_730),
.B(n_52),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_788),
.B(n_53),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_796),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_54),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_789),
.B(n_798),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_719),
.A2(n_748),
.B1(n_783),
.B2(n_777),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_796),
.B(n_838),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_789),
.B(n_691),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_838),
.A2(n_737),
.B(n_774),
.C(n_768),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_741),
.A2(n_763),
.B1(n_711),
.B2(n_810),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_712),
.A2(n_732),
.B(n_714),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_836),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_836),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_811),
.B(n_777),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_759),
.B(n_803),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_791),
.A2(n_728),
.B(n_694),
.C(n_699),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_713),
.A2(n_720),
.B(n_727),
.Y(n_953)
);

AO22x1_ASAP7_75t_L g954 ( 
.A1(n_840),
.A2(n_706),
.B1(n_764),
.B2(n_834),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_728),
.A2(n_842),
.B(n_839),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_786),
.B(n_796),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_804),
.B(n_808),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_780),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_813),
.B(n_796),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_741),
.A2(n_763),
.B1(n_812),
.B2(n_835),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_742),
.B(n_744),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_785),
.A2(n_795),
.B(n_799),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_687),
.A2(n_783),
.B(n_770),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_752),
.A2(n_766),
.B(n_773),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_693),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_811),
.B(n_816),
.Y(n_966)
);

OAI321xp33_ASAP7_75t_L g967 ( 
.A1(n_726),
.A2(n_820),
.A3(n_828),
.B1(n_844),
.B2(n_745),
.C(n_696),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_822),
.A2(n_829),
.B(n_757),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_725),
.B(n_765),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_840),
.A2(n_749),
.B(n_781),
.C(n_776),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_836),
.B(n_708),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_756),
.A2(n_767),
.B(n_825),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_725),
.B(n_765),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_815),
.A2(n_847),
.B(n_697),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_794),
.A2(n_825),
.B(n_708),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_739),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_708),
.B(n_794),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_765),
.B(n_734),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_708),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_722),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_764),
.B(n_724),
.C(n_769),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_743),
.B(n_769),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_743),
.A2(n_735),
.B(n_841),
.C(n_800),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_724),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_707),
.A2(n_747),
.B(n_593),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_753),
.B(n_554),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_707),
.A2(n_593),
.B(n_821),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_707),
.B(n_758),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_764),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_761),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_735),
.A2(n_841),
.B(n_800),
.C(n_703),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_729),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_698),
.A2(n_821),
.B(n_613),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_707),
.A2(n_593),
.B(n_821),
.Y(n_994)
);

CKINVDCx10_ASAP7_75t_R g995 ( 
.A(n_769),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_761),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_707),
.A2(n_593),
.B(n_821),
.Y(n_997)
);

BUFx12f_ASAP7_75t_L g998 ( 
.A(n_764),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_762),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_707),
.B(n_758),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_717),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_707),
.A2(n_747),
.B(n_593),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_845),
.A2(n_747),
.B(n_821),
.Y(n_1003)
);

OAI321xp33_ASAP7_75t_L g1004 ( 
.A1(n_686),
.A2(n_546),
.A3(n_673),
.B1(n_541),
.B2(n_595),
.C(n_711),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_794),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_707),
.B(n_758),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_761),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_753),
.B(n_554),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_707),
.B(n_758),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_753),
.B(n_554),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_707),
.A2(n_747),
.B(n_593),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_786),
.B(n_759),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_761),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_786),
.B(n_759),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_755),
.B(n_790),
.Y(n_1016)
);

AND2x6_ASAP7_75t_L g1017 ( 
.A(n_802),
.B(n_805),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_836),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_735),
.A2(n_841),
.B(n_800),
.C(n_703),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_1003),
.A2(n_968),
.B(n_888),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_905),
.B(n_991),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_885),
.A2(n_925),
.B(n_879),
.C(n_1004),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_993),
.A2(n_877),
.B(n_850),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_972),
.A2(n_904),
.B(n_971),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_857),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_871),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1004),
.A2(n_930),
.B(n_946),
.C(n_1019),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_913),
.B(n_988),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_992),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_985),
.A2(n_1011),
.B(n_1002),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_863),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_908),
.B(n_934),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1016),
.B(n_917),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_SL g1035 ( 
.A(n_1005),
.B(n_864),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_971),
.A2(n_975),
.B(n_979),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_865),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_910),
.B(n_923),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_875),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_979),
.A2(n_852),
.B(n_977),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_961),
.B(n_907),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_987),
.A2(n_997),
.B(n_994),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_957),
.B(n_898),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_946),
.A2(n_950),
.B(n_960),
.C(n_872),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_874),
.A2(n_890),
.B(n_884),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_1013),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_SL g1047 ( 
.A1(n_985),
.A2(n_1011),
.B(n_1002),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_932),
.B(n_976),
.Y(n_1048)
);

AOI221xp5_ASAP7_75t_SL g1049 ( 
.A1(n_960),
.A2(n_931),
.B1(n_912),
.B2(n_920),
.C(n_881),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_980),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_944),
.A2(n_942),
.B1(n_986),
.B2(n_1010),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_929),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_911),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_869),
.A2(n_955),
.B(n_883),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_977),
.A2(n_962),
.B(n_876),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_853),
.A2(n_860),
.B(n_866),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_849),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_966),
.A2(n_967),
.B(n_887),
.C(n_938),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_869),
.A2(n_883),
.B(n_945),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_911),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_952),
.A2(n_896),
.A3(n_894),
.B(n_926),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_963),
.A2(n_924),
.B(n_955),
.C(n_854),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1008),
.A2(n_851),
.B1(n_893),
.B2(n_943),
.Y(n_1063)
);

AOI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_970),
.A2(n_870),
.B(n_859),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_1013),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_867),
.A2(n_964),
.B(n_878),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_909),
.B(n_916),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_990),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_909),
.B(n_941),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_963),
.A2(n_922),
.B(n_983),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_959),
.A2(n_951),
.B(n_953),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_899),
.B(n_924),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_947),
.A2(n_1005),
.B(n_901),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_1015),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_889),
.A2(n_1018),
.B(n_948),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_886),
.A2(n_935),
.B(n_928),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_911),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_996),
.B(n_1014),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_903),
.A2(n_974),
.B(n_902),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_967),
.A2(n_940),
.B(n_937),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_892),
.B(n_954),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_956),
.A2(n_1015),
.B(n_982),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_SL g1083 ( 
.A(n_873),
.B(n_927),
.C(n_914),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_L g1084 ( 
.A1(n_958),
.A2(n_891),
.B(n_862),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_921),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1007),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_889),
.A2(n_948),
.B(n_949),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_858),
.A2(n_919),
.B(n_956),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_858),
.A2(n_939),
.B(n_936),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1012),
.B(n_1017),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1017),
.B(n_856),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_918),
.B(n_906),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_868),
.B(n_973),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_999),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1017),
.B(n_969),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_880),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_936),
.B(n_939),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1017),
.B(n_897),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_900),
.A2(n_848),
.B(n_931),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_978),
.A2(n_864),
.B(n_981),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_936),
.A2(n_1001),
.B1(n_939),
.B2(n_933),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1001),
.A2(n_984),
.B(n_864),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1001),
.A2(n_965),
.B(n_989),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_965),
.A2(n_882),
.B(n_995),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_965),
.A2(n_861),
.A3(n_945),
.B(n_952),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_880),
.A2(n_709),
.B(n_869),
.C(n_963),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_998),
.A2(n_1003),
.B(n_904),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_885),
.A2(n_807),
.B(n_755),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_885),
.B(n_913),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_855),
.A2(n_707),
.B(n_593),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1016),
.B(n_755),
.Y(n_1111)
);

INVx6_ASAP7_75t_L g1112 ( 
.A(n_965),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_862),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_855),
.A2(n_707),
.B(n_593),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_988),
.A2(n_1006),
.B1(n_1009),
.B2(n_1000),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_885),
.B(n_913),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_855),
.A2(n_707),
.B(n_593),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_885),
.A2(n_925),
.B(n_879),
.C(n_1004),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_885),
.B(n_913),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_885),
.B(n_913),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1016),
.B(n_755),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_885),
.A2(n_755),
.B(n_946),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1016),
.B(n_755),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_885),
.B(n_913),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1016),
.B(n_755),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_988),
.A2(n_1006),
.B1(n_1009),
.B2(n_1000),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_885),
.B(n_913),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_993),
.A2(n_877),
.B(n_850),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_857),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_885),
.B(n_913),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_885),
.A2(n_925),
.B(n_879),
.C(n_1004),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_885),
.B(n_913),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_885),
.B(n_913),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_861),
.A2(n_945),
.A3(n_952),
.B(n_960),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1003),
.A2(n_968),
.B(n_845),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_993),
.A2(n_877),
.B(n_850),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_885),
.B(n_913),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_885),
.B(n_913),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1016),
.B(n_755),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_857),
.B(n_832),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_998),
.B(n_693),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_855),
.A2(n_1019),
.B(n_991),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1016),
.B(n_755),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_885),
.B(n_913),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1016),
.B(n_755),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_993),
.A2(n_877),
.B(n_850),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_885),
.B(n_913),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_862),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1003),
.A2(n_968),
.B(n_845),
.Y(n_1149)
);

AOI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_885),
.A2(n_755),
.B(n_946),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_863),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1003),
.A2(n_968),
.B(n_845),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_855),
.A2(n_1019),
.B(n_991),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_863),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_885),
.A2(n_925),
.B(n_879),
.C(n_1004),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1003),
.A2(n_968),
.B(n_845),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_855),
.A2(n_707),
.B(n_593),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_991),
.A2(n_1019),
.B(n_930),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_862),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_861),
.A2(n_945),
.A3(n_952),
.B(n_960),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_857),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1003),
.A2(n_904),
.B(n_1011),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1016),
.B(n_755),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1122),
.A2(n_1150),
.B1(n_1083),
.B2(n_1108),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1032),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1022),
.A2(n_1131),
.B(n_1118),
.C(n_1155),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1041),
.A2(n_1132),
.B1(n_1147),
.B2(n_1124),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1022),
.A2(n_1131),
.B1(n_1118),
.B2(n_1155),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1028),
.A2(n_1044),
.B(n_1058),
.C(n_1106),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1024),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1024),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1046),
.B(n_1074),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1129),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1033),
.B(n_1050),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1052),
.Y(n_1176)
);

AOI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_1044),
.A2(n_1028),
.B(n_1021),
.Y(n_1177)
);

AND2x2_ASAP7_75t_SL g1178 ( 
.A(n_1081),
.B(n_1101),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1143),
.B(n_1140),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1119),
.A2(n_1127),
.B(n_1120),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_L g1181 ( 
.A(n_1161),
.B(n_1067),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1111),
.B(n_1121),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1057),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_1130),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1033),
.B(n_1069),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1027),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1026),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1133),
.B(n_1137),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1068),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_1102),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1086),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1060),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1143),
.B(n_1123),
.Y(n_1193)
);

OR2x6_ASAP7_75t_SL g1194 ( 
.A(n_1048),
.B(n_1138),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1144),
.A2(n_1029),
.B1(n_1058),
.B2(n_1126),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1096),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1115),
.B(n_1038),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1042),
.A2(n_1142),
.B(n_1153),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1030),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1125),
.B(n_1139),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1021),
.A2(n_1073),
.B(n_1047),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1145),
.B(n_1163),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1096),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1034),
.B(n_1038),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_1112),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1151),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1141),
.B(n_1103),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1112),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1037),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1039),
.B(n_1037),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1094),
.B(n_1049),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1112),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1051),
.B(n_1064),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1078),
.B(n_1154),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1104),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_1053),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1104),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1101),
.A2(n_1059),
.B1(n_1157),
.B2(n_1110),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1100),
.B(n_1081),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1053),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1077),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1085),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1114),
.B(n_1117),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1113),
.B(n_1148),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1095),
.B(n_1158),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1148),
.B(n_1159),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1141),
.B(n_1035),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1063),
.B(n_1080),
.Y(n_1228)
);

NAND2x1_ASAP7_75t_L g1229 ( 
.A(n_1159),
.B(n_1089),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1097),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1080),
.B(n_1160),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1084),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1080),
.B(n_1099),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1134),
.B(n_1160),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1097),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1141),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1107),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1091),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1062),
.A2(n_1072),
.B(n_1106),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1088),
.B(n_1090),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_L g1241 ( 
.A(n_1098),
.B(n_1083),
.C(n_1076),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1134),
.B(n_1160),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1134),
.B(n_1160),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1075),
.B(n_1087),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1107),
.B(n_1105),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1079),
.B(n_1031),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1134),
.B(n_1031),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1105),
.B(n_1061),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1082),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1072),
.A2(n_1070),
.B(n_1079),
.Y(n_1251)
);

AO21x1_ASAP7_75t_L g1252 ( 
.A1(n_1070),
.A2(n_1071),
.B(n_1054),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1082),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1054),
.A2(n_1020),
.B(n_1066),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_L g1255 ( 
.A(n_1061),
.B(n_1045),
.Y(n_1255)
);

NAND2x1_ASAP7_75t_L g1256 ( 
.A(n_1040),
.B(n_1056),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1061),
.B(n_1162),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1061),
.B(n_1162),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1055),
.A2(n_1156),
.B1(n_1152),
.B2(n_1135),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1025),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1149),
.A2(n_1023),
.B(n_1128),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1136),
.Y(n_1262)
);

INVx3_ASAP7_75t_SL g1263 ( 
.A(n_1146),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1092),
.B(n_1109),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1092),
.B(n_1109),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1141),
.B(n_693),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1036),
.A2(n_1040),
.B(n_1025),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1129),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1032),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1111),
.B(n_1121),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1024),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1032),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1024),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1024),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1129),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1032),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1022),
.A2(n_1118),
.B(n_1155),
.C(n_1131),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1024),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1112),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1141),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1032),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1032),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1129),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1129),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1060),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1032),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1111),
.B(n_1121),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1041),
.B(n_755),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1024),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1111),
.B(n_1121),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1032),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1024),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1022),
.A2(n_1131),
.B(n_1155),
.C(n_1118),
.Y(n_1298)
);

AOI21xp33_ASAP7_75t_L g1299 ( 
.A1(n_1022),
.A2(n_1131),
.B(n_1118),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1111),
.B(n_1121),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1032),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1024),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_L g1306 ( 
.A(n_1022),
.B(n_1118),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1041),
.A2(n_844),
.B1(n_755),
.B2(n_685),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1032),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1275),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1168),
.A2(n_1219),
.B1(n_1306),
.B2(n_1178),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1186),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1225),
.B(n_1234),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1168),
.A2(n_1299),
.B1(n_1164),
.B2(n_1177),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1167),
.B(n_1307),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1256),
.A2(n_1239),
.B(n_1254),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1211),
.B(n_1204),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1291),
.A2(n_1215),
.B1(n_1193),
.B2(n_1213),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1303),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1232),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1165),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1187),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1216),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1189),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1261),
.A2(n_1267),
.B(n_1251),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1187),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1190),
.B(n_1185),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1166),
.B(n_1298),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1188),
.B(n_1304),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1276),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1201),
.B(n_1198),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1224),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1269),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1205),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1192),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1276),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1190),
.B(n_1185),
.Y(n_1336)
);

AO21x1_ASAP7_75t_L g1337 ( 
.A1(n_1278),
.A2(n_1195),
.B(n_1299),
.Y(n_1337)
);

AO21x1_ASAP7_75t_L g1338 ( 
.A1(n_1195),
.A2(n_1177),
.B(n_1218),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1226),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1180),
.A2(n_1184),
.B1(n_1179),
.B2(n_1241),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1180),
.A2(n_1241),
.B1(n_1293),
.B2(n_1202),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1287),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1282),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1295),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1182),
.A2(n_1270),
.B1(n_1301),
.B2(n_1290),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1250),
.B(n_1245),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1200),
.A2(n_1283),
.B1(n_1300),
.B2(n_1271),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1302),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1176),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1183),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1191),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1192),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1223),
.A2(n_1169),
.B(n_1228),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1248),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1268),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1206),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1294),
.A2(n_1305),
.B1(n_1253),
.B2(n_1218),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1273),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1264),
.A2(n_1265),
.B(n_1257),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1199),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1250),
.B(n_1245),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1214),
.B(n_1194),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1243),
.B(n_1249),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1208),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1199),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1209),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1238),
.B(n_1225),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1277),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1181),
.A2(n_1174),
.B1(n_1272),
.B2(n_1172),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1285),
.B(n_1308),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1289),
.B(n_1197),
.Y(n_1371)
);

BUFx2_ASAP7_75t_SL g1372 ( 
.A(n_1170),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1250),
.B(n_1246),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1274),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1279),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1286),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1292),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1240),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1171),
.B(n_1271),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1196),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1296),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1220),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1171),
.A2(n_1300),
.B1(n_1283),
.B2(n_1284),
.Y(n_1384)
);

INVx8_ASAP7_75t_L g1385 ( 
.A(n_1207),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1210),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1235),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1197),
.A2(n_1297),
.B1(n_1284),
.B2(n_1281),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1234),
.B(n_1242),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1262),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1203),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1280),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1297),
.A2(n_1240),
.B1(n_1173),
.B2(n_1175),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1244),
.A2(n_1259),
.B(n_1257),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1247),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1173),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1229),
.A2(n_1233),
.B(n_1231),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1231),
.A2(n_1258),
.B(n_1230),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1227),
.B(n_1221),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1255),
.A2(n_1263),
.B(n_1247),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1175),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1280),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1260),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1236),
.A2(n_1266),
.B1(n_1212),
.B2(n_1221),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1266),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1212),
.B(n_1266),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1288),
.A2(n_1041),
.B1(n_1188),
.B2(n_1118),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1164),
.B(n_1211),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1306),
.A2(n_879),
.B1(n_656),
.B2(n_925),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1237),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1275),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1188),
.A2(n_844),
.B1(n_1041),
.B2(n_685),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1222),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1190),
.B(n_1185),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1192),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1306),
.A2(n_879),
.B1(n_656),
.B2(n_925),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1261),
.A2(n_1025),
.B(n_1267),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1190),
.B(n_1185),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1186),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1363),
.B(n_1316),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1318),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1324),
.A2(n_1315),
.B(n_1418),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1324),
.A2(n_1315),
.B(n_1418),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1385),
.B(n_1330),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1318),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1412),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1319),
.Y(n_1428)
);

AND2x2_ASAP7_75t_SL g1429 ( 
.A(n_1313),
.B(n_1410),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1417),
.B(n_1314),
.C(n_1357),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1412),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1354),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1328),
.B(n_1386),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1322),
.Y(n_1434)
);

NAND2x1_ASAP7_75t_L g1435 ( 
.A(n_1380),
.B(n_1330),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1329),
.Y(n_1436)
);

AND2x2_ASAP7_75t_SL g1437 ( 
.A(n_1327),
.B(n_1404),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1330),
.B(n_1380),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1335),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1394),
.B(n_1396),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1399),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1409),
.B(n_1367),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1322),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1389),
.B(n_1312),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1394),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1396),
.Y(n_1446)
);

AO21x1_ASAP7_75t_SL g1447 ( 
.A1(n_1340),
.A2(n_1362),
.B(n_1312),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1389),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1413),
.A2(n_1317),
.B(n_1408),
.Y(n_1449)
);

INVx4_ASAP7_75t_SL g1450 ( 
.A(n_1380),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1398),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1359),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1365),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1360),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1353),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1353),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1353),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1409),
.B(n_1367),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1390),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1321),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1390),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1416),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1327),
.B(n_1310),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1371),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1371),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1370),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1401),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1325),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1339),
.B(n_1378),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1378),
.B(n_1404),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1366),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1380),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1395),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1309),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1338),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1388),
.B(n_1341),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1331),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1331),
.B(n_1342),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1345),
.B(n_1347),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1330),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1383),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1337),
.A2(n_1351),
.B(n_1358),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1416),
.B(n_1326),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1349),
.A2(n_1368),
.B(n_1356),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1350),
.A2(n_1387),
.B(n_1343),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1326),
.B(n_1336),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1382),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1403),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1374),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1320),
.A2(n_1344),
.B(n_1348),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1402),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1415),
.B(n_1419),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1455),
.B(n_1411),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1434),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1434),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1482),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1448),
.B(n_1411),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1361),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1438),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1457),
.B(n_1361),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1448),
.B(n_1323),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1441),
.Y(n_1503)
);

INVx2_ASAP7_75t_R g1504 ( 
.A(n_1467),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1435),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1482),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1450),
.B(n_1419),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1452),
.B(n_1346),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1464),
.B(n_1332),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1428),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1484),
.Y(n_1512)
);

AND2x4_ASAP7_75t_SL g1513 ( 
.A(n_1425),
.B(n_1416),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1484),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1442),
.B(n_1373),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1458),
.B(n_1480),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1443),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1432),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1425),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1458),
.B(n_1480),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1429),
.A2(n_1333),
.B1(n_1364),
.B2(n_1406),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1465),
.B(n_1373),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1465),
.B(n_1414),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1444),
.B(n_1372),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1451),
.B(n_1402),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1438),
.B(n_1400),
.Y(n_1528)
);

XOR2x2_ASAP7_75t_L g1529 ( 
.A(n_1430),
.B(n_1384),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1444),
.B(n_1459),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1516),
.B(n_1421),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1496),
.A2(n_1424),
.B(n_1423),
.Y(n_1532)
);

NAND4xp25_ASAP7_75t_L g1533 ( 
.A(n_1522),
.B(n_1449),
.C(n_1433),
.D(n_1460),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1525),
.B(n_1474),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1529),
.A2(n_1429),
.B(n_1476),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_L g1536 ( 
.A(n_1522),
.B(n_1429),
.C(n_1475),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1475),
.C(n_1470),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1529),
.B(n_1437),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1517),
.B(n_1422),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1516),
.B(n_1521),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1426),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1502),
.B(n_1427),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1528),
.A2(n_1437),
.B1(n_1463),
.B2(n_1393),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1529),
.A2(n_1479),
.B1(n_1488),
.B2(n_1470),
.C(n_1471),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1528),
.A2(n_1437),
.B1(n_1405),
.B2(n_1483),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1502),
.A2(n_1489),
.B(n_1379),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1431),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1497),
.B(n_1468),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_SL g1550 ( 
.A(n_1520),
.B(n_1391),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1515),
.B(n_1436),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1333),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1500),
.A2(n_1369),
.B(n_1435),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_L g1554 ( 
.A(n_1520),
.B(n_1462),
.C(n_1478),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.B(n_1440),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_1440),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1519),
.A2(n_1483),
.B(n_1466),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1493),
.B(n_1440),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1509),
.B(n_1439),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1509),
.B(n_1453),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1513),
.A2(n_1407),
.B(n_1492),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1477),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1493),
.B(n_1440),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1507),
.B(n_1364),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1508),
.B(n_1438),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1524),
.B(n_1481),
.Y(n_1566)
);

NAND3xp33_ASAP7_75t_L g1567 ( 
.A(n_1506),
.B(n_1446),
.C(n_1445),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1510),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1508),
.B(n_1523),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1508),
.B(n_1438),
.Y(n_1570)
);

OAI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1500),
.A2(n_1454),
.B1(n_1486),
.B2(n_1420),
.C(n_1311),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1523),
.B(n_1472),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1506),
.B(n_1446),
.C(n_1445),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1524),
.B(n_1469),
.Y(n_1574)
);

OAI221xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1528),
.A2(n_1425),
.B1(n_1447),
.B2(n_1487),
.C(n_1472),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1520),
.B(n_1450),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1507),
.B(n_1311),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1499),
.B(n_1501),
.Y(n_1578)
);

AOI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1518),
.A2(n_1459),
.B(n_1461),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1494),
.B(n_1469),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1494),
.B(n_1490),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1495),
.B(n_1490),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1527),
.B(n_1473),
.C(n_1491),
.Y(n_1583)
);

AND2x4_ASAP7_75t_SL g1584 ( 
.A(n_1576),
.B(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1578),
.B(n_1504),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1578),
.B(n_1504),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1549),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1569),
.B(n_1504),
.Y(n_1589)
);

AND2x4_ASAP7_75t_SL g1590 ( 
.A(n_1576),
.B(n_1528),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1569),
.B(n_1504),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1568),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1568),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1579),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1579),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1581),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1582),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1557),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1567),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1548),
.B(n_1547),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1534),
.B(n_1530),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1540),
.B(n_1530),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1532),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1532),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1539),
.B(n_1530),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1566),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1520),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1577),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1503),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1503),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1560),
.B(n_1503),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1562),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1505),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1542),
.B(n_1511),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1556),
.B(n_1498),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1585),
.Y(n_1620)
);

NOR2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1614),
.B(n_1533),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1616),
.B(n_1614),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1541),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1598),
.A2(n_1535),
.B1(n_1536),
.B2(n_1538),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1610),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1607),
.B(n_1531),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1588),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1531),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1570),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1584),
.B(n_1554),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1558),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1552),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1616),
.A2(n_1538),
.B1(n_1545),
.B2(n_1543),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1615),
.B(n_1558),
.Y(n_1637)
);

NOR2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1614),
.B(n_1616),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1592),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1602),
.B(n_1574),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1601),
.A2(n_1575),
.B(n_1553),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1563),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1570),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1601),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1606),
.B(n_1563),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1616),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1589),
.B(n_1555),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1615),
.B(n_1571),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1572),
.Y(n_1651)
);

AOI33xp33_ASAP7_75t_L g1652 ( 
.A1(n_1596),
.A2(n_1377),
.A3(n_1375),
.B1(n_1526),
.B2(n_1514),
.B3(n_1512),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1592),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1555),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1584),
.B(n_1505),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1618),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1544),
.C(n_1546),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1638),
.B(n_1608),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1620),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1633),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1608),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1608),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1644),
.B(n_1655),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1644),
.B(n_1589),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1597),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1624),
.A2(n_1537),
.B(n_1583),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1650),
.B(n_1597),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1655),
.B(n_1589),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1639),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1650),
.B(n_1617),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1655),
.B(n_1591),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1632),
.B(n_1391),
.C(n_1561),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1646),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1651),
.B(n_1617),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1632),
.B(n_1505),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1633),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1626),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1623),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1657),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1642),
.B(n_1652),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1612),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1629),
.B(n_1586),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1637),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1629),
.B(n_1586),
.Y(n_1693)
);

NAND2x1_ASAP7_75t_L g1694 ( 
.A(n_1631),
.B(n_1593),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1656),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1587),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1635),
.B(n_1613),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1635),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1649),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1641),
.B(n_1611),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1660),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1660),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1661),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1669),
.B(n_1634),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1661),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1665),
.B(n_1648),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1686),
.A2(n_1636),
.B1(n_1631),
.B2(n_1520),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1671),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1700),
.B(n_1625),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1665),
.B(n_1631),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1686),
.B(n_1625),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1694),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1672),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1700),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1694),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1700),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1687),
.A2(n_1584),
.B1(n_1590),
.B2(n_1500),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1698),
.Y(n_1721)
);

AOI222xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1698),
.A2(n_1668),
.B1(n_1684),
.B2(n_1685),
.C1(n_1683),
.C2(n_1682),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1669),
.B(n_1658),
.Y(n_1723)
);

AO21x1_ASAP7_75t_L g1724 ( 
.A1(n_1687),
.A2(n_1594),
.B(n_1595),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1681),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1663),
.B(n_1654),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1689),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1689),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1663),
.B(n_1587),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1659),
.B(n_1590),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1664),
.B(n_1587),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1699),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1677),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1666),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1677),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1682),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1659),
.B(n_1590),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1673),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1727),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1713),
.B(n_1673),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1711),
.B(n_1697),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1664),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1727),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1702),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1702),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1703),
.Y(n_1746)
);

OAI31xp33_ASAP7_75t_L g1747 ( 
.A1(n_1728),
.A2(n_1688),
.A3(n_1697),
.B(n_1685),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1711),
.B(n_1668),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1704),
.Y(n_1751)
);

AOI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1719),
.A2(n_1688),
.B(n_1667),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1722),
.A2(n_1684),
.B1(n_1667),
.B2(n_1676),
.C(n_1692),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1670),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1717),
.A2(n_1676),
.B(n_1683),
.C(n_1699),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1717),
.B(n_1381),
.Y(n_1756)
);

AOI33xp33_ASAP7_75t_L g1757 ( 
.A1(n_1720),
.A2(n_1699),
.A3(n_1662),
.B1(n_1695),
.B2(n_1678),
.B3(n_1675),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1679),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1708),
.A2(n_1717),
.B(n_1707),
.C(n_1714),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_L g1760 ( 
.A(n_1714),
.B(n_1381),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1706),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1724),
.A2(n_1630),
.B(n_1662),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1706),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1749),
.B(n_1709),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1744),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1740),
.B(n_1709),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1740),
.B(n_1710),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1754),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1745),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1742),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1746),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1739),
.B(n_1714),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1738),
.B(n_1723),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1705),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1742),
.B(n_1707),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1741),
.B(n_1734),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1747),
.B(n_1734),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1748),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1743),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1730),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1750),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1782),
.A2(n_1760),
.B(n_1755),
.Y(n_1784)
);

NAND2x1_ASAP7_75t_L g1785 ( 
.A(n_1773),
.B(n_1714),
.Y(n_1785)
);

OAI21xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1764),
.A2(n_1757),
.B(n_1753),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1764),
.A2(n_1759),
.B(n_1752),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1779),
.A2(n_1759),
.B(n_1724),
.C(n_1762),
.Y(n_1788)
);

AOI32xp33_ASAP7_75t_L g1789 ( 
.A1(n_1777),
.A2(n_1743),
.A3(n_1725),
.B1(n_1718),
.B2(n_1751),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1770),
.A2(n_1730),
.B1(n_1737),
.B2(n_1718),
.Y(n_1790)
);

NOR4xp25_ASAP7_75t_L g1791 ( 
.A(n_1781),
.B(n_1761),
.C(n_1763),
.D(n_1757),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_SL g1792 ( 
.A(n_1772),
.B(n_1716),
.C(n_1715),
.Y(n_1792)
);

OAI211xp5_ASAP7_75t_L g1793 ( 
.A1(n_1766),
.A2(n_1715),
.B(n_1733),
.C(n_1716),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1776),
.Y(n_1794)
);

AOI21xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1775),
.A2(n_1735),
.B(n_1733),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1775),
.B(n_1730),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_L g1797 ( 
.A1(n_1778),
.A2(n_1732),
.B(n_1735),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1786),
.B(n_1776),
.C(n_1767),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1792),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1785),
.Y(n_1800)
);

OAI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1791),
.A2(n_1768),
.B(n_1774),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1788),
.B(n_1767),
.C(n_1766),
.Y(n_1802)
);

OAI211xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1787),
.A2(n_1765),
.B(n_1771),
.C(n_1769),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1793),
.Y(n_1804)
);

NOR3xp33_ASAP7_75t_L g1805 ( 
.A(n_1784),
.B(n_1783),
.C(n_1780),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1794),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1789),
.B(n_1730),
.Y(n_1807)
);

NOR4xp25_ASAP7_75t_L g1808 ( 
.A(n_1797),
.B(n_1796),
.C(n_1795),
.D(n_1732),
.Y(n_1808)
);

NAND4xp75_ASAP7_75t_L g1809 ( 
.A(n_1790),
.B(n_1732),
.C(n_1736),
.D(n_1729),
.Y(n_1809)
);

NAND4xp25_ASAP7_75t_L g1810 ( 
.A(n_1798),
.B(n_1736),
.C(n_1737),
.D(n_1420),
.Y(n_1810)
);

NOR4xp25_ASAP7_75t_L g1811 ( 
.A(n_1801),
.B(n_1662),
.C(n_1392),
.D(n_1729),
.Y(n_1811)
);

NAND4xp25_ASAP7_75t_L g1812 ( 
.A(n_1802),
.B(n_1737),
.C(n_1376),
.D(n_1731),
.Y(n_1812)
);

NOR4xp75_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1809),
.C(n_1808),
.D(n_1805),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1803),
.B(n_1406),
.C(n_1392),
.Y(n_1814)
);

AOI322xp5_ASAP7_75t_L g1815 ( 
.A1(n_1799),
.A2(n_1737),
.A3(n_1731),
.B1(n_1726),
.B2(n_1695),
.C1(n_1670),
.C2(n_1674),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1810),
.B(n_1800),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1813),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1812),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1814),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1811),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1810),
.Y(n_1822)
);

NAND4xp75_ASAP7_75t_L g1823 ( 
.A(n_1816),
.B(n_1804),
.C(n_1806),
.D(n_1803),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1817),
.Y(n_1824)
);

NAND4xp25_ASAP7_75t_L g1825 ( 
.A(n_1821),
.B(n_1376),
.C(n_1726),
.D(n_1564),
.Y(n_1825)
);

NAND2x1_ASAP7_75t_L g1826 ( 
.A(n_1819),
.B(n_1674),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1822),
.B(n_1818),
.Y(n_1827)
);

XNOR2xp5_ASAP7_75t_L g1828 ( 
.A(n_1817),
.B(n_1397),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1824),
.Y(n_1829)
);

XNOR2xp5_ASAP7_75t_L g1830 ( 
.A(n_1828),
.B(n_1820),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1826),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1831),
.Y(n_1832)
);

OAI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1829),
.B1(n_1830),
.B2(n_1827),
.C1(n_1823),
.C2(n_1825),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1695),
.B1(n_1678),
.B2(n_1675),
.C(n_1666),
.Y(n_1834)
);

AOI221x1_ASAP7_75t_L g1835 ( 
.A1(n_1833),
.A2(n_1690),
.B1(n_1691),
.B2(n_1693),
.C(n_1604),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1701),
.B(n_1690),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1834),
.A2(n_1693),
.B(n_1691),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1701),
.B(n_1696),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1696),
.B(n_1680),
.Y(n_1839)
);

NAND4xp25_ASAP7_75t_L g1840 ( 
.A(n_1838),
.B(n_1355),
.C(n_1462),
.D(n_1680),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1840),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1839),
.B1(n_1355),
.B2(n_1605),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1416),
.B(n_1334),
.C(n_1352),
.Y(n_1843)
);


endmodule