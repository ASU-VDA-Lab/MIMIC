module real_jpeg_30858_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_0),
.Y(n_392)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_0),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_1),
.A2(n_75),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_1),
.A2(n_75),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_1),
.A2(n_75),
.B1(n_395),
.B2(n_398),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_109),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_2),
.A2(n_109),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_2),
.A2(n_109),
.B1(n_335),
.B2(n_338),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_3),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_4),
.A2(n_77),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_4),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_4),
.A2(n_353),
.B1(n_455),
.B2(n_459),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_4),
.A2(n_353),
.B1(n_549),
.B2(n_551),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_4),
.A2(n_353),
.B1(n_617),
.B2(n_621),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_6),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_124),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_124),
.B1(n_223),
.B2(n_226),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_6),
.A2(n_124),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_7),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_7),
.A2(n_276),
.B1(n_381),
.B2(n_385),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_7),
.A2(n_223),
.B1(n_276),
.B2(n_503),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_7),
.A2(n_276),
.B1(n_595),
.B2(n_596),
.Y(n_594)
);

OAI22x1_ASAP7_75t_SL g259 ( 
.A1(n_8),
.A2(n_107),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_8),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_8),
.A2(n_260),
.B1(n_360),
.B2(n_362),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_8),
.A2(n_260),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_8),
.A2(n_260),
.B1(n_530),
.B2(n_535),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_9),
.A2(n_60),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_9),
.A2(n_60),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_11),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_12),
.Y(n_238)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_12),
.Y(n_534)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_13),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_14),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_14),
.A2(n_189),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_14),
.A2(n_189),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_14),
.A2(n_189),
.B1(n_474),
.B2(n_477),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_20),
.B(n_657),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_15),
.B(n_658),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_16),
.B(n_93),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_16),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_16),
.B(n_113),
.Y(n_481)
);

OAI32xp33_ASAP7_75t_L g507 ( 
.A1(n_16),
.A2(n_508),
.A3(n_511),
.B1(n_513),
.B2(n_520),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_16),
.A2(n_450),
.B1(n_543),
.B2(n_546),
.Y(n_542)
);

OAI21xp33_ASAP7_75t_L g632 ( 
.A1(n_16),
.A2(n_298),
.B(n_598),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_17),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_18),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_18),
.Y(n_128)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_203),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_202),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_177),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_24),
.B(n_177),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_165),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_67),
.C(n_114),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_26),
.A2(n_27),
.B1(n_114),
.B2(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_27),
.B(n_182),
.C(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_27),
.B(n_193),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_44),
.B(n_57),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_28),
.A2(n_44),
.B1(n_57),
.B2(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_28),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_28),
.A2(n_44),
.B1(n_438),
.B2(n_444),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_28),
.B(n_438),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_46),
.Y(n_45)
);

OAI22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_32),
.Y(n_242)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_32),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_47),
.B1(n_50),
.B2(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_37),
.Y(n_399)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_37),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_38),
.Y(n_245)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_38),
.Y(n_397)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_38),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_38),
.Y(n_537)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_44),
.B(n_587),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_44),
.B(n_438),
.Y(n_603)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_45),
.A2(n_222),
.B1(n_248),
.B2(n_255),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_45),
.A2(n_248),
.B1(n_255),
.B2(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_45),
.A2(n_255),
.B1(n_303),
.B2(n_345),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g501 ( 
.A1(n_45),
.A2(n_502),
.B(n_505),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_45),
.A2(n_255),
.B1(n_502),
.B2(n_548),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_47),
.Y(n_249)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_49),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_49),
.Y(n_512)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_55),
.Y(n_441)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_56),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_56),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_59),
.Y(n_347)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_59),
.Y(n_443)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_66),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_67),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_80),
.B1(n_105),
.B2(n_112),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_69),
.A2(n_81),
.B1(n_113),
.B2(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_74),
.Y(n_265)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_79),
.Y(n_449)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_113),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_83),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_83),
.B(n_275),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g351 ( 
.A1(n_83),
.A2(n_113),
.B1(n_275),
.B2(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_83),
.B(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_85),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_86),
.Y(n_384)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_88),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_88),
.Y(n_419)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_91),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_99),
.B2(n_103),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_100),
.Y(n_356)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g190 ( 
.A(n_108),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_113),
.B(n_184),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_113),
.B(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_113),
.B(n_352),
.Y(n_376)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22x1_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_129),
.B1(n_154),
.B2(n_161),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_116),
.A2(n_131),
.B1(n_161),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_122),
.Y(n_287)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_122),
.Y(n_361)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_123),
.Y(n_545)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_127),
.Y(n_546)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_128),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_154),
.B(n_161),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_129),
.A2(n_161),
.B1(n_194),
.B2(n_216),
.Y(n_215)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_129),
.A2(n_161),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22x1_ASAP7_75t_L g357 ( 
.A1(n_130),
.A2(n_162),
.B1(n_358),
.B2(n_363),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_130),
.A2(n_380),
.B(n_387),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_130),
.A2(n_387),
.B(n_542),
.Y(n_541)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_131),
.A2(n_163),
.B1(n_216),
.B2(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_131),
.B(n_359),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_139),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_137),
.B1(n_139),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_136),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_145),
.B1(n_148),
.B2(n_153),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_143),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_144),
.Y(n_463)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_162),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_162),
.B(n_450),
.Y(n_601)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_163),
.B(n_359),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_175),
.B2(n_176),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_174),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_191),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_212),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_183),
.A2(n_212),
.B(n_213),
.C(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_183),
.Y(n_318)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_319),
.B(n_652),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_267),
.Y(n_205)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_206),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_207),
.B(n_210),
.Y(n_656)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_229),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_211),
.A2(n_213),
.B(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_212),
.A2(n_214),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_215),
.B(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx4f_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_229),
.B(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_246),
.B(n_256),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_230),
.A2(n_231),
.B1(n_257),
.B2(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_230),
.A2(n_231),
.B1(n_247),
.B2(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_247),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_235),
.B(n_241),
.Y(n_231)
);

BUFx2_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_233),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_234),
.Y(n_630)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

AO22x1_ASAP7_75t_SL g390 ( 
.A1(n_235),
.A2(n_334),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_235),
.B(n_529),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_235),
.A2(n_391),
.B1(n_615),
.B2(n_623),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_238),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_238),
.Y(n_479)
);

INVx4_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g527 ( 
.A(n_240),
.Y(n_527)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_247),
.Y(n_365)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_253),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_254),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_254),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_255),
.A2(n_548),
.B(n_603),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_255),
.B(n_450),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_257),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_258),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_314),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_268),
.B(n_314),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.C(n_310),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_270),
.B(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2x2_ASAP7_75t_L g366 ( 
.A(n_272),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_283),
.C(n_290),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_273),
.A2(n_284),
.B1(n_285),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_282),
.B(n_446),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_292),
.B(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_298),
.B1(n_333),
.B2(n_341),
.Y(n_332)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_294),
.Y(n_577)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_298),
.A2(n_341),
.B1(n_394),
.B2(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_298),
.A2(n_594),
.B(n_598),
.Y(n_593)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_300),
.Y(n_599)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_309),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2x1_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_491),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_425),
.B(n_487),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_322),
.B(n_649),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_366),
.B(n_368),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_323),
.B(n_366),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_323),
.B(n_366),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.C(n_364),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_325),
.A2(n_326),
.B1(n_364),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_351),
.C(n_357),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_331),
.B(n_424),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_344),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_332),
.B(n_344),
.Y(n_434)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_345),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_351),
.B(n_357),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_364),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_369),
.B(n_372),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_420),
.C(n_422),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.C(n_388),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_374),
.A2(n_375),
.B1(n_378),
.B2(n_379),
.Y(n_432)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_384),
.Y(n_386)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_388),
.A2(n_389),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_400),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_390),
.A2(n_400),
.B1(n_401),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_397),
.Y(n_640)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AOI32xp33_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_405),
.A3(n_409),
.B1(n_413),
.B2(n_414),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_413),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_423),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.C(n_464),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_SL g649 ( 
.A1(n_427),
.A2(n_650),
.B(n_651),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_429),
.Y(n_650)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.C(n_435),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_433),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_445),
.C(n_452),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_452),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_467),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_450),
.B(n_451),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_450),
.B(n_521),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_450),
.B(n_511),
.Y(n_575)
);

OAI21xp33_ASAP7_75t_SL g587 ( 
.A1(n_450),
.A2(n_575),
.B(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_450),
.B(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_454),
.Y(n_483)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_485),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_465),
.B(n_485),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_468),
.C(n_470),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_466),
.B(n_558),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_468),
.A2(n_470),
.B1(n_471),
.B2(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_468),
.Y(n_559)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_480),
.C(n_482),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_480),
.B1(n_481),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_473),
.A2(n_525),
.B(n_528),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2x2_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B(n_490),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_648),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_560),
.B(n_646),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_553),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_538),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_495),
.B(n_538),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_496),
.B(n_500),
.C(n_556),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_506),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_505),
.B(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_524),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_507),
.B(n_524),
.Y(n_539)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx2_ASAP7_75t_SL g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx3_ASAP7_75t_SL g521 ( 
.A(n_522),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_526),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_528),
.A2(n_616),
.B(n_629),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_529),
.B(n_599),
.Y(n_598)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_531),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx6_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

MAJx2_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.C(n_547),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_539),
.B(n_610),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_541),
.B(n_547),
.Y(n_610)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_557),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_555),
.B(n_647),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_557),
.Y(n_647)
);

AOI211x1_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_611),
.B(n_643),
.C(n_645),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_562),
.A2(n_604),
.B(n_605),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_562),
.B(n_612),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_592),
.Y(n_562)
);

NOR2x1_ASAP7_75t_SL g604 ( 
.A(n_563),
.B(n_592),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_585),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_564),
.B(n_585),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_574),
.B1(n_576),
.B2(n_578),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_570),
.Y(n_565)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_571),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_573),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_582),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

XNOR2x1_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_600),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_607),
.C(n_608),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_594),
.Y(n_623)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_601),
.B(n_602),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_601),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_602),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_609),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_606),
.B(n_609),
.Y(n_644)
);

AOI21xp33_ASAP7_75t_L g612 ( 
.A1(n_613),
.A2(n_625),
.B(n_642),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_614),
.B(n_624),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_614),
.B(n_624),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

BUFx2_ASAP7_75t_SL g619 ( 
.A(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_626),
.A2(n_631),
.B(n_641),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_627),
.B(n_628),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_627),
.B(n_628),
.Y(n_641)
);

INVx8_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_634),
.B(n_639),
.Y(n_633)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_653),
.A2(n_654),
.B(n_655),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_656),
.Y(n_655)
);


endmodule