module fake_jpeg_32061_n_36 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_36);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_5),
.A2(n_4),
.B1(n_1),
.B2(n_12),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_17),
.C(n_13),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_2),
.C(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_22),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_17),
.B(n_13),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.C(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_31),
.B(n_9),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_11),
.C(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_10),
.Y(n_36)
);


endmodule