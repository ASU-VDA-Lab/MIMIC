module fake_jpeg_9415_n_45 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_21),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_5),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_2),
.B(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_39),
.B1(n_32),
.B2(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_44)
);

OAI221xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.C(n_15),
.Y(n_45)
);


endmodule