module fake_jpeg_6196_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_31),
.Y(n_48)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_35),
.B1(n_39),
.B2(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_26),
.C(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_15),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_28),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_16),
.B1(n_44),
.B2(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_3),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_19),
.B1(n_17),
.B2(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_43),
.B1(n_17),
.B2(n_12),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_38),
.B2(n_22),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_60),
.C(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_4),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_13),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_86),
.B1(n_63),
.B2(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_60),
.C(n_50),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_71),
.C(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_102),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_90),
.C(n_86),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_72),
.C(n_78),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_93),
.B(n_94),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_63),
.B1(n_72),
.B2(n_59),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_79),
.C(n_82),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_101),
.B1(n_100),
.B2(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_23),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_113),
.A2(n_114),
.B(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_23),
.C(n_6),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_23),
.B(n_7),
.C(n_5),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_117),
.B(n_118),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_122),
.B(n_55),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_7),
.Y(n_125)
);


endmodule