module fake_jpeg_31120_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_10),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_1),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_49),
.C(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_83),
.B1(n_59),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_57),
.B1(n_50),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_88),
.B1(n_64),
.B2(n_52),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_50),
.B1(n_67),
.B2(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_108),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_106),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_29),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_58),
.B1(n_53),
.B2(n_51),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_2),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_116),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_42),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_4),
.C(n_6),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_48),
.B1(n_28),
.B2(n_30),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_121),
.B1(n_127),
.B2(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_27),
.B1(n_46),
.B2(n_45),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_7),
.B(n_8),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_8),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_38),
.B1(n_19),
.B2(n_20),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_136),
.C(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_12),
.B1(n_23),
.B2(n_24),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_141),
.Y(n_148)
);

AND2x4_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_32),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_144),
.C(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_119),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_154),
.C(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_121),
.C(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_135),
.B1(n_144),
.B2(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_134),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_139),
.B1(n_129),
.B2(n_131),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_155),
.C(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_160),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_149),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_147),
.Y(n_167)
);


endmodule