module fake_jpeg_29057_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_SL g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_22),
.B1(n_26),
.B2(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_3),
.B1(n_9),
.B2(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_17),
.C(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.C(n_28),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_37),
.B1(n_31),
.B2(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_19),
.B1(n_25),
.B2(n_20),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_36),
.C(n_28),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_24),
.A3(n_20),
.B1(n_10),
.B2(n_25),
.C1(n_16),
.C2(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_24),
.C(n_52),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_24),
.C(n_10),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_54),
.B(n_10),
.C(n_16),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_16),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);


endmodule