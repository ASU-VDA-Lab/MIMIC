module fake_aes_7802_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_9), .B(n_2), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_7), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_3), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
NOR2xp67_ASAP7_75t_SL g20 ( .A(n_14), .B(n_10), .Y(n_20) );
AOI221x1_ASAP7_75t_L g21 ( .A1(n_14), .A2(n_8), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_15), .B(n_7), .Y(n_22) );
NAND2xp33_ASAP7_75t_SL g23 ( .A(n_20), .B(n_13), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_19), .B(n_16), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_22), .Y(n_26) );
INVxp33_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_24), .B1(n_20), .B2(n_16), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_23), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_26), .B1(n_28), .B2(n_12), .C(n_21), .Y(n_31) );
OAI31xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_12), .A3(n_0), .B(n_6), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_6), .Y(n_33) );
BUFx12f_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_31), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_33), .Y(n_36) );
AOI22xp5_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_33), .B1(n_35), .B2(n_34), .Y(n_37) );
endmodule