module fake_ariane_678_n_1892 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1892);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1892;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g171 ( 
.A(n_58),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_20),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_98),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_54),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_7),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_37),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_75),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_71),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_70),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_87),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_62),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_64),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_74),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_43),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_58),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_55),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_40),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_14),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_41),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_81),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_145),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_103),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_48),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_146),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_47),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_139),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_61),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_80),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_129),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_97),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_17),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_151),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_104),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_50),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_23),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_60),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_46),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_36),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_163),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_121),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_25),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_0),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_149),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_29),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_53),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_59),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_162),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_26),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_60),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_94),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_142),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_22),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_82),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_120),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_8),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_29),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_113),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_44),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_110),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_31),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_168),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_65),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_65),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_16),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_26),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_116),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_28),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_52),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_93),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_56),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_11),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_122),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_35),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_144),
.Y(n_308)
);

BUFx8_ASAP7_75t_SL g309 ( 
.A(n_138),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_91),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_132),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_128),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_92),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_28),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_83),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_88),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_3),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_150),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_12),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_153),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_127),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_78),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_156),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_67),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_133),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_68),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_66),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_84),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_15),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_119),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_32),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_17),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_137),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_38),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_135),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_52),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_4),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_173),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_319),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_254),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_309),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_180),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_240),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_311),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_262),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_262),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_226),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_180),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_185),
.B(n_1),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_208),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_185),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_174),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_248),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_248),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_179),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_266),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_319),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_298),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_331),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_266),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_187),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_187),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_195),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_198),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_198),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_171),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_176),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_298),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_248),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_183),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_200),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_200),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_212),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_186),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_340),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_248),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_207),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_301),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_220),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_231),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_190),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_231),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_192),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_232),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_194),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_232),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_260),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_202),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_178),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_235),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_205),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_235),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_236),
.B(n_1),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_301),
.B(n_108),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_206),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_238),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_216),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_216),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_225),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_243),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_238),
.B(n_2),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_260),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_300),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_244),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_210),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_211),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_215),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_244),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_251),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_251),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_196),
.B(n_3),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_340),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_341),
.B(n_300),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_228),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_358),
.A2(n_283),
.B1(n_280),
.B2(n_318),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_345),
.A2(n_263),
.B(n_259),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_341),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_359),
.A2(n_263),
.B(n_259),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_353),
.B(n_305),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_346),
.B(n_305),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_274),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_349),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_357),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_369),
.B(n_370),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_371),
.B(n_274),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

BUFx8_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_372),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_373),
.B(n_178),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_373),
.B(n_216),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_380),
.B(n_181),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_382),
.A2(n_230),
.B(n_199),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_383),
.B(n_181),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_383),
.B(n_277),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_277),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_306),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_395),
.B(n_306),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_397),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_403),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_410),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_478),
.B(n_366),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_436),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_462),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_478),
.B(n_366),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_429),
.B(n_377),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_410),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_379),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_R g517 ( 
.A(n_433),
.B(n_350),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_451),
.B(n_347),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_469),
.B(n_342),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_462),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_469),
.B(n_310),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_463),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_462),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_445),
.B(n_405),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_426),
.B(n_347),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_427),
.A2(n_389),
.B1(n_377),
.B2(n_423),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_431),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_427),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_437),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_429),
.B(n_389),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_462),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_463),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_451),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_473),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_469),
.B(n_376),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_423),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_482),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_433),
.B(n_356),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_SL g549 ( 
.A(n_439),
.B(n_223),
.C(n_219),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_482),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_451),
.B(n_445),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_445),
.B(n_384),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_476),
.B(n_406),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_426),
.A2(n_348),
.B1(n_404),
.B2(n_355),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_458),
.B(n_399),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_473),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_482),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_426),
.A2(n_413),
.B1(n_329),
.B2(n_270),
.Y(n_560)
);

OAI21xp33_ASAP7_75t_L g561 ( 
.A1(n_465),
.A2(n_416),
.B(n_408),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_445),
.B(n_347),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_433),
.B(n_356),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_477),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_496),
.B(n_408),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_473),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

INVx8_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_469),
.B(n_392),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_476),
.B(n_416),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_483),
.A2(n_312),
.B(n_310),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_473),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_496),
.B(n_420),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_473),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_480),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_496),
.B(n_420),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_473),
.B(n_394),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_426),
.A2(n_265),
.B1(n_291),
.B2(n_295),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_480),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_480),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_496),
.B(n_396),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_453),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_458),
.B(n_402),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_498),
.B(n_407),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_495),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_426),
.B(n_417),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_495),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_452),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_455),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_498),
.B(n_422),
.C(n_421),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_476),
.B(n_481),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_455),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_498),
.B(n_418),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_495),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_498),
.B(n_421),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_477),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_465),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_452),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_477),
.B(n_335),
.C(n_250),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_476),
.B(n_365),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_452),
.B(n_419),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_441),
.B(n_344),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_L g616 ( 
.A(n_441),
.B(n_221),
.C(n_201),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_457),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_476),
.B(n_422),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_467),
.B(n_367),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_467),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_464),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_457),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_468),
.B(n_386),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_468),
.B(n_361),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_468),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_472),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_450),
.B(n_400),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_472),
.B(n_361),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_464),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_472),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_474),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_450),
.B(n_234),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_457),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_481),
.B(n_234),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_474),
.B(n_362),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_481),
.B(n_381),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_457),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_481),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_481),
.B(n_343),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_471),
.A2(n_362),
.B1(n_414),
.B2(n_398),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_464),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_464),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_466),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_466),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_481),
.A2(n_201),
.B1(n_284),
.B2(n_288),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_485),
.B(n_234),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_474),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_485),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_475),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_475),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_485),
.B(n_234),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_600),
.B(n_475),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_591),
.A2(n_556),
.B1(n_600),
.B2(n_500),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_551),
.A2(n_486),
.B(n_471),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_639),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_514),
.B(n_479),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_568),
.Y(n_658)
);

INVx8_ASAP7_75t_L g659 ( 
.A(n_568),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_639),
.B(n_479),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_510),
.B(n_479),
.Y(n_661)
);

BUFx4_ASAP7_75t_L g662 ( 
.A(n_530),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_639),
.B(n_487),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_613),
.B(n_487),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_548),
.B(n_490),
.C(n_487),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_650),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_535),
.B(n_490),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_490),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_650),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_613),
.B(n_491),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_507),
.B(n_491),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_613),
.B(n_491),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_608),
.B(n_519),
.C(n_609),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_613),
.B(n_492),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_609),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_639),
.B(n_492),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_546),
.A2(n_492),
.B1(n_499),
.B2(n_494),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_521),
.A2(n_446),
.B1(n_443),
.B2(n_485),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_649),
.B(n_499),
.Y(n_679)
);

OAI221xp5_ASAP7_75t_L g680 ( 
.A1(n_555),
.A2(n_264),
.B1(n_221),
.B2(n_222),
.C(n_229),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_649),
.B(n_499),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_519),
.B(n_485),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_649),
.B(n_533),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_564),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_622),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_622),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_428),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_629),
.B(n_485),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_619),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_630),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_636),
.B(n_466),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_562),
.B(n_466),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_630),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_513),
.B(n_470),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_630),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_649),
.B(n_470),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_532),
.B(n_470),
.Y(n_697)
);

OA22x2_ASAP7_75t_L g698 ( 
.A1(n_560),
.A2(n_439),
.B1(n_414),
.B2(n_398),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_532),
.B(n_534),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_534),
.B(n_620),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_545),
.B(n_486),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_533),
.B(n_470),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_533),
.B(n_484),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_600),
.B(n_484),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_569),
.B(n_489),
.Y(n_705)
);

OAI221xp5_ASAP7_75t_L g706 ( 
.A1(n_555),
.A2(n_288),
.B1(n_229),
.B2(n_233),
.C(n_253),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_594),
.B(n_489),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_572),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_596),
.B(n_493),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_624),
.B(n_587),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_572),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_607),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_596),
.B(n_484),
.Y(n_713)
);

NAND3x1_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_585),
.C(n_611),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_568),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_619),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_528),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_610),
.B(n_484),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_646),
.A2(n_222),
.B1(n_294),
.B2(n_297),
.C(n_233),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_581),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_488),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_600),
.B(n_488),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_542),
.B(n_488),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_600),
.B(n_488),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_600),
.A2(n_546),
.B1(n_525),
.B2(n_527),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_581),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_621),
.Y(n_727)
);

HB1xp67_ASAP7_75t_SL g728 ( 
.A(n_522),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_517),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_626),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_600),
.B(n_497),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_522),
.B(n_493),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_526),
.B(n_497),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_541),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_548),
.B(n_563),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_563),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_521),
.A2(n_546),
.B1(n_561),
.B2(n_443),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_554),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_628),
.B(n_439),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_626),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_627),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_542),
.B(n_497),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_644),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_558),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_614),
.B(n_494),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_497),
.C(n_239),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_627),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_541),
.B(n_428),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_589),
.B(n_592),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_568),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_554),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_637),
.B(n_428),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_558),
.B(n_443),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_521),
.A2(n_443),
.B1(n_446),
.B2(n_428),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_542),
.B(n_483),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_631),
.Y(n_757)
);

BUFx6f_ASAP7_75t_SL g758 ( 
.A(n_526),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_637),
.B(n_456),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_640),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_631),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_521),
.A2(n_443),
.B1(n_446),
.B2(n_456),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_526),
.B(n_456),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_573),
.B(n_483),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_644),
.Y(n_765)
);

BUFx8_ASAP7_75t_L g766 ( 
.A(n_640),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_546),
.A2(n_456),
.B1(n_312),
.B2(n_313),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_603),
.B(n_224),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_632),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_584),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_635),
.B(n_242),
.Y(n_772)
);

AO22x2_ASAP7_75t_L g773 ( 
.A1(n_583),
.A2(n_253),
.B1(n_261),
.B2(n_264),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_584),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_632),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_526),
.B(n_443),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_518),
.B(n_443),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_546),
.A2(n_313),
.B1(n_325),
.B2(n_336),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_590),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_641),
.B(n_273),
.C(n_261),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_573),
.B(n_483),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_573),
.B(n_325),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_571),
.B(n_446),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_571),
.B(n_446),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_566),
.B(n_364),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_590),
.Y(n_788)
);

INVx8_ASAP7_75t_L g789 ( 
.A(n_554),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_571),
.B(n_336),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_648),
.B(n_199),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_554),
.A2(n_570),
.B1(n_618),
.B2(n_648),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_521),
.B(n_245),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_642),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_579),
.B(n_275),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_579),
.B(n_275),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_570),
.Y(n_797)
);

NOR2xp67_ASAP7_75t_L g798 ( 
.A(n_566),
.B(n_415),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_579),
.B(n_230),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_521),
.A2(n_247),
.B1(n_255),
.B2(n_249),
.Y(n_800)
);

INVx8_ASAP7_75t_L g801 ( 
.A(n_570),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_597),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_651),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_651),
.A2(n_446),
.B(n_425),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_570),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_588),
.B(n_593),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_577),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_647),
.B(n_252),
.Y(n_808)
);

BUFx6f_ASAP7_75t_SL g809 ( 
.A(n_521),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_585),
.B(n_415),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_586),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_595),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_588),
.B(n_446),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_616),
.B(n_388),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_570),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_618),
.A2(n_257),
.B1(n_256),
.B2(n_267),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_540),
.B(n_268),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_618),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_595),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_618),
.B(n_281),
.C(n_271),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_675),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_707),
.B(n_618),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_657),
.A2(n_606),
.B(n_593),
.Y(n_823)
);

OAI321xp33_ASAP7_75t_L g824 ( 
.A1(n_680),
.A2(n_304),
.A3(n_273),
.B1(n_276),
.B2(n_307),
.C(n_303),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_707),
.A2(n_576),
.B(n_565),
.Y(n_825)
);

NOR2x1_ASAP7_75t_L g826 ( 
.A(n_684),
.B(n_543),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_654),
.A2(n_593),
.B1(n_601),
.B2(n_604),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_792),
.A2(n_601),
.B1(n_588),
.B2(n_604),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_601),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_694),
.A2(n_756),
.B(n_764),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_706),
.A2(n_580),
.B(n_605),
.C(n_606),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_756),
.A2(n_604),
.B(n_511),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_659),
.B(n_575),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_764),
.A2(n_511),
.B(n_506),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_709),
.B(n_575),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_785),
.A2(n_813),
.B(n_786),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_745),
.B(n_652),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_783),
.A2(n_516),
.B(n_506),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_783),
.A2(n_520),
.B(n_516),
.Y(n_839)
);

BUFx12f_ASAP7_75t_L g840 ( 
.A(n_734),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_745),
.B(n_501),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_689),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_701),
.A2(n_574),
.B(n_598),
.C(n_561),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_725),
.A2(n_598),
.B(n_502),
.C(n_503),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_716),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_701),
.B(n_501),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_735),
.A2(n_285),
.B(n_282),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_655),
.A2(n_523),
.B(n_520),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_685),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_714),
.A2(n_578),
.B1(n_633),
.B2(n_508),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_727),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_659),
.Y(n_852)
);

OAI22x1_ASAP7_75t_L g853 ( 
.A1(n_739),
.A2(n_411),
.B1(n_412),
.B2(n_549),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_778),
.A2(n_537),
.B(n_523),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_732),
.A2(n_505),
.B1(n_536),
.B2(n_531),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_789),
.B(n_502),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_705),
.B(n_503),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_760),
.B(n_284),
.C(n_276),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_738),
.A2(n_512),
.B1(n_536),
.B2(n_531),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_685),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_686),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_688),
.A2(n_512),
.B(n_505),
.C(n_508),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_705),
.B(n_557),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_668),
.B(n_557),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_712),
.B(n_642),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_806),
.A2(n_538),
.B(n_537),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_692),
.A2(n_539),
.B(n_538),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_717),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_729),
.B(n_509),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_749),
.B(n_509),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_661),
.A2(n_645),
.B(n_643),
.C(n_509),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_665),
.B(n_515),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_704),
.A2(n_547),
.B(n_539),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_668),
.B(n_643),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_730),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_687),
.B(n_279),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_777),
.B(n_645),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_653),
.B(n_737),
.Y(n_878)
);

OAI22x1_ASAP7_75t_L g879 ( 
.A1(n_810),
.A2(n_315),
.B1(n_287),
.B2(n_302),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_671),
.B(n_515),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_659),
.B(n_540),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_550),
.B(n_547),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_702),
.A2(n_550),
.B(n_559),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_736),
.Y(n_884)
);

BUFx4f_ASAP7_75t_L g885 ( 
.A(n_767),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_703),
.A2(n_567),
.B(n_559),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_703),
.A2(n_567),
.B(n_524),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_738),
.A2(n_515),
.B1(n_524),
.B2(n_553),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_671),
.B(n_524),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_723),
.A2(n_553),
.B(n_544),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_661),
.B(n_553),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_667),
.B(n_597),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_667),
.A2(n_294),
.B(n_307),
.C(n_304),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_686),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_723),
.A2(n_544),
.B(n_540),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_682),
.B(n_599),
.Y(n_896)
);

CKINVDCx10_ASAP7_75t_R g897 ( 
.A(n_662),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_746),
.B(n_599),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_818),
.A2(n_750),
.B1(n_758),
.B2(n_805),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_795),
.A2(n_638),
.B(n_634),
.C(n_623),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_763),
.B(n_602),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_742),
.A2(n_638),
.B(n_612),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_700),
.A2(n_303),
.B(n_299),
.C(n_297),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_738),
.B(n_540),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_742),
.A2(n_612),
.B(n_602),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_690),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_664),
.B(n_617),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_L g908 ( 
.A(n_738),
.B(n_540),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_670),
.B(n_617),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_697),
.A2(n_299),
.B(n_293),
.C(n_289),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_672),
.B(n_623),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_673),
.A2(n_293),
.B(n_289),
.C(n_634),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_658),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_767),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_674),
.B(n_710),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_740),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_750),
.B(n_296),
.C(n_333),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_691),
.B(n_544),
.Y(n_918)
);

O2A1O1Ixp5_ASAP7_75t_L g919 ( 
.A1(n_795),
.A2(n_438),
.B(n_435),
.C(n_424),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_779),
.A2(n_544),
.B(n_582),
.C(n_460),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_699),
.B(n_544),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_736),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_660),
.A2(n_582),
.B(n_438),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_781),
.B(n_582),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_660),
.A2(n_582),
.B(n_438),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_815),
.B(n_582),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_753),
.B(n_759),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_690),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_666),
.B(n_321),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_334),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_815),
.B(n_460),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_767),
.B(n_442),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_663),
.A2(n_424),
.B(n_425),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_693),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_747),
.B(n_337),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_820),
.B(n_769),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_757),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_761),
.B(n_339),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_767),
.B(n_797),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_L g940 ( 
.A(n_789),
.B(n_801),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_770),
.B(n_440),
.Y(n_941)
);

BUFx4f_ASAP7_75t_L g942 ( 
.A(n_797),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_775),
.B(n_440),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_752),
.B(n_279),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_663),
.A2(n_424),
.B(n_425),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_803),
.B(n_440),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_677),
.A2(n_444),
.B(n_447),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_676),
.A2(n_424),
.B(n_425),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_728),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_676),
.A2(n_435),
.B(n_438),
.Y(n_950)
);

BUFx12f_ASAP7_75t_L g951 ( 
.A(n_766),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_435),
.B(n_459),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_818),
.A2(n_175),
.B1(n_172),
.B2(n_177),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_679),
.A2(n_435),
.B(n_290),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_698),
.A2(n_279),
.B1(n_216),
.B2(n_459),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_768),
.A2(n_460),
.B(n_444),
.C(n_459),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_797),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_789),
.B(n_444),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_679),
.A2(n_286),
.B(n_184),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_715),
.B(n_279),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_807),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_814),
.B(n_460),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_801),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_769),
.B(n_460),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_693),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_698),
.A2(n_447),
.B1(n_454),
.B2(n_460),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_772),
.B(n_808),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_811),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_787),
.B(n_447),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_796),
.A2(n_454),
.B(n_461),
.C(n_449),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_797),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_715),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_801),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_772),
.B(n_454),
.C(n_217),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_713),
.B(n_182),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_748),
.B(n_442),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_681),
.A2(n_292),
.B(n_189),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_681),
.A2(n_308),
.B(n_191),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_696),
.A2(n_314),
.B(n_193),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_658),
.A2(n_316),
.B1(n_197),
.B2(n_203),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_696),
.A2(n_317),
.B(n_209),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_812),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_819),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_718),
.B(n_188),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_808),
.B(n_6),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_683),
.A2(n_322),
.B(n_214),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_721),
.B(n_213),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_798),
.B(n_7),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_733),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_683),
.A2(n_323),
.B(n_227),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_816),
.B(n_218),
.C(n_237),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_669),
.B(n_241),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_695),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_758),
.B(n_9),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_773),
.B(n_246),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_773),
.B(n_722),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_748),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_695),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_724),
.A2(n_461),
.B(n_449),
.C(n_448),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_731),
.A2(n_330),
.B(n_278),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_784),
.A2(n_338),
.B(n_320),
.Y(n_1001)
);

AO21x1_ASAP7_75t_L g1002 ( 
.A1(n_754),
.A2(n_461),
.B(n_449),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_751),
.B(n_10),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_751),
.B(n_11),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_766),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_743),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_678),
.A2(n_272),
.B(n_269),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_773),
.A2(n_328),
.B1(n_258),
.B2(n_326),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_967),
.A2(n_790),
.B(n_784),
.C(n_799),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_822),
.A2(n_793),
.B(n_744),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_821),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_918),
.A2(n_656),
.B(n_782),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_854),
.A2(n_830),
.B(n_829),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_967),
.A2(n_835),
.B(n_837),
.C(n_893),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_846),
.A2(n_863),
.B(n_857),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_852),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_842),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_878),
.A2(n_915),
.B1(n_870),
.B2(n_1003),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_841),
.A2(n_656),
.B(n_782),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_917),
.A2(n_809),
.B1(n_719),
.B2(n_791),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_845),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_947),
.A2(n_804),
.B(n_796),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_852),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_951),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_851),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_927),
.B(n_868),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_974),
.A2(n_754),
.B(n_799),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_876),
.B(n_791),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_960),
.B(n_800),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_840),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_960),
.B(n_737),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_1002),
.A2(n_790),
.B(n_765),
.C(n_743),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_850),
.B(n_809),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_858),
.A2(n_678),
.B1(n_755),
.B2(n_762),
.C(n_765),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_852),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_870),
.B(n_791),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_856),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_985),
.A2(n_755),
.B(n_762),
.C(n_794),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_949),
.B(n_794),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_1005),
.B(n_791),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_858),
.B(n_791),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_963),
.B(n_817),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_852),
.B(n_708),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_865),
.B(n_802),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_885),
.B(n_788),
.Y(n_1045)
);

AND2x4_ASAP7_75t_SL g1046 ( 
.A(n_963),
.B(n_780),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_856),
.B(n_774),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_834),
.A2(n_771),
.B(n_726),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_955),
.B(n_711),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_875),
.Y(n_1050)
);

OAI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_824),
.A2(n_720),
.B1(n_220),
.B2(n_327),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_974),
.A2(n_461),
.B(n_449),
.C(n_448),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_973),
.B(n_449),
.Y(n_1053)
);

CKINVDCx10_ASAP7_75t_R g1054 ( 
.A(n_897),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_955),
.B(n_13),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_917),
.A2(n_461),
.B1(n_449),
.B2(n_448),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_916),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_885),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_843),
.A2(n_434),
.B(n_430),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_L g1060 ( 
.A1(n_1008),
.A2(n_899),
.B1(n_994),
.B2(n_884),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_836),
.A2(n_434),
.B(n_430),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_838),
.A2(n_461),
.B(n_449),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_937),
.B(n_15),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_914),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_893),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_991),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_878),
.A2(n_461),
.B1(n_449),
.B2(n_448),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_856),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_SL g1069 ( 
.A1(n_1003),
.A2(n_24),
.B(n_27),
.C(n_30),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_922),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_849),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_914),
.B(n_461),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_936),
.A2(n_461),
.B(n_449),
.C(n_448),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_926),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_913),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_942),
.B(n_448),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_942),
.B(n_448),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_949),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_839),
.A2(n_448),
.B(n_442),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_860),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_962),
.B(n_32),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_931),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_966),
.B(n_864),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_833),
.B(n_99),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_861),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_913),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_972),
.Y(n_1087)
);

INVx3_ASAP7_75t_SL g1088 ( 
.A(n_931),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_972),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_847),
.B(n_34),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_957),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_926),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_991),
.A2(n_34),
.B(n_37),
.C(n_42),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_SL g1094 ( 
.A(n_825),
.B(n_42),
.C(n_44),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_961),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_45),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_994),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_944),
.B(n_826),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1004),
.A2(n_983),
.B1(n_982),
.B2(n_968),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1004),
.A2(n_997),
.B1(n_828),
.B2(n_889),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_879),
.A2(n_448),
.B1(n_442),
.B2(n_327),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_969),
.B(n_45),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_972),
.B(n_442),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_957),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_853),
.A2(n_220),
.B1(n_324),
.B2(n_327),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_944),
.B(n_46),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_906),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_973),
.B(n_49),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_869),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_971),
.B(n_49),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_L g1113 ( 
.A1(n_844),
.A2(n_442),
.B(n_53),
.C(n_55),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_928),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_988),
.A2(n_442),
.B1(n_327),
.B2(n_324),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_872),
.A2(n_442),
.B(n_327),
.C(n_324),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_877),
.B(n_51),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_848),
.A2(n_434),
.B(n_430),
.Y(n_1118)
);

AOI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1007),
.A2(n_324),
.B(n_220),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_934),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_997),
.A2(n_324),
.B1(n_220),
.B2(n_63),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1006),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_872),
.A2(n_434),
.B(n_430),
.C(n_63),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_972),
.B(n_434),
.Y(n_1124)
);

AND2x2_ASAP7_75t_SL g1125 ( 
.A(n_940),
.B(n_908),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_880),
.A2(n_51),
.B1(n_57),
.B2(n_64),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_873),
.A2(n_434),
.B(n_430),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_SL g1128 ( 
.A(n_930),
.B(n_57),
.C(n_66),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_869),
.B(n_434),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_939),
.B(n_434),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_891),
.A2(n_434),
.B1(n_430),
.B2(n_79),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_831),
.A2(n_430),
.B(n_76),
.C(n_86),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_939),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_996),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_998),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_941),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_989),
.B(n_430),
.C(n_89),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_904),
.B(n_430),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_953),
.B(n_73),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_943),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_929),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_823),
.A2(n_90),
.B(n_96),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_912),
.A2(n_100),
.B(n_102),
.C(n_105),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_946),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_921),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_896),
.A2(n_112),
.B1(n_117),
.B2(n_124),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_976),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_976),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_L g1150 ( 
.A(n_903),
.B(n_125),
.C(n_136),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_844),
.A2(n_143),
.B(n_147),
.C(n_157),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_827),
.A2(n_158),
.B1(n_169),
.B2(n_170),
.Y(n_1152)
);

NOR2x1p5_ASAP7_75t_L g1153 ( 
.A(n_935),
.B(n_938),
.Y(n_1153)
);

AOI222xp33_ASAP7_75t_L g1154 ( 
.A1(n_995),
.A2(n_874),
.B1(n_901),
.B2(n_892),
.C1(n_909),
.C2(n_907),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_859),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_964),
.B(n_924),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_904),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_992),
.B(n_958),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_932),
.B(n_920),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_862),
.A2(n_910),
.B(n_855),
.C(n_898),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_911),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_975),
.A2(n_987),
.B1(n_984),
.B2(n_888),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_867),
.A2(n_832),
.B(n_866),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_980),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1062),
.A2(n_900),
.B(n_886),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_1064),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_932),
.B1(n_986),
.B2(n_990),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_1018),
.A2(n_1014),
.B(n_1100),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1014),
.A2(n_871),
.B1(n_981),
.B2(n_979),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1107),
.A2(n_881),
.B1(n_952),
.B2(n_977),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1031),
.A2(n_1051),
.B1(n_1090),
.B2(n_1033),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1013),
.A2(n_900),
.B(n_999),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1058),
.B(n_956),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1026),
.B(n_978),
.Y(n_1174)
);

NOR4xp25_ASAP7_75t_L g1175 ( 
.A(n_1065),
.B(n_902),
.C(n_905),
.D(n_970),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_1026),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1082),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1027),
.A2(n_895),
.A3(n_883),
.B(n_925),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1079),
.A2(n_923),
.B(n_919),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1108),
.A2(n_959),
.B1(n_1001),
.B2(n_882),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1066),
.A2(n_919),
.B(n_970),
.C(n_1000),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1011),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1090),
.A2(n_890),
.B1(n_887),
.B2(n_954),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1052),
.A2(n_933),
.A3(n_945),
.B(n_948),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1020),
.B(n_950),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1091),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1058),
.B(n_1092),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1015),
.A2(n_1101),
.B(n_1119),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1009),
.A2(n_1032),
.B(n_1113),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1009),
.A2(n_1066),
.B(n_1093),
.C(n_1041),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1163),
.A2(n_1116),
.A3(n_1038),
.B(n_1073),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1059),
.A2(n_1061),
.B(n_1118),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1024),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1048),
.A2(n_1127),
.B(n_1022),
.Y(n_1194)
);

NOR2x1_ASAP7_75t_L g1195 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1047),
.B(n_1064),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_SL g1197 ( 
.A1(n_1132),
.A2(n_1123),
.B(n_1162),
.C(n_1036),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1142),
.B(n_1088),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1093),
.A2(n_1094),
.B(n_1153),
.C(n_1065),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1017),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1148),
.B(n_1064),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1054),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1010),
.A2(n_1129),
.B(n_1019),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1012),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1125),
.A2(n_1155),
.B(n_1141),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1064),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1106),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1125),
.A2(n_1155),
.B(n_1137),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1044),
.B(n_1158),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1098),
.B(n_1088),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1021),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1094),
.A2(n_1033),
.B(n_1111),
.C(n_1160),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1044),
.B(n_1145),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1035),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1032),
.A2(n_1143),
.B(n_1151),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1051),
.A2(n_1097),
.B1(n_1083),
.B2(n_1055),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1159),
.A2(n_1111),
.B(n_1152),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1078),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1035),
.B(n_1087),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1159),
.A2(n_1156),
.B(n_1151),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1025),
.Y(n_1221)
);

NAND2x1_ASAP7_75t_L g1222 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1028),
.A2(n_1029),
.B(n_1103),
.C(n_1113),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1067),
.A2(n_1139),
.B(n_1076),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1030),
.Y(n_1225)
);

NOR4xp25_ASAP7_75t_L g1226 ( 
.A(n_1126),
.B(n_1102),
.C(n_1121),
.D(n_1063),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1146),
.A2(n_1161),
.B(n_1042),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_1072),
.B(n_1154),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1050),
.B(n_1096),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1112),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1139),
.A2(n_1124),
.B(n_1105),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1099),
.B(n_1081),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1161),
.A2(n_1115),
.B(n_1104),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1122),
.A2(n_1077),
.B(n_1147),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1034),
.Y(n_1235)
);

INVx8_ASAP7_75t_L g1236 ( 
.A(n_1035),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1057),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_1074),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1138),
.A2(n_1049),
.B(n_1144),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1110),
.B(n_1157),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1130),
.A2(n_1086),
.B(n_1075),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1148),
.B(n_1039),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1130),
.A2(n_1043),
.B(n_1150),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1077),
.A2(n_1117),
.B(n_1045),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1112),
.A2(n_1128),
.B1(n_1056),
.B2(n_1102),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1047),
.A2(n_1148),
.B(n_1069),
.Y(n_1246)
);

OAI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1128),
.A2(n_1040),
.B1(n_1068),
.B2(n_1037),
.C(n_1047),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1133),
.A2(n_1149),
.B(n_1046),
.C(n_1135),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1136),
.A2(n_1134),
.B(n_1053),
.C(n_1074),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1037),
.B(n_1068),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1134),
.B(n_1060),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1053),
.A2(n_1085),
.B(n_1120),
.C(n_1114),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1148),
.B(n_1035),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1071),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1084),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1023),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1023),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1080),
.A2(n_1095),
.B(n_1109),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1089),
.Y(n_1259)
);

AOI31xp67_ASAP7_75t_L g1260 ( 
.A1(n_1084),
.A2(n_1089),
.A3(n_1023),
.B(n_1016),
.Y(n_1260)
);

OAI22x1_ASAP7_75t_L g1261 ( 
.A1(n_1016),
.A2(n_1008),
.B1(n_560),
.B2(n_967),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1089),
.B(n_1023),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1164),
.A2(n_967),
.B1(n_560),
.B2(n_654),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1062),
.A2(n_1079),
.B(n_1059),
.Y(n_1265)
);

INVxp67_ASAP7_75t_SL g1266 ( 
.A(n_1026),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1058),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1094),
.B(n_967),
.C(n_1014),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1026),
.B(n_735),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1026),
.B(n_735),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1078),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1164),
.B(n_522),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1164),
.B(n_522),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1018),
.A2(n_967),
.B1(n_714),
.B2(n_822),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1014),
.A2(n_967),
.B(n_917),
.C(n_1018),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1163),
.A2(n_1119),
.B(n_1013),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1027),
.A2(n_1002),
.A3(n_947),
.B(n_1052),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1026),
.B(n_735),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1027),
.A2(n_1002),
.A3(n_947),
.B(n_1052),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1058),
.B(n_963),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1011),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1018),
.A2(n_967),
.B(n_1014),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1027),
.A2(n_1002),
.A3(n_947),
.B(n_1052),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1011),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1058),
.B(n_963),
.Y(n_1286)
);

NOR4xp25_ASAP7_75t_L g1287 ( 
.A(n_1065),
.B(n_1066),
.C(n_1093),
.D(n_1014),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1054),
.Y(n_1288)
);

NAND3x1_ASAP7_75t_L g1289 ( 
.A(n_1090),
.B(n_967),
.C(n_917),
.Y(n_1289)
);

AOI31xp67_ASAP7_75t_L g1290 ( 
.A1(n_1156),
.A2(n_1159),
.A3(n_1115),
.B(n_1056),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1026),
.B(n_735),
.Y(n_1291)
);

OAI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1090),
.A2(n_1008),
.B1(n_560),
.B2(n_967),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1051),
.B(n_878),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1026),
.B(n_735),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1018),
.A2(n_967),
.B1(n_822),
.B2(n_654),
.Y(n_1295)
);

INVx8_ASAP7_75t_L g1296 ( 
.A(n_1024),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1058),
.B(n_963),
.Y(n_1298)
);

BUFx2_ASAP7_75t_R g1299 ( 
.A(n_1070),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1026),
.B(n_735),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1027),
.A2(n_1002),
.A3(n_947),
.B(n_1052),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_1026),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1026),
.B(n_735),
.Y(n_1304)
);

CKINVDCx14_ASAP7_75t_R g1305 ( 
.A(n_1024),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1014),
.B(n_967),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1058),
.B(n_963),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1027),
.A2(n_1002),
.A3(n_947),
.B(n_1052),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1026),
.B(n_735),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_SL g1310 ( 
.A1(n_1108),
.A2(n_985),
.B(n_822),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1026),
.B(n_735),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1018),
.A2(n_967),
.B(n_1014),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1119),
.A2(n_1027),
.B(n_854),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1079),
.A2(n_1163),
.B(n_1013),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1026),
.B(n_735),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1070),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1026),
.B(n_735),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1024),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1018),
.A2(n_967),
.B1(n_822),
.B2(n_654),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1018),
.A2(n_1015),
.B(n_822),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1062),
.A2(n_1079),
.B(n_1059),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1062),
.A2(n_1079),
.B(n_1059),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1026),
.B(n_735),
.Y(n_1325)
);

CKINVDCx6p67_ASAP7_75t_R g1326 ( 
.A(n_1202),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1296),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1236),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1296),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1238),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1263),
.A2(n_1276),
.B(n_1274),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1293),
.A2(n_1216),
.B1(n_1268),
.B2(n_1245),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1236),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1182),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1293),
.A2(n_1292),
.B1(n_1171),
.B2(n_1261),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1275),
.A2(n_1289),
.B1(n_1230),
.B2(n_1312),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1200),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1291),
.B(n_1316),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1218),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1211),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1275),
.A2(n_1268),
.B1(n_1283),
.B2(n_1312),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1221),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_SL g1343 ( 
.A(n_1253),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1283),
.A2(n_1321),
.B1(n_1295),
.B2(n_1311),
.Y(n_1344)
);

INVx5_ASAP7_75t_L g1345 ( 
.A(n_1236),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1273),
.A2(n_1306),
.B1(n_1212),
.B2(n_1199),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1269),
.A2(n_1325),
.B1(n_1309),
.B2(n_1294),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1296),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1305),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1237),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1216),
.A2(n_1168),
.B1(n_1232),
.B2(n_1251),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1166),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1271),
.A2(n_1319),
.B1(n_1279),
.B2(n_1300),
.Y(n_1353)
);

BUFx4f_ASAP7_75t_SL g1354 ( 
.A(n_1255),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1288),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1174),
.A2(n_1266),
.B1(n_1209),
.B2(n_1240),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1193),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1320),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1225),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1304),
.A2(n_1198),
.B1(n_1247),
.B2(n_1302),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1213),
.B(n_1186),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1228),
.A2(n_1254),
.B1(n_1217),
.B2(n_1235),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1282),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1205),
.A2(n_1208),
.B1(n_1189),
.B2(n_1270),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1272),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1210),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1285),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1176),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1190),
.A2(n_1207),
.B1(n_1322),
.B2(n_1303),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1258),
.A2(n_1302),
.B1(n_1176),
.B2(n_1170),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1317),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1250),
.A2(n_1173),
.B1(n_1189),
.B2(n_1239),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1287),
.A2(n_1297),
.B1(n_1264),
.B2(n_1313),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1318),
.A2(n_1173),
.B1(n_1223),
.B2(n_1224),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1239),
.A2(n_1177),
.B1(n_1196),
.B2(n_1242),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1259),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1287),
.A2(n_1226),
.B1(n_1220),
.B2(n_1314),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1166),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1267),
.A2(n_1167),
.B1(n_1241),
.B2(n_1246),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1227),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1299),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1314),
.B2(n_1169),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1187),
.B(n_1267),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1195),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1188),
.A2(n_1196),
.B1(n_1183),
.B2(n_1166),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1249),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1201),
.A2(n_1180),
.B1(n_1185),
.B2(n_1233),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1262),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1183),
.A2(n_1204),
.B1(n_1298),
.B2(n_1281),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1248),
.A2(n_1222),
.B1(n_1307),
.B2(n_1286),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1226),
.A2(n_1277),
.B1(n_1243),
.B2(n_1215),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_SL g1392 ( 
.A(n_1286),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1206),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1206),
.A2(n_1214),
.B1(n_1231),
.B2(n_1219),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1252),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1257),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_1206),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1256),
.Y(n_1398)
);

CKINVDCx11_ASAP7_75t_R g1399 ( 
.A(n_1256),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1307),
.A2(n_1244),
.B1(n_1256),
.B2(n_1172),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1277),
.A2(n_1290),
.B1(n_1172),
.B2(n_1234),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1197),
.A2(n_1310),
.B1(n_1214),
.B2(n_1260),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1219),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1178),
.Y(n_1404)
);

BUFx8_ASAP7_75t_L g1405 ( 
.A(n_1175),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1278),
.Y(n_1406)
);

BUFx10_ASAP7_75t_L g1407 ( 
.A(n_1175),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1194),
.B(n_1179),
.Y(n_1408)
);

BUFx8_ASAP7_75t_L g1409 ( 
.A(n_1278),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1280),
.B(n_1284),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1203),
.A2(n_1192),
.B1(n_1165),
.B2(n_1324),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1280),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1265),
.A2(n_1323),
.B1(n_1181),
.B2(n_1191),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1284),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1315),
.A2(n_1191),
.B1(n_1284),
.B2(n_1301),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1308),
.A2(n_967),
.B(n_1018),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1184),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1184),
.A2(n_967),
.B1(n_1275),
.B2(n_1289),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1202),
.Y(n_1419)
);

AOI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1292),
.A2(n_967),
.B(n_1276),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1289),
.A2(n_967),
.B(n_1276),
.Y(n_1421)
);

BUFx10_ASAP7_75t_L g1422 ( 
.A(n_1288),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1202),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1202),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1229),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1229),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1293),
.A2(n_698),
.B1(n_439),
.B2(n_1216),
.Y(n_1427)
);

INVx6_ASAP7_75t_L g1428 ( 
.A(n_1166),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1166),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1275),
.A2(n_967),
.B1(n_1289),
.B2(n_1263),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1275),
.A2(n_967),
.B1(n_1289),
.B2(n_1263),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1229),
.Y(n_1432)
);

INVx8_ASAP7_75t_L g1433 ( 
.A(n_1236),
.Y(n_1433)
);

BUFx2_ASAP7_75t_SL g1434 ( 
.A(n_1255),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1291),
.B(n_1316),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1293),
.A2(n_439),
.B1(n_698),
.B2(n_1292),
.Y(n_1436)
);

BUFx8_ASAP7_75t_SL g1437 ( 
.A(n_1193),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1293),
.A2(n_698),
.B1(n_439),
.B2(n_1216),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1202),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1293),
.A2(n_439),
.B1(n_698),
.B2(n_1292),
.Y(n_1440)
);

OAI22x1_ASAP7_75t_L g1441 ( 
.A1(n_1275),
.A2(n_1008),
.B1(n_1240),
.B2(n_967),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1168),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1291),
.B(n_1316),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1288),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1275),
.A2(n_967),
.B1(n_1289),
.B2(n_1263),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1236),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1293),
.A2(n_698),
.B1(n_439),
.B2(n_1216),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1209),
.B(n_1291),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1293),
.A2(n_698),
.B1(n_439),
.B2(n_1216),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1229),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1166),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1293),
.A2(n_439),
.B1(n_698),
.B2(n_1292),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1229),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1330),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1410),
.B(n_1407),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1368),
.B(n_1354),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1361),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1338),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1404),
.Y(n_1462)
);

NAND2x1_ASAP7_75t_L g1463 ( 
.A(n_1416),
.B(n_1374),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1407),
.B(n_1442),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1380),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1334),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_1413),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1337),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1415),
.A2(n_1385),
.B(n_1418),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1415),
.A2(n_1385),
.B(n_1364),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1340),
.Y(n_1472)
);

AO21x1_ASAP7_75t_SL g1473 ( 
.A1(n_1421),
.A2(n_1372),
.B(n_1420),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1342),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1417),
.A2(n_1387),
.B(n_1362),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1350),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_SL g1477 ( 
.A1(n_1430),
.A2(n_1431),
.B(n_1445),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1363),
.Y(n_1478)
);

BUFx4f_ASAP7_75t_L g1479 ( 
.A(n_1428),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1437),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1388),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1367),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1409),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1339),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1378),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1409),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1354),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1417),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1369),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1408),
.A2(n_1379),
.B(n_1389),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1414),
.Y(n_1491)
);

CKINVDCx6p67_ASAP7_75t_R g1492 ( 
.A(n_1327),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1386),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1377),
.B(n_1435),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1425),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1428),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1426),
.Y(n_1497)
);

AO21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1351),
.A2(n_1400),
.B(n_1382),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1405),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1432),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1429),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1450),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1335),
.A2(n_1395),
.B(n_1370),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1405),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1429),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1429),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1377),
.B(n_1443),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1336),
.B(n_1448),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1453),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1364),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1341),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1396),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1341),
.B(n_1356),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1451),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1366),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1365),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1346),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1441),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1344),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1344),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1391),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1391),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1375),
.A2(n_1390),
.B(n_1383),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1373),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1373),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1329),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1401),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1333),
.Y(n_1528)
);

CKINVDCx12_ASAP7_75t_R g1529 ( 
.A(n_1343),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1401),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1332),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1345),
.B(n_1446),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1402),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1331),
.B(n_1447),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1345),
.B(n_1446),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1352),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1402),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1427),
.B(n_1438),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1360),
.B(n_1452),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1381),
.B(n_1349),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1394),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1394),
.Y(n_1542)
);

AO22x2_ASAP7_75t_L g1543 ( 
.A1(n_1427),
.A2(n_1449),
.B1(n_1447),
.B2(n_1438),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1484),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1534),
.A2(n_1436),
.B1(n_1440),
.B2(n_1449),
.C(n_1434),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1527),
.A2(n_1403),
.B(n_1384),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1534),
.B(n_1365),
.C(n_1393),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1460),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1457),
.B(n_1484),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1458),
.B(n_1326),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1457),
.B(n_1376),
.Y(n_1551)
);

AOI22x1_ASAP7_75t_SL g1552 ( 
.A1(n_1526),
.A2(n_1439),
.B1(n_1424),
.B2(n_1355),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1470),
.B(n_1399),
.Y(n_1553)
);

BUFx5_ASAP7_75t_L g1554 ( 
.A(n_1489),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1499),
.A2(n_1504),
.B1(n_1516),
.B2(n_1517),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1484),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_SL g1557 ( 
.A(n_1492),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_SL g1558 ( 
.A1(n_1477),
.A2(n_1392),
.B(n_1348),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1470),
.B(n_1398),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1470),
.B(n_1345),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1481),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1455),
.B(n_1397),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1494),
.B(n_1328),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_R g1564 ( 
.A(n_1538),
.B(n_1357),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_SL g1565 ( 
.A(n_1473),
.B(n_1328),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1471),
.B(n_1371),
.Y(n_1566)
);

BUFx8_ASAP7_75t_L g1567 ( 
.A(n_1516),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1462),
.B(n_1358),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1538),
.A2(n_1433),
.B(n_1359),
.C(n_1422),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_SL g1570 ( 
.A1(n_1463),
.A2(n_1489),
.B(n_1513),
.C(n_1511),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1468),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1467),
.A2(n_1433),
.B(n_1422),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1463),
.A2(n_1433),
.B(n_1423),
.C(n_1419),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1461),
.B(n_1444),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1513),
.A2(n_1531),
.B(n_1539),
.C(n_1519),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1507),
.B(n_1515),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1543),
.A2(n_1510),
.B(n_1469),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1511),
.A2(n_1519),
.B(n_1520),
.Y(n_1578)
);

INVx5_ASAP7_75t_SL g1579 ( 
.A(n_1492),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1472),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1543),
.A2(n_1531),
.B1(n_1524),
.B2(n_1525),
.C(n_1521),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1468),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1543),
.A2(n_1520),
.B1(n_1524),
.B2(n_1525),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1464),
.B(n_1485),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1508),
.B(n_1472),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1543),
.A2(n_1539),
.B1(n_1499),
.B2(n_1504),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_SL g1587 ( 
.A1(n_1487),
.A2(n_1510),
.B(n_1533),
.C(n_1537),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1464),
.B(n_1485),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1518),
.A2(n_1522),
.B(n_1521),
.C(n_1533),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1495),
.B(n_1497),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1474),
.B(n_1478),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1503),
.A2(n_1498),
.B1(n_1473),
.B2(n_1522),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1518),
.A2(n_1537),
.B(n_1530),
.C(n_1527),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1474),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1530),
.A2(n_1456),
.B1(n_1459),
.B2(n_1479),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1469),
.A2(n_1503),
.B1(n_1493),
.B2(n_1491),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1467),
.A2(n_1490),
.B(n_1523),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1523),
.A2(n_1490),
.B(n_1542),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1466),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1491),
.B(n_1482),
.Y(n_1600)
);

A2O1A1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1541),
.A2(n_1542),
.B(n_1479),
.C(n_1493),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1541),
.A2(n_1503),
.B(n_1475),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1476),
.B(n_1469),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1496),
.A2(n_1514),
.A3(n_1506),
.B1(n_1505),
.B2(n_1501),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1571),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1545),
.A2(n_1581),
.B1(n_1583),
.B2(n_1503),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1582),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1603),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1554),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1495),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1564),
.A2(n_1475),
.B1(n_1529),
.B2(n_1509),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1560),
.B(n_1465),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1594),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1548),
.B(n_1500),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1465),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1577),
.A2(n_1498),
.B1(n_1475),
.B2(n_1502),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1561),
.B(n_1488),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1553),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1512),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1590),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1560),
.B(n_1475),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1488),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1604),
.Y(n_1626)
);

NOR2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1592),
.A2(n_1497),
.B1(n_1500),
.B2(n_1502),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1544),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1566),
.B(n_1540),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1599),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1549),
.B(n_1454),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1576),
.B(n_1454),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1609),
.B(n_1559),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1605),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1621),
.B(n_1626),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

INVx5_ASAP7_75t_L g1639 ( 
.A(n_1609),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1619),
.Y(n_1640)
);

CKINVDCx16_ASAP7_75t_R g1641 ( 
.A(n_1619),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1622),
.B(n_1598),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1619),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1626),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1611),
.A2(n_1602),
.B(n_1593),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1606),
.A2(n_1586),
.B1(n_1592),
.B2(n_1596),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1597),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1626),
.B(n_1604),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

OAI31xp33_ASAP7_75t_L g1651 ( 
.A1(n_1606),
.A2(n_1575),
.A3(n_1589),
.B(n_1593),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1622),
.B(n_1584),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1597),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1619),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1612),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1630),
.A2(n_1550),
.B(n_1566),
.C(n_1573),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1616),
.A2(n_1578),
.B1(n_1562),
.B2(n_1547),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1607),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1607),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1617),
.B(n_1572),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1616),
.A2(n_1575),
.B1(n_1589),
.B2(n_1564),
.C(n_1587),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1632),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1628),
.A2(n_1587),
.B1(n_1570),
.B2(n_1569),
.C(n_1595),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1615),
.B(n_1588),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1634),
.B(n_1620),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1624),
.A2(n_1570),
.B(n_1601),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1613),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1674)
);

INVxp33_ASAP7_75t_SL g1675 ( 
.A(n_1667),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1645),
.B(n_1618),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1636),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_1625),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1638),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1638),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1650),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1640),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1650),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1661),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1627),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1662),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1625),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1652),
.B(n_1625),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1662),
.Y(n_1694)
);

INVx4_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1640),
.B(n_1633),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1670),
.B(n_1611),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1663),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1633),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1646),
.A2(n_1624),
.B1(n_1611),
.B2(n_1546),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1644),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1663),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1637),
.B(n_1614),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1654),
.B(n_1633),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1648),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1665),
.A2(n_1631),
.B(n_1555),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1671),
.Y(n_1709)
);

AND3x2_ASAP7_75t_L g1710 ( 
.A(n_1651),
.B(n_1631),
.C(n_1568),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1673),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1684),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1673),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1679),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1667),
.C(n_1658),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1674),
.B(n_1637),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1684),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1675),
.B(n_1649),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1687),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1685),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1675),
.A2(n_1658),
.B(n_1649),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1698),
.A2(n_1665),
.B1(n_1647),
.B2(n_1659),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1677),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1687),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1678),
.B(n_1657),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1669),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1698),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1678),
.B(n_1657),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1692),
.B(n_1693),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1677),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1696),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1690),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1690),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1691),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1691),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1694),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_SL g1744 ( 
.A1(n_1686),
.A2(n_1573),
.B(n_1569),
.C(n_1670),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1702),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1708),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1708),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

OAI31xp33_ASAP7_75t_L g1750 ( 
.A1(n_1698),
.A2(n_1651),
.A3(n_1647),
.B(n_1659),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1709),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1697),
.B(n_1669),
.Y(n_1753)
);

OAI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1716),
.A2(n_1701),
.B(n_1706),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1672),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1750),
.B(n_1723),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1717),
.B(n_1695),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1750),
.B(n_1697),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1726),
.B(n_1672),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1737),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1723),
.B(n_1700),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1711),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1728),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1711),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1739),
.B(n_1557),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1713),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1737),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1713),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.B(n_1676),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1676),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1724),
.A2(n_1480),
.B(n_1689),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1736),
.B(n_1653),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1714),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1557),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1725),
.B(n_1695),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1712),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1746),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1725),
.B(n_1695),
.Y(n_1778)
);

NAND2x1_ASAP7_75t_L g1779 ( 
.A(n_1728),
.B(n_1689),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1718),
.B(n_1700),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1714),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_SL g1782 ( 
.A(n_1732),
.B(n_1721),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1746),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1715),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1715),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1721),
.B(n_1722),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1731),
.B(n_1705),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1722),
.B(n_1705),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1733),
.B(n_1653),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1776),
.B(n_1753),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1768),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1784),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1756),
.A2(n_1646),
.B1(n_1710),
.B2(n_1656),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1784),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1755),
.B(n_1730),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1758),
.B(n_1655),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1762),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1732),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1755),
.B(n_1730),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1763),
.B(n_1751),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1754),
.B(n_1579),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1782),
.A2(n_1653),
.B(n_1720),
.Y(n_1803)
);

AOI222xp33_ASAP7_75t_L g1804 ( 
.A1(n_1761),
.A2(n_1656),
.B1(n_1655),
.B2(n_1743),
.C1(n_1742),
.C2(n_1720),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1782),
.A2(n_1646),
.B1(n_1656),
.B2(n_1655),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1767),
.B(n_1751),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1779),
.B(n_1734),
.C(n_1727),
.Y(n_1808)
);

AOI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1777),
.A2(n_1734),
.B(n_1727),
.Y(n_1809)
);

OAI32xp33_ASAP7_75t_L g1810 ( 
.A1(n_1774),
.A2(n_1752),
.A3(n_1749),
.B1(n_1748),
.B2(n_1747),
.Y(n_1810)
);

AOI322xp5_ASAP7_75t_L g1811 ( 
.A1(n_1786),
.A2(n_1729),
.A3(n_1664),
.B1(n_1623),
.B2(n_1628),
.C1(n_1745),
.C2(n_1743),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1760),
.B(n_1735),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1764),
.Y(n_1813)
);

AOI222xp33_ASAP7_75t_L g1814 ( 
.A1(n_1786),
.A2(n_1752),
.B1(n_1749),
.B2(n_1748),
.C1(n_1747),
.C2(n_1745),
.Y(n_1814)
);

INVxp67_ASAP7_75t_L g1815 ( 
.A(n_1765),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1800),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1799),
.B(n_1760),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1812),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1805),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1800),
.Y(n_1820)
);

AOI21xp33_ASAP7_75t_L g1821 ( 
.A1(n_1810),
.A2(n_1783),
.B(n_1777),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1806),
.A2(n_1771),
.B(n_1799),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1791),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1792),
.Y(n_1825)
);

AO21x1_ASAP7_75t_SL g1826 ( 
.A1(n_1807),
.A2(n_1787),
.B(n_1773),
.Y(n_1826)
);

AOI311xp33_ASAP7_75t_L g1827 ( 
.A1(n_1790),
.A2(n_1766),
.A3(n_1785),
.B(n_1781),
.C(n_1788),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1802),
.A2(n_1779),
.B(n_1757),
.C(n_1775),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1796),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1811),
.B(n_1814),
.C(n_1794),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1801),
.B(n_1780),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1805),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1759),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1793),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1802),
.A2(n_1772),
.B1(n_1759),
.B2(n_1769),
.C(n_1770),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1831),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1830),
.A2(n_1823),
.B1(n_1829),
.B2(n_1820),
.Y(n_1837)
);

AOI32xp33_ASAP7_75t_L g1838 ( 
.A1(n_1827),
.A2(n_1801),
.A3(n_1795),
.B1(n_1813),
.B2(n_1798),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1831),
.B(n_1775),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1816),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1829),
.A2(n_1804),
.B1(n_1646),
.B2(n_1778),
.Y(n_1841)
);

XNOR2xp5_ASAP7_75t_L g1842 ( 
.A(n_1817),
.B(n_1552),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1816),
.A2(n_1815),
.B1(n_1803),
.B2(n_1778),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1817),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1820),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1819),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1819),
.Y(n_1847)
);

OAI21xp33_ASAP7_75t_L g1848 ( 
.A1(n_1822),
.A2(n_1757),
.B(n_1808),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1836),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1846),
.B(n_1835),
.C(n_1821),
.Y(n_1850)
);

AOI211x1_ASAP7_75t_L g1851 ( 
.A1(n_1848),
.A2(n_1828),
.B(n_1818),
.C(n_1809),
.Y(n_1851)
);

NOR3x1_ASAP7_75t_L g1852 ( 
.A(n_1847),
.B(n_1833),
.C(n_1825),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1842),
.B(n_1832),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1839),
.Y(n_1854)
);

NAND4xp25_ASAP7_75t_SL g1855 ( 
.A(n_1837),
.B(n_1833),
.C(n_1826),
.D(n_1834),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1843),
.A2(n_1832),
.B(n_1824),
.Y(n_1856)
);

NOR3xp33_ASAP7_75t_L g1857 ( 
.A(n_1840),
.B(n_1783),
.C(n_1772),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1844),
.B(n_1769),
.Y(n_1858)
);

AOI322xp5_ASAP7_75t_L g1859 ( 
.A1(n_1841),
.A2(n_1826),
.A3(n_1623),
.B1(n_1664),
.B2(n_1742),
.C1(n_1741),
.C2(n_1740),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1845),
.A2(n_1646),
.B1(n_1789),
.B2(n_1770),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1850),
.A2(n_1789),
.B1(n_1843),
.B2(n_1740),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1853),
.A2(n_1838),
.B(n_1579),
.C(n_1738),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1855),
.A2(n_1741),
.B(n_1738),
.C(n_1735),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1856),
.A2(n_1551),
.B(n_1568),
.C(n_1664),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1854),
.B(n_1666),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

OAI211xp5_ASAP7_75t_SL g1867 ( 
.A1(n_1862),
.A2(n_1861),
.B(n_1863),
.C(n_1859),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1864),
.B(n_1857),
.Y(n_1868)
);

AOI21xp33_ASAP7_75t_SL g1869 ( 
.A1(n_1861),
.A2(n_1858),
.B(n_1849),
.Y(n_1869)
);

AOI21xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1861),
.A2(n_1852),
.B(n_1860),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1861),
.A2(n_1851),
.B1(n_1666),
.B2(n_1702),
.C(n_1568),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1867),
.B(n_1579),
.Y(n_1872)
);

NAND4xp75_ASAP7_75t_L g1873 ( 
.A(n_1866),
.B(n_1623),
.C(n_1574),
.D(n_1562),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1868),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1871),
.A2(n_1567),
.B1(n_1635),
.B2(n_1546),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1869),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1874),
.A2(n_1870),
.B1(n_1567),
.B2(n_1635),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1876),
.Y(n_1878)
);

AOI322xp5_ASAP7_75t_L g1879 ( 
.A1(n_1872),
.A2(n_1608),
.A3(n_1660),
.B1(n_1635),
.B2(n_1612),
.C1(n_1614),
.C2(n_1563),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1878),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1877),
.B1(n_1875),
.B2(n_1873),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1881),
.B(n_1879),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1881),
.A2(n_1567),
.B1(n_1529),
.B2(n_1683),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1882),
.B(n_1669),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1883),
.B(n_1660),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_SL g1886 ( 
.A1(n_1884),
.A2(n_1558),
.B(n_1565),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1885),
.A2(n_1703),
.B1(n_1699),
.B2(n_1682),
.Y(n_1887)
);

AOI21xp33_ASAP7_75t_L g1888 ( 
.A1(n_1887),
.A2(n_1885),
.B(n_1486),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1888),
.A2(n_1886),
.B(n_1635),
.Y(n_1889)
);

XNOR2xp5_ASAP7_75t_L g1890 ( 
.A(n_1889),
.B(n_1483),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_R g1891 ( 
.A1(n_1890),
.A2(n_1639),
.B1(n_1681),
.B2(n_1635),
.C(n_1668),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_1556),
.B(n_1532),
.C(n_1535),
.Y(n_1892)
);


endmodule