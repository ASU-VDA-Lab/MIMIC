module fake_jpeg_16155_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_41),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_28),
.B1(n_14),
.B2(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_30),
.B1(n_28),
.B2(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_15),
.B1(n_22),
.B2(n_26),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_22),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_39),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_2),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_23),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_72),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_20),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_39),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_76),
.C(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_56),
.B1(n_53),
.B2(n_2),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_36),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_15),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_2),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_41),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_66),
.C(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_71),
.B1(n_77),
.B2(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

XOR2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_68),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_32),
.B(n_29),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_110),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_74),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_85),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_78),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.C(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_69),
.B1(n_72),
.B2(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_116),
.B1(n_101),
.B2(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_91),
.B1(n_93),
.B2(n_97),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_40),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_113),
.Y(n_129)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_104),
.B1(n_105),
.B2(n_8),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_115),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

AOI31xp67_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_118),
.A3(n_112),
.B(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_5),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_40),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.C(n_29),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_41),
.C(n_29),
.Y(n_133)
);

AOI21x1_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_126),
.B(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_128),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_6),
.B(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_6),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_139),
.B(n_12),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_32),
.CI(n_135),
.CON(n_145),
.SN(n_145)
);


endmodule