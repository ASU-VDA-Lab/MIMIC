module fake_jpeg_5883_n_101 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_12),
.B(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_10),
.B1(n_12),
.B2(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_18),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_42),
.B(n_25),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_29),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_49),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_31),
.B1(n_35),
.B2(n_27),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_37),
.B1(n_42),
.B2(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_47),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_20),
.C(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_45),
.B1(n_44),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_54),
.B1(n_59),
.B2(n_61),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_20),
.C(n_1),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_76),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_54),
.B(n_1),
.Y(n_71)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_0),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_16),
.B1(n_11),
.B2(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NAND4xp25_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_24),
.C(n_20),
.D(n_11),
.Y(n_74)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_69),
.B(n_66),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_9),
.C(n_3),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_67),
.A3(n_9),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_84),
.C(n_77),
.Y(n_86)
);

XNOR2x1_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_74),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.C(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_73),
.B1(n_83),
.B2(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_70),
.C(n_80),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_92),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_2),
.B(n_6),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_93),
.Y(n_101)
);


endmodule