module fake_jpeg_12943_n_97 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_54),
.B1(n_39),
.B2(n_20),
.Y(n_61)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_40),
.B1(n_41),
.B2(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_57),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_36),
.B(n_39),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_72),
.B(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_2),
.B(n_3),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_30),
.B(n_28),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_50),
.C(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_49),
.B1(n_7),
.B2(n_10),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_13),
.B1(n_21),
.B2(n_22),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_70),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_63),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_79),
.B1(n_81),
.B2(n_73),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_85),
.B(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_88),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_87),
.Y(n_97)
);


endmodule