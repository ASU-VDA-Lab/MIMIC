module fake_jpeg_9830_n_110 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_51),
.B(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_38),
.B1(n_17),
.B2(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_57),
.C(n_11),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_58),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_13),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_61),
.B(n_65),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_19),
.B(n_39),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_39),
.B(n_32),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_2),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_54),
.C(n_57),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.C(n_12),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_21),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_55),
.B(n_44),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_15),
.B1(n_13),
.B2(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_82),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_51),
.B(n_2),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_81),
.B(n_64),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_30),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_65),
.B(n_63),
.C(n_66),
.D(n_12),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_1),
.C(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_81),
.B1(n_66),
.B2(n_82),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_80),
.C(n_69),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_63),
.B(n_3),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_3),
.B(n_5),
.C(n_7),
.D(n_10),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_60),
.B1(n_15),
.B2(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_84),
.B1(n_40),
.B2(n_88),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_97),
.B(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_93),
.C(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_26),
.C(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_96),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_53),
.C(n_40),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_5),
.B(n_7),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.C(n_104),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_52),
.Y(n_110)
);


endmodule