module real_aes_15767_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_16;
wire n_13;
wire n_15;
wire n_7;
wire n_9;
wire n_8;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
AOI221xp5_ASAP7_75t_R g6 ( .A1(n_0), .A2(n_5), .B1(n_7), .B2(n_9), .C(n_11), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g7 ( .A(n_2), .B(n_8), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_2), .B(n_3), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_2), .B(n_3), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_3), .Y(n_8) );
NOR2xp33_ASAP7_75t_R g9 ( .A(n_3), .B(n_10), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
OAI22xp33_ASAP7_75t_SL g11 ( .A1(n_12), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
endmodule