module fake_aes_695_n_1666 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_296, n_157, n_79, n_202, n_386, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_389, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_387, n_163, n_105, n_227, n_384, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_381, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_388, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_385, n_257, n_269, n_1666);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_386;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_389;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_387;
input n_163;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_381;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_388;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1666;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_1663;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_1657;
wire n_1655;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_659;
wire n_432;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1659;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVxp67_ASAP7_75t_L g390 ( .A(n_108), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_222), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_163), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_29), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_180), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_123), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_78), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_89), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_383), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_388), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_317), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_203), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_121), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_274), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_199), .Y(n_405) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_284), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_55), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_362), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_19), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_27), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_147), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_7), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_47), .Y(n_413) );
BUFx10_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_204), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_280), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_218), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_141), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_257), .Y(n_419) );
NOR2xp67_ASAP7_75t_L g420 ( .A(n_71), .B(n_304), .Y(n_420) );
BUFx5_ASAP7_75t_L g421 ( .A(n_118), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_282), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_35), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_26), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_39), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_344), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_50), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_119), .Y(n_428) );
INVx4_ASAP7_75t_R g429 ( .A(n_197), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_272), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_34), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_45), .B(n_333), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_104), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_50), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_379), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_135), .Y(n_436) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_318), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_0), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_101), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_21), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_309), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_226), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_292), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_370), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_360), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_366), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_386), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_42), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_352), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_0), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_99), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_252), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_269), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_316), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_266), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_117), .B(n_42), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_163), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_189), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g459 ( .A(n_192), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_220), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_112), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_140), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_212), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_129), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_251), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_70), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_306), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_55), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_160), .B(n_334), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_57), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_261), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_51), .Y(n_472) );
INVxp33_ASAP7_75t_L g473 ( .A(n_169), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_53), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_250), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_198), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_1), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_363), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_15), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_187), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_215), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_26), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_353), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_384), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_123), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_299), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_287), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_14), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_361), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_20), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_234), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_270), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_305), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_96), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_313), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_247), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_164), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_225), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_98), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_6), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_111), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_324), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_389), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_185), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_256), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_210), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_275), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_268), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_186), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_346), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_327), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_188), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_291), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_36), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_254), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_8), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_314), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_321), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_358), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_349), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_57), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_331), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_147), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_378), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_48), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_43), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_140), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_281), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_224), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_355), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_53), .Y(n_531) );
INVxp33_ASAP7_75t_L g532 ( .A(n_308), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_124), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_206), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_136), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_223), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_246), .Y(n_537) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_143), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_76), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_289), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_312), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_155), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_82), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_99), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_330), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_193), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_75), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_211), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_89), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_66), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_86), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_301), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_377), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_102), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_342), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_190), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_77), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_58), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_153), .B(n_255), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_267), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_124), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_347), .Y(n_562) );
INVxp33_ASAP7_75t_L g563 ( .A(n_191), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_231), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_92), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_61), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_260), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_87), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_290), .Y(n_569) );
BUFx3_ASAP7_75t_L g570 ( .A(n_241), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_86), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_178), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_70), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_43), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_387), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_235), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_21), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g578 ( .A(n_90), .Y(n_578) );
CKINVDCx14_ASAP7_75t_R g579 ( .A(n_213), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_67), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_72), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_340), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_264), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_296), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_357), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_183), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_136), .Y(n_587) );
BUFx3_ASAP7_75t_L g588 ( .A(n_121), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_35), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_295), .Y(n_590) );
INVx5_ASAP7_75t_L g591 ( .A(n_402), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_558), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g593 ( .A1(n_411), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_402), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_413), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_402), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_558), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_479), .B(n_4), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_566), .B(n_5), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_558), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_402), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_473), .B(n_5), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_421), .Y(n_603) );
INVx6_ASAP7_75t_L g604 ( .A(n_414), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_421), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_473), .B(n_6), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_421), .Y(n_607) );
OA21x2_ASAP7_75t_L g608 ( .A1(n_415), .A2(n_173), .B(n_172), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_421), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_421), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_455), .B(n_8), .Y(n_611) );
INVxp33_ASAP7_75t_SL g612 ( .A(n_410), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_421), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_486), .B(n_9), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_562), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_414), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_421), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_578), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_589), .Y(n_621) );
OAI22xp5_ASAP7_75t_SL g622 ( .A1(n_411), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_525), .B(n_12), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_393), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g625 ( .A1(n_485), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_532), .B(n_13), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_414), .B(n_582), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_582), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_393), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_543), .B(n_16), .Y(n_630) );
CKINVDCx6p67_ASAP7_75t_R g631 ( .A(n_446), .Y(n_631) );
AND2x6_ASAP7_75t_L g632 ( .A(n_623), .B(n_517), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_617), .B(n_525), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_603), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_603), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_605), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_605), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_607), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_620), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_617), .B(n_532), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_607), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
OR2x6_ASAP7_75t_L g643 ( .A(n_593), .B(n_456), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_593), .B(n_433), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_623), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_604), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_602), .A2(n_396), .B1(n_398), .B2(n_397), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_609), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_631), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_610), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_621), .Y(n_651) );
INVx6_ASAP7_75t_L g652 ( .A(n_604), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_604), .B(n_563), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_610), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_617), .B(n_453), .Y(n_655) );
CKINVDCx6p67_ASAP7_75t_R g656 ( .A(n_631), .Y(n_656) );
INVx5_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_614), .Y(n_658) );
OAI22xp33_ASAP7_75t_SL g659 ( .A1(n_619), .A2(n_440), .B1(n_501), .B2(n_418), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_618), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_618), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_592), .Y(n_663) );
BUFx3_ASAP7_75t_L g664 ( .A(n_604), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_621), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_617), .B(n_563), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_592), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_597), .Y(n_668) );
INVx4_ASAP7_75t_L g669 ( .A(n_623), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_602), .A2(n_403), .B1(n_409), .B2(n_407), .Y(n_670) );
INVx8_ASAP7_75t_L g671 ( .A(n_632), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_663), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_640), .B(n_626), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_633), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_651), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_666), .B(n_606), .Y(n_676) );
NOR2x1p5_ASAP7_75t_L g677 ( .A(n_656), .B(n_615), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_633), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_655), .B(n_606), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_633), .Y(n_680) );
NAND2x1_ASAP7_75t_L g681 ( .A(n_645), .B(n_429), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_667), .A2(n_623), .B(n_600), .C(n_597), .Y(n_682) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_665), .B(n_619), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_645), .B(n_612), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_653), .B(n_627), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_649), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_669), .B(n_635), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_667), .A2(n_600), .B(n_611), .C(n_599), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_633), .B(n_615), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_669), .B(n_506), .Y(n_690) );
AOI21x1_ASAP7_75t_L g691 ( .A1(n_635), .A2(n_608), .B(n_599), .Y(n_691) );
INVx6_ASAP7_75t_L g692 ( .A(n_652), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_668), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_632), .A2(n_629), .B1(n_624), .B2(n_412), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_668), .A2(n_598), .B(n_630), .C(n_629), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_634), .Y(n_696) );
AND2x4_ASAP7_75t_SL g697 ( .A(n_656), .B(n_430), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_652), .Y(n_698) );
BUFx3_ASAP7_75t_L g699 ( .A(n_632), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_634), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_637), .A2(n_598), .B(n_624), .C(n_588), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_632), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_652), .B(n_510), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_652), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_632), .B(n_417), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_632), .B(n_419), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_636), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_636), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_641), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_632), .Y(n_710) );
INVxp67_ASAP7_75t_L g711 ( .A(n_646), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_641), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_664), .B(n_419), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_664), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_647), .B(n_454), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_670), .B(n_454), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_638), .B(n_642), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_643), .A2(n_424), .B1(n_427), .B2(n_425), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_638), .B(n_524), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_648), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_642), .B(n_524), .Y(n_721) );
INVx4_ASAP7_75t_L g722 ( .A(n_648), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_650), .B(n_540), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_662), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_650), .B(n_540), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_654), .B(n_546), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_654), .Y(n_727) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_657), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_658), .B(n_546), .Y(n_729) );
AND2x6_ASAP7_75t_SL g730 ( .A(n_644), .B(n_622), .Y(n_730) );
NAND2xp33_ASAP7_75t_L g731 ( .A(n_658), .B(n_548), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_644), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_660), .B(n_391), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_660), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_661), .B(n_394), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_661), .B(n_548), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_662), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_659), .B(n_406), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_657), .B(n_564), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_657), .B(n_564), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_657), .B(n_590), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_643), .B(n_430), .Y(n_742) );
BUFx4_ASAP7_75t_L g743 ( .A(n_644), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_657), .B(n_395), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_643), .B(n_437), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_643), .B(n_437), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_644), .B(n_595), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_673), .B(n_418), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_676), .B(n_440), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_710), .B(n_406), .Y(n_750) );
NOR2xp67_ASAP7_75t_SL g751 ( .A(n_710), .B(n_501), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_L g752 ( .A1(n_695), .A2(n_688), .B(n_701), .C(n_682), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_689), .B(n_527), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_710), .B(n_435), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_694), .A2(n_435), .B1(n_447), .B2(n_443), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_687), .A2(n_608), .B(n_432), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_675), .Y(n_757) );
AO32x2_ASAP7_75t_L g758 ( .A1(n_698), .A2(n_622), .A3(n_625), .B1(n_595), .B2(n_608), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_674), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_678), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_710), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_679), .B(n_527), .Y(n_762) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_671), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_687), .A2(n_608), .B(n_536), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_679), .B(n_531), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_722), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_680), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_693), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_684), .B(n_644), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_699), .B(n_443), .Y(n_770) );
BUFx4f_ASAP7_75t_L g771 ( .A(n_697), .Y(n_771) );
OR2x6_ASAP7_75t_L g772 ( .A(n_686), .B(n_625), .Y(n_772) );
OR2x6_ASAP7_75t_L g773 ( .A(n_677), .B(n_390), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_743), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_722), .B(n_547), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_742), .Y(n_776) );
OR2x6_ASAP7_75t_L g777 ( .A(n_742), .B(n_461), .Y(n_777) );
CKINVDCx11_ASAP7_75t_R g778 ( .A(n_730), .Y(n_778) );
BUFx3_ASAP7_75t_L g779 ( .A(n_692), .Y(n_779) );
OR2x6_ASAP7_75t_SL g780 ( .A(n_747), .B(n_547), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_699), .B(n_447), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_734), .Y(n_782) );
BUFx12f_ASAP7_75t_L g783 ( .A(n_702), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_734), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_717), .A2(n_404), .B(n_401), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_690), .B(n_549), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_683), .B(n_485), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_719), .B(n_549), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_738), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_732), .B(n_523), .C(n_450), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_694), .A2(n_475), .B1(n_522), .B2(n_496), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_671), .A2(n_475), .B1(n_522), .B2(n_496), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_724), .B(n_537), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_716), .B(n_537), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_723), .B(n_550), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_L g796 ( .A1(n_715), .A2(n_538), .B(n_436), .C(n_438), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_717), .A2(n_408), .B(n_405), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_725), .B(n_550), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_685), .A2(n_588), .B(n_577), .C(n_431), .Y(n_799) );
INVx5_ASAP7_75t_L g800 ( .A(n_671), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_724), .A2(n_576), .B1(n_579), .B2(n_459), .Y(n_801) );
O2A1O1Ixp5_ASAP7_75t_L g802 ( .A1(n_685), .A2(n_559), .B(n_416), .C(n_422), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_728), .Y(n_803) );
OR2x6_ASAP7_75t_SL g804 ( .A(n_745), .B(n_392), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_736), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_672), .Y(n_806) );
NAND2x1p5_ASAP7_75t_L g807 ( .A(n_727), .B(n_516), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_727), .B(n_576), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_737), .B(n_423), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g810 ( .A(n_705), .B(n_399), .Y(n_810) );
O2A1O1Ixp5_ASAP7_75t_L g811 ( .A1(n_691), .A2(n_415), .B(n_422), .C(n_416), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_706), .A2(n_442), .B(n_441), .Y(n_812) );
BUFx12f_ASAP7_75t_L g813 ( .A(n_728), .Y(n_813) );
AND2x6_ASAP7_75t_L g814 ( .A(n_714), .B(n_517), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_696), .A2(n_445), .B(n_444), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_700), .A2(n_452), .B(n_449), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_700), .A2(n_465), .B(n_463), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_713), .Y(n_818) );
INVx1_ASAP7_75t_SL g819 ( .A(n_739), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_746), .B(n_428), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_733), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_731), .B(n_439), .Y(n_822) );
NAND2x1p5_ASAP7_75t_L g823 ( .A(n_714), .B(n_544), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_738), .A2(n_468), .B1(n_494), .B2(n_464), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_718), .B(n_568), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_733), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_718), .A2(n_459), .B1(n_579), .B2(n_469), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_721), .B(n_726), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_703), .B(n_497), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_703), .B(n_499), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_735), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_681), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_707), .A2(n_462), .B1(n_466), .B2(n_448), .Y(n_833) );
INVx5_ASAP7_75t_L g834 ( .A(n_728), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_708), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_709), .A2(n_482), .B1(n_490), .B2(n_477), .Y(n_836) );
NOR2xp33_ASAP7_75t_R g837 ( .A(n_704), .B(n_580), .Y(n_837) );
AO32x2_ASAP7_75t_L g838 ( .A1(n_735), .A2(n_420), .A3(n_628), .B1(n_620), .B2(n_582), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_712), .A2(n_471), .B(n_467), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_729), .Y(n_840) );
OAI21xp33_ASAP7_75t_L g841 ( .A1(n_712), .A2(n_581), .B(n_514), .Y(n_841) );
OAI21xp33_ASAP7_75t_SL g842 ( .A1(n_720), .A2(n_521), .B(n_500), .Y(n_842) );
A2O1A1Ixp33_ASAP7_75t_L g843 ( .A1(n_720), .A2(n_533), .B(n_535), .C(n_526), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_L g844 ( .A1(n_711), .A2(n_542), .B(n_551), .C(n_539), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_728), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g846 ( .A(n_741), .B(n_400), .Y(n_846) );
INVx4_ASAP7_75t_L g847 ( .A(n_692), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_740), .B(n_557), .Y(n_848) );
OAI22xp5_ASAP7_75t_SL g849 ( .A1(n_692), .A2(n_565), .B1(n_573), .B2(n_561), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_744), .B(n_574), .Y(n_850) );
A2O1A1Ixp33_ASAP7_75t_SL g851 ( .A1(n_744), .A2(n_594), .B(n_601), .C(n_596), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_683), .A2(n_587), .B1(n_478), .B2(n_480), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_687), .A2(n_481), .B(n_476), .Y(n_853) );
A2O1A1Ixp33_ASAP7_75t_L g854 ( .A1(n_717), .A2(n_433), .B(n_451), .C(n_434), .Y(n_854) );
O2A1O1Ixp33_ASAP7_75t_L g855 ( .A1(n_695), .A2(n_434), .B(n_457), .C(n_451), .Y(n_855) );
O2A1O1Ixp33_ASAP7_75t_L g856 ( .A1(n_695), .A2(n_457), .B(n_472), .C(n_470), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_722), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_674), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_674), .Y(n_859) );
AOI21x1_ASAP7_75t_L g860 ( .A1(n_691), .A2(n_487), .B(n_484), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_722), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_687), .A2(n_493), .B(n_491), .Y(n_862) );
OR2x6_ASAP7_75t_L g863 ( .A(n_686), .B(n_470), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_717), .A2(n_472), .B(n_554), .C(n_488), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_687), .A2(n_498), .B(n_495), .Y(n_865) );
AOI221xp5_ASAP7_75t_SL g866 ( .A1(n_695), .A2(n_488), .B1(n_571), .B2(n_554), .C(n_545), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_683), .A2(n_503), .B1(n_504), .B2(n_502), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g868 ( .A1(n_717), .A2(n_508), .B(n_507), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_674), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_693), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_755), .A2(n_571), .B1(n_474), .B2(n_458), .Y(n_871) );
INVx4_ASAP7_75t_L g872 ( .A(n_813), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_782), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_768), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_757), .B(n_474), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_771), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_807), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_870), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_787), .B(n_426), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_SL g880 ( .A1(n_799), .A2(n_513), .B(n_518), .C(n_512), .Y(n_880) );
A2O1A1Ixp33_ASAP7_75t_L g881 ( .A1(n_752), .A2(n_520), .B(n_528), .C(n_519), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_823), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_870), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_834), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_759), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_771), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_760), .Y(n_887) );
AND2x4_ASAP7_75t_L g888 ( .A(n_800), .B(n_541), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_767), .Y(n_889) );
INVx5_ASAP7_75t_L g890 ( .A(n_834), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_784), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_756), .A2(n_553), .B(n_552), .Y(n_892) );
INVxp67_ASAP7_75t_L g893 ( .A(n_863), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_764), .A2(n_560), .B(n_555), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_778), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_835), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_L g897 ( .A1(n_855), .A2(n_856), .B(n_802), .C(n_812), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_777), .A2(n_474), .B1(n_572), .B2(n_567), .Y(n_898) );
AOI31xp67_ASAP7_75t_L g899 ( .A1(n_845), .A2(n_596), .A3(n_601), .B(n_594), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_769), .B(n_474), .Y(n_900) );
O2A1O1Ixp33_ASAP7_75t_L g901 ( .A1(n_854), .A2(n_585), .B(n_583), .C(n_530), .Y(n_901) );
NAND2x1p5_ASAP7_75t_L g902 ( .A(n_834), .B(n_556), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_806), .A2(n_530), .B(n_529), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_777), .B(n_505), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_791), .A2(n_483), .B1(n_489), .B2(n_460), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_766), .Y(n_906) );
INVx5_ASAP7_75t_L g907 ( .A(n_814), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_805), .B(n_492), .Y(n_908) );
AND2x2_ASAP7_75t_SL g909 ( .A(n_792), .B(n_529), .Y(n_909) );
CKINVDCx11_ASAP7_75t_R g910 ( .A(n_774), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_780), .B(n_16), .Y(n_911) );
A2O1A1Ixp33_ASAP7_75t_L g912 ( .A1(n_785), .A2(n_569), .B(n_584), .C(n_534), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_809), .A2(n_569), .B(n_534), .Y(n_913) );
A2O1A1Ixp33_ASAP7_75t_L g914 ( .A1(n_797), .A2(n_584), .B(n_570), .C(n_556), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_857), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_825), .B(n_515), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_827), .A2(n_794), .B1(n_801), .B2(n_868), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_858), .Y(n_918) );
AO32x2_ASAP7_75t_L g919 ( .A1(n_833), .A2(n_628), .A3(n_620), .B1(n_594), .B2(n_613), .Y(n_919) );
AO31x2_ASAP7_75t_L g920 ( .A1(n_864), .A2(n_601), .A3(n_613), .B(n_596), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_859), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_863), .B(n_17), .Y(n_922) );
AOI21xp5_ASAP7_75t_L g923 ( .A1(n_821), .A2(n_511), .B(n_509), .Y(n_923) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_803), .Y(n_924) );
O2A1O1Ixp33_ASAP7_75t_SL g925 ( .A1(n_851), .A2(n_575), .B(n_616), .C(n_613), .Y(n_925) );
BUFx2_ASAP7_75t_L g926 ( .A(n_837), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_793), .A2(n_586), .B1(n_570), .B2(n_582), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_789), .B(n_18), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_779), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_844), .A2(n_628), .B1(n_620), .B2(n_591), .C(n_639), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_772), .B(n_18), .Y(n_931) );
INVx1_ASAP7_75t_SL g932 ( .A(n_808), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_869), .Y(n_933) );
AOI21xp5_ASAP7_75t_L g934 ( .A1(n_826), .A2(n_639), .B(n_591), .Y(n_934) );
OAI21x1_ASAP7_75t_L g935 ( .A1(n_815), .A2(n_628), .B(n_175), .Y(n_935) );
OAI21x1_ASAP7_75t_L g936 ( .A1(n_816), .A2(n_628), .B(n_176), .Y(n_936) );
A2O1A1Ixp33_ASAP7_75t_L g937 ( .A1(n_866), .A2(n_591), .B(n_639), .C(n_22), .Y(n_937) );
O2A1O1Ixp33_ASAP7_75t_L g938 ( .A1(n_843), .A2(n_22), .B(n_19), .C(n_20), .Y(n_938) );
BUFx4f_ASAP7_75t_SL g939 ( .A(n_783), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_861), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_776), .A2(n_591), .B1(n_639), .B2(n_25), .Y(n_941) );
A2O1A1Ixp33_ASAP7_75t_L g942 ( .A1(n_796), .A2(n_591), .B(n_639), .C(n_27), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_831), .Y(n_943) );
AND2x4_ASAP7_75t_L g944 ( .A(n_800), .B(n_23), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_842), .A2(n_29), .B(n_24), .C(n_28), .Y(n_945) );
AO21x2_ASAP7_75t_L g946 ( .A1(n_817), .A2(n_177), .B(n_174), .Y(n_946) );
INVx4_ASAP7_75t_SL g947 ( .A(n_814), .Y(n_947) );
AO31x2_ASAP7_75t_L g948 ( .A1(n_839), .A2(n_31), .A3(n_24), .B(n_30), .Y(n_948) );
BUFx2_ASAP7_75t_R g949 ( .A(n_804), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_850), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_775), .Y(n_951) );
AO31x2_ASAP7_75t_L g952 ( .A1(n_836), .A2(n_32), .A3(n_30), .B(n_31), .Y(n_952) );
INVx4_ASAP7_75t_L g953 ( .A(n_800), .Y(n_953) );
OAI21x1_ASAP7_75t_L g954 ( .A1(n_853), .A2(n_181), .B(n_179), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_788), .A2(n_184), .B(n_182), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_830), .B(n_32), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_848), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_803), .Y(n_958) );
CKINVDCx11_ASAP7_75t_R g959 ( .A(n_773), .Y(n_959) );
INVx6_ASAP7_75t_L g960 ( .A(n_773), .Y(n_960) );
BUFx2_ASAP7_75t_R g961 ( .A(n_770), .Y(n_961) );
O2A1O1Ixp5_ASAP7_75t_L g962 ( .A1(n_750), .A2(n_195), .B(n_196), .C(n_194), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_849), .A2(n_36), .B1(n_33), .B2(n_34), .Y(n_963) );
O2A1O1Ixp33_ASAP7_75t_L g964 ( .A1(n_786), .A2(n_38), .B(n_33), .C(n_37), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_852), .B(n_37), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g966 ( .A1(n_790), .A2(n_40), .B1(n_38), .B2(n_39), .Y(n_966) );
NOR3xp33_ASAP7_75t_L g967 ( .A(n_829), .B(n_40), .C(n_41), .Y(n_967) );
INVx2_ASAP7_75t_SL g968 ( .A(n_828), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_762), .B(n_41), .Y(n_969) );
AO31x2_ASAP7_75t_L g970 ( .A1(n_862), .A2(n_46), .A3(n_44), .B(n_45), .Y(n_970) );
AO31x2_ASAP7_75t_L g971 ( .A1(n_865), .A2(n_47), .A3(n_44), .B(n_46), .Y(n_971) );
INVx6_ASAP7_75t_L g972 ( .A(n_847), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_765), .A2(n_51), .B1(n_48), .B2(n_49), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_803), .Y(n_974) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_867), .A2(n_54), .B(n_49), .C(n_52), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_758), .Y(n_976) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_761), .Y(n_977) );
OAI22xp5_ASAP7_75t_SL g978 ( .A1(n_840), .A2(n_56), .B1(n_52), .B2(n_54), .Y(n_978) );
O2A1O1Ixp33_ASAP7_75t_L g979 ( .A1(n_748), .A2(n_59), .B(n_56), .C(n_58), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_824), .B(n_59), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_749), .B(n_60), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_758), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g983 ( .A(n_818), .Y(n_983) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_761), .Y(n_984) );
BUFx3_ASAP7_75t_L g985 ( .A(n_832), .Y(n_985) );
AO32x2_ASAP7_75t_L g986 ( .A1(n_838), .A2(n_60), .A3(n_61), .B1(n_62), .B2(n_63), .Y(n_986) );
O2A1O1Ixp33_ASAP7_75t_L g987 ( .A1(n_795), .A2(n_64), .B(n_62), .C(n_63), .Y(n_987) );
BUFx8_ASAP7_75t_L g988 ( .A(n_758), .Y(n_988) );
AO32x2_ASAP7_75t_L g989 ( .A1(n_838), .A2(n_64), .A3(n_65), .B1(n_66), .B2(n_67), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_753), .Y(n_990) );
A2O1A1Ixp33_ASAP7_75t_L g991 ( .A1(n_820), .A2(n_69), .B(n_65), .C(n_68), .Y(n_991) );
AOI21xp5_ASAP7_75t_L g992 ( .A1(n_798), .A2(n_201), .B(n_200), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g993 ( .A1(n_841), .A2(n_71), .B(n_68), .C(n_69), .Y(n_993) );
AOI21xp5_ASAP7_75t_L g994 ( .A1(n_810), .A2(n_205), .B(n_202), .Y(n_994) );
OAI21xp5_ASAP7_75t_L g995 ( .A1(n_819), .A2(n_208), .B(n_207), .Y(n_995) );
INVx2_ASAP7_75t_SL g996 ( .A(n_828), .Y(n_996) );
BUFx2_ASAP7_75t_R g997 ( .A(n_781), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g998 ( .A1(n_846), .A2(n_214), .B(n_209), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_754), .B(n_72), .Y(n_999) );
OAI21x1_ASAP7_75t_L g1000 ( .A1(n_822), .A2(n_217), .B(n_216), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_761), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_847), .Y(n_1002) );
OR2x6_ASAP7_75t_L g1003 ( .A(n_763), .B(n_73), .Y(n_1003) );
A2O1A1Ixp33_ASAP7_75t_L g1004 ( .A1(n_751), .A2(n_75), .B(n_73), .C(n_74), .Y(n_1004) );
AOI21xp5_ASAP7_75t_L g1005 ( .A1(n_763), .A2(n_221), .B(n_219), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_763), .Y(n_1006) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_814), .B(n_74), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_769), .B(n_76), .Y(n_1008) );
BUFx2_ASAP7_75t_SL g1009 ( .A(n_834), .Y(n_1009) );
O2A1O1Ixp33_ASAP7_75t_SL g1010 ( .A1(n_799), .A2(n_228), .B(n_229), .C(n_227), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_756), .A2(n_232), .B(n_230), .Y(n_1011) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_811), .A2(n_236), .B(n_233), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_769), .B(n_77), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_782), .Y(n_1014) );
INVx2_ASAP7_75t_L g1015 ( .A(n_782), .Y(n_1015) );
O2A1O1Ixp33_ASAP7_75t_L g1016 ( .A1(n_799), .A2(n_78), .B(n_79), .C(n_80), .Y(n_1016) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_756), .A2(n_238), .B(n_237), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_756), .A2(n_240), .B(n_239), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_768), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_755), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_787), .B(n_81), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_769), .B(n_82), .Y(n_1022) );
INVx2_ASAP7_75t_L g1023 ( .A(n_782), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_787), .B(n_83), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g1025 ( .A1(n_756), .A2(n_243), .B(n_242), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_755), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1026) );
OAI21x1_ASAP7_75t_L g1027 ( .A1(n_860), .A2(n_245), .B(n_244), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_874), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_890), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_947), .B(n_84), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g1031 ( .A1(n_892), .A2(n_249), .B(n_248), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1019), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_878), .Y(n_1033) );
AO31x2_ASAP7_75t_L g1034 ( .A1(n_976), .A2(n_85), .A3(n_87), .B(n_88), .Y(n_1034) );
INVxp67_ASAP7_75t_SL g1035 ( .A(n_1006), .Y(n_1035) );
A2O1A1Ixp33_ASAP7_75t_L g1036 ( .A1(n_1021), .A2(n_88), .B(n_90), .C(n_91), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_885), .Y(n_1037) );
AO21x2_ASAP7_75t_L g1038 ( .A1(n_1012), .A2(n_258), .B(n_253), .Y(n_1038) );
OAI21xp5_ASAP7_75t_L g1039 ( .A1(n_897), .A2(n_93), .B(n_94), .Y(n_1039) );
INVx3_ASAP7_75t_L g1040 ( .A(n_890), .Y(n_1040) );
A2O1A1Ixp33_ASAP7_75t_L g1041 ( .A1(n_1024), .A2(n_917), .B(n_1016), .C(n_901), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_887), .Y(n_1042) );
NOR2xp33_ASAP7_75t_SL g1043 ( .A(n_907), .B(n_93), .Y(n_1043) );
AOI21xp5_ASAP7_75t_L g1044 ( .A1(n_894), .A2(n_262), .B(n_259), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_988), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_883), .Y(n_1046) );
AO31x2_ASAP7_75t_L g1047 ( .A1(n_982), .A2(n_95), .A3(n_97), .B(n_98), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_909), .B(n_97), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_877), .B(n_100), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_988), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_889), .Y(n_1051) );
AOI21xp5_ASAP7_75t_L g1052 ( .A1(n_925), .A2(n_265), .B(n_263), .Y(n_1052) );
OAI221xp5_ASAP7_75t_SL g1053 ( .A1(n_911), .A2(n_103), .B1(n_104), .B2(n_105), .C(n_106), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_918), .Y(n_1054) );
A2O1A1Ixp33_ASAP7_75t_L g1055 ( .A1(n_969), .A2(n_103), .B(n_105), .C(n_106), .Y(n_1055) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_872), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g1057 ( .A(n_890), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_1003), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_990), .B(n_107), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_980), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1061 ( .A1(n_898), .A2(n_110), .B1(n_112), .B2(n_113), .C(n_114), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_921), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_933), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_1011), .A2(n_273), .B(n_271), .Y(n_1064) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_959), .Y(n_1065) );
INVx4_ASAP7_75t_L g1066 ( .A(n_872), .Y(n_1066) );
OAI22x1_ASAP7_75t_L g1067 ( .A1(n_926), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_873), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_891), .Y(n_1069) );
OA21x2_ASAP7_75t_L g1070 ( .A1(n_1027), .A2(n_277), .B(n_276), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_983), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1014), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_957), .B(n_115), .Y(n_1073) );
AO21x2_ASAP7_75t_L g1074 ( .A1(n_937), .A2(n_294), .B(n_385), .Y(n_1074) );
AO21x2_ASAP7_75t_L g1075 ( .A1(n_900), .A2(n_293), .B(n_382), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_947), .B(n_116), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_922), .B(n_116), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1015), .Y(n_1078) );
AO21x2_ASAP7_75t_L g1079 ( .A1(n_1017), .A2(n_297), .B(n_381), .Y(n_1079) );
OAI21xp5_ASAP7_75t_L g1080 ( .A1(n_881), .A2(n_117), .B(n_118), .Y(n_1080) );
CKINVDCx11_ASAP7_75t_R g1081 ( .A(n_910), .Y(n_1081) );
AO21x2_ASAP7_75t_L g1082 ( .A1(n_1018), .A2(n_298), .B(n_380), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1003), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_960), .B(n_119), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_951), .B(n_120), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_950), .B(n_120), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_950), .B(n_122), .Y(n_1087) );
OA21x2_ASAP7_75t_L g1088 ( .A1(n_935), .A2(n_300), .B(n_376), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_956), .B(n_125), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_943), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1023), .B(n_125), .Y(n_1091) );
OR2x6_ASAP7_75t_L g1092 ( .A(n_1009), .B(n_126), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_875), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_882), .Y(n_1094) );
AOI21xp5_ASAP7_75t_L g1095 ( .A1(n_1025), .A2(n_303), .B(n_375), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_896), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g1097 ( .A1(n_942), .A2(n_127), .B(n_128), .Y(n_1097) );
OR2x6_ASAP7_75t_L g1098 ( .A(n_960), .B(n_130), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_907), .B(n_130), .Y(n_1099) );
OR2x6_ASAP7_75t_L g1100 ( .A(n_1007), .B(n_131), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_1007), .Y(n_1101) );
OA21x2_ASAP7_75t_L g1102 ( .A1(n_936), .A2(n_307), .B(n_374), .Y(n_1102) );
AOI21xp5_ASAP7_75t_L g1103 ( .A1(n_934), .A2(n_302), .B(n_373), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_978), .A2(n_131), .B1(n_132), .B2(n_133), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_1020), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_906), .Y(n_1106) );
OR2x6_ASAP7_75t_L g1107 ( .A(n_944), .B(n_134), .Y(n_1107) );
OAI21x1_ASAP7_75t_L g1108 ( .A1(n_1000), .A2(n_311), .B(n_369), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_915), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_970), .Y(n_1110) );
OA21x2_ASAP7_75t_L g1111 ( .A1(n_954), .A2(n_310), .B(n_368), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_931), .B(n_135), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_968), .B(n_137), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_932), .B(n_137), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_928), .A2(n_138), .B1(n_139), .B2(n_141), .Y(n_1115) );
INVxp67_ASAP7_75t_L g1116 ( .A(n_949), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_1010), .A2(n_913), .B(n_981), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_996), .B(n_138), .Y(n_1118) );
AO31x2_ASAP7_75t_L g1119 ( .A1(n_914), .A2(n_139), .A3(n_142), .B(n_143), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_940), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_880), .A2(n_319), .B(n_367), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_893), .B(n_142), .Y(n_1122) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_955), .A2(n_320), .B(n_365), .Y(n_1123) );
A2O1A1Ixp33_ASAP7_75t_L g1124 ( .A1(n_987), .A2(n_144), .B(n_145), .C(n_146), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_879), .B(n_144), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_967), .A2(n_145), .B1(n_146), .B2(n_148), .Y(n_1126) );
OAI21xp5_ASAP7_75t_L g1127 ( .A1(n_912), .A2(n_148), .B(n_149), .Y(n_1127) );
AOI21xp33_ASAP7_75t_L g1128 ( .A1(n_1008), .A2(n_149), .B(n_150), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1013), .B(n_150), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_992), .A2(n_325), .B(n_364), .Y(n_1130) );
A2O1A1Ixp33_ASAP7_75t_L g1131 ( .A1(n_964), .A2(n_151), .B(n_152), .C(n_153), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_999), .A2(n_151), .B1(n_152), .B2(n_154), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_920), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1134 ( .A(n_939), .Y(n_1134) );
NAND2xp5_ASAP7_75t_SL g1135 ( .A(n_907), .B(n_154), .Y(n_1135) );
AO31x2_ASAP7_75t_L g1136 ( .A1(n_993), .A2(n_155), .A3(n_156), .B(n_157), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_899), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1138 ( .A1(n_1026), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_1138) );
AOI21xp5_ASAP7_75t_L g1139 ( .A1(n_1001), .A2(n_326), .B(n_359), .Y(n_1139) );
AOI21xp5_ASAP7_75t_L g1140 ( .A1(n_1001), .A2(n_323), .B(n_356), .Y(n_1140) );
AOI21x1_ASAP7_75t_L g1141 ( .A1(n_903), .A2(n_322), .B(n_354), .Y(n_1141) );
AO31x2_ASAP7_75t_L g1142 ( .A1(n_1004), .A2(n_158), .A3(n_159), .B(n_160), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_970), .Y(n_1143) );
AOI21xp5_ASAP7_75t_L g1144 ( .A1(n_984), .A2(n_328), .B(n_351), .Y(n_1144) );
CKINVDCx11_ASAP7_75t_R g1145 ( .A(n_929), .Y(n_1145) );
AO31x2_ASAP7_75t_L g1146 ( .A1(n_945), .A2(n_159), .A3(n_161), .B(n_162), .Y(n_1146) );
INVx3_ASAP7_75t_L g1147 ( .A(n_953), .Y(n_1147) );
OAI22xp33_ASAP7_75t_SL g1148 ( .A1(n_966), .A2(n_161), .B1(n_162), .B2(n_164), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_971), .Y(n_1149) );
INVxp33_ASAP7_75t_L g1150 ( .A(n_904), .Y(n_1150) );
AOI21xp5_ASAP7_75t_L g1151 ( .A1(n_1022), .A2(n_329), .B(n_350), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_971), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_871), .A2(n_165), .B1(n_166), .B2(n_167), .C(n_168), .Y(n_1153) );
OA21x2_ASAP7_75t_L g1154 ( .A1(n_995), .A2(n_962), .B(n_994), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_944), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_965), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_952), .Y(n_1157) );
OAI21x1_ASAP7_75t_L g1158 ( .A1(n_958), .A2(n_335), .B(n_348), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_916), .B(n_170), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_952), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_908), .B(n_171), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_938), .A2(n_171), .B1(n_278), .B2(n_279), .C(n_283), .Y(n_1162) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_953), .B(n_285), .Y(n_1163) );
OA21x2_ASAP7_75t_L g1164 ( .A1(n_998), .A2(n_286), .B(n_288), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1165 ( .A(n_876), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_948), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_952), .Y(n_1167) );
OAI21xp33_ASAP7_75t_SL g1168 ( .A1(n_973), .A2(n_315), .B(n_332), .Y(n_1168) );
OAI22x1_ASAP7_75t_L g1169 ( .A1(n_886), .A2(n_336), .B1(n_337), .B2(n_338), .Y(n_1169) );
INVx3_ASAP7_75t_SL g1170 ( .A(n_895), .Y(n_1170) );
NAND2x1p5_ASAP7_75t_L g1171 ( .A(n_884), .B(n_339), .Y(n_1171) );
A2O1A1Ixp33_ASAP7_75t_L g1172 ( .A1(n_979), .A2(n_341), .B(n_343), .C(n_345), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_961), .B(n_997), .Y(n_1173) );
OAI21x1_ASAP7_75t_SL g1174 ( .A1(n_974), .A2(n_1005), .B(n_923), .Y(n_1174) );
AOI21xp5_ASAP7_75t_L g1175 ( .A1(n_946), .A2(n_977), .B(n_924), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_905), .B(n_884), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_888), .A2(n_963), .B1(n_930), .B2(n_1002), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_888), .B(n_985), .Y(n_1178) );
OAI22xp33_ASAP7_75t_L g1179 ( .A1(n_927), .A2(n_941), .B1(n_902), .B2(n_972), .Y(n_1179) );
OA21x2_ASAP7_75t_L g1180 ( .A1(n_991), .A2(n_975), .B(n_919), .Y(n_1180) );
OA21x2_ASAP7_75t_L g1181 ( .A1(n_919), .A2(n_986), .B(n_989), .Y(n_1181) );
AOI21xp5_ASAP7_75t_L g1182 ( .A1(n_977), .A2(n_924), .B(n_919), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_972), .Y(n_1183) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_1057), .Y(n_1184) );
BUFx6f_ASAP7_75t_L g1185 ( .A(n_1057), .Y(n_1185) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1137), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1056), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1028), .Y(n_1188) );
BUFx3_ASAP7_75t_L g1189 ( .A(n_1057), .Y(n_1189) );
AO21x2_ASAP7_75t_L g1190 ( .A1(n_1157), .A2(n_986), .B(n_989), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1032), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1107), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1037), .B(n_948), .Y(n_1193) );
NOR2x1_ASAP7_75t_R g1194 ( .A(n_1081), .B(n_924), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1042), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1051), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1054), .Y(n_1197) );
OAI21xp5_ASAP7_75t_L g1198 ( .A1(n_1041), .A2(n_986), .B(n_989), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1068), .B(n_977), .Y(n_1199) );
CKINVDCx16_ASAP7_75t_R g1200 ( .A(n_1134), .Y(n_1200) );
AO21x2_ASAP7_75t_L g1201 ( .A1(n_1160), .A2(n_1167), .B(n_1143), .Y(n_1201) );
AOI21xp5_ASAP7_75t_SL g1202 ( .A1(n_1100), .A2(n_1101), .B(n_1107), .Y(n_1202) );
AOI21x1_ASAP7_75t_L g1203 ( .A1(n_1175), .A2(n_1182), .B(n_1149), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1033), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1205 ( .A(n_1100), .B(n_1046), .Y(n_1205) );
AOI221xp5_ASAP7_75t_L g1206 ( .A1(n_1105), .A2(n_1148), .B1(n_1053), .B2(n_1156), .C(n_1058), .Y(n_1206) );
INVxp67_ASAP7_75t_SL g1207 ( .A(n_1043), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1069), .B(n_1072), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1062), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1210 ( .A(n_1040), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1078), .B(n_1096), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1100), .B(n_1063), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1110), .B(n_1152), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_1107), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1161), .B(n_1048), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1086), .B(n_1087), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1147), .B(n_1040), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1086), .B(n_1087), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_1150), .A2(n_1177), .B1(n_1092), .B2(n_1058), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_1092), .A2(n_1050), .B1(n_1098), .B2(n_1155), .Y(n_1220) );
BUFx3_ASAP7_75t_L g1221 ( .A(n_1145), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1091), .Y(n_1222) );
INVx3_ASAP7_75t_L g1223 ( .A(n_1163), .Y(n_1223) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_1105), .A2(n_1148), .B1(n_1156), .B2(n_1155), .C(n_1128), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1166), .B(n_1176), .Y(n_1225) );
INVx1_ASAP7_75t_SL g1226 ( .A(n_1071), .Y(n_1226) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_1043), .Y(n_1227) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_1104), .B(n_1055), .C(n_1050), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1029), .Y(n_1229) );
OA21x2_ASAP7_75t_L g1230 ( .A1(n_1133), .A2(n_1039), .B(n_1117), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_1092), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1232 ( .A1(n_1060), .A2(n_1115), .B(n_1045), .C(n_1125), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1106), .B(n_1109), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1083), .B(n_1035), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1088), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_1098), .A2(n_1077), .B1(n_1080), .B2(n_1138), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1120), .B(n_1146), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1146), .B(n_1127), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_1098), .A2(n_1112), .B1(n_1114), .B2(n_1084), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1127), .B(n_1080), .Y(n_1240) );
OAI21xp33_ASAP7_75t_L g1241 ( .A1(n_1126), .A2(n_1089), .B(n_1132), .Y(n_1241) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_1147), .Y(n_1242) );
NOR2xp33_ASAP7_75t_L g1243 ( .A(n_1066), .B(n_1178), .Y(n_1243) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_1124), .A2(n_1131), .B1(n_1097), .B2(n_1036), .C(n_1159), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1119), .B(n_1142), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_1094), .Y(n_1246) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1102), .Y(n_1247) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_1173), .A2(n_1059), .B1(n_1085), .B2(n_1093), .Y(n_1248) );
INVx4_ASAP7_75t_L g1249 ( .A(n_1163), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1113), .Y(n_1250) );
AND2x4_ASAP7_75t_L g1251 ( .A(n_1099), .B(n_1030), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1113), .Y(n_1252) );
OA21x2_ASAP7_75t_L g1253 ( .A1(n_1052), .A2(n_1108), .B(n_1097), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1119), .B(n_1142), .Y(n_1254) );
AO21x2_ASAP7_75t_L g1255 ( .A1(n_1038), .A2(n_1172), .B(n_1074), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1073), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1034), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1119), .B(n_1142), .Y(n_1258) );
AOI21xp5_ASAP7_75t_SL g1259 ( .A1(n_1099), .A2(n_1169), .B(n_1076), .Y(n_1259) );
BUFx3_ASAP7_75t_L g1260 ( .A(n_1066), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_1065), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1034), .B(n_1047), .Y(n_1262) );
NAND2xp5_ASAP7_75t_SL g1263 ( .A(n_1168), .B(n_1179), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1183), .Y(n_1264) );
NOR2x1_ASAP7_75t_L g1265 ( .A(n_1030), .B(n_1076), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1034), .Y(n_1266) );
AO21x2_ASAP7_75t_L g1267 ( .A1(n_1074), .A2(n_1174), .B(n_1121), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1047), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1129), .B(n_1181), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1047), .B(n_1181), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1271 ( .A(n_1049), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1136), .B(n_1129), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1118), .Y(n_1273) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_1171), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1122), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1165), .B(n_1128), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1061), .A2(n_1153), .B1(n_1067), .B2(n_1162), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1116), .B(n_1170), .Y(n_1278) );
NAND2x1p5_ASAP7_75t_L g1279 ( .A(n_1135), .B(n_1111), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_1075), .B(n_1158), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1136), .B(n_1180), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1180), .B(n_1082), .Y(n_1282) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1111), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1079), .B(n_1082), .Y(n_1284) );
BUFx3_ASAP7_75t_L g1285 ( .A(n_1079), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1070), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1141), .B(n_1070), .Y(n_1287) );
INVx3_ASAP7_75t_L g1288 ( .A(n_1164), .Y(n_1288) );
AND2x4_ASAP7_75t_L g1289 ( .A(n_1144), .B(n_1151), .Y(n_1289) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_1164), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1154), .B(n_1140), .Y(n_1291) );
NAND4xp25_ASAP7_75t_L g1292 ( .A(n_1044), .B(n_1031), .C(n_1103), .D(n_1123), .Y(n_1292) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1154), .Y(n_1293) );
OAI21xp5_ASAP7_75t_L g1294 ( .A1(n_1130), .A2(n_1064), .B(n_1095), .Y(n_1294) );
AO21x2_ASAP7_75t_L g1295 ( .A1(n_1139), .A2(n_1160), .B(n_1157), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_1048), .A2(n_988), .B1(n_909), .B2(n_917), .Y(n_1296) );
AND2x4_ASAP7_75t_L g1297 ( .A(n_1090), .B(n_1101), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1028), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1028), .B(n_747), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1028), .B(n_747), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1028), .Y(n_1301) );
AO21x2_ASAP7_75t_L g1302 ( .A1(n_1157), .A2(n_1167), .B(n_1160), .Y(n_1302) );
OR2x6_ASAP7_75t_L g1303 ( .A(n_1100), .B(n_1107), .Y(n_1303) );
BUFx3_ASAP7_75t_L g1304 ( .A(n_1057), .Y(n_1304) );
OR2x6_ASAP7_75t_L g1305 ( .A(n_1100), .B(n_1107), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1068), .B(n_1069), .Y(n_1306) );
AO21x2_ASAP7_75t_L g1307 ( .A1(n_1157), .A2(n_1167), .B(n_1160), .Y(n_1307) );
INVx2_ASAP7_75t_SL g1308 ( .A(n_1057), .Y(n_1308) );
HB1xp67_ASAP7_75t_L g1309 ( .A(n_1107), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1310 ( .A(n_1150), .B(n_960), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_1048), .A2(n_988), .B1(n_909), .B2(n_917), .Y(n_1311) );
BUFx2_ASAP7_75t_L g1312 ( .A(n_1101), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1068), .B(n_1069), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1137), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1028), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1068), .B(n_1069), .Y(n_1316) );
AOI21x1_ASAP7_75t_L g1317 ( .A1(n_1175), .A2(n_1182), .B(n_1160), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1028), .Y(n_1318) );
BUFx3_ASAP7_75t_L g1319 ( .A(n_1260), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1237), .B(n_1272), .Y(n_1320) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_1229), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1188), .B(n_1191), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1225), .B(n_1269), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1237), .B(n_1272), .Y(n_1324) );
HB1xp67_ASAP7_75t_L g1325 ( .A(n_1312), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1195), .Y(n_1326) );
OAI321xp33_ASAP7_75t_L g1327 ( .A1(n_1220), .A2(n_1228), .A3(n_1303), .B1(n_1305), .B2(n_1206), .C(n_1198), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1196), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1245), .B(n_1254), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1245), .B(n_1254), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1225), .B(n_1269), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1258), .B(n_1270), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1197), .B(n_1209), .Y(n_1333) );
BUFx2_ASAP7_75t_L g1334 ( .A(n_1303), .Y(n_1334) );
AND2x4_ASAP7_75t_L g1335 ( .A(n_1249), .B(n_1223), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1258), .B(n_1270), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_1296), .A2(n_1311), .B1(n_1303), .B2(n_1305), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1298), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1262), .B(n_1238), .Y(n_1339) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1226), .B(n_1310), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1301), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1262), .B(n_1238), .Y(n_1342) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_1249), .B(n_1223), .Y(n_1343) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1193), .B(n_1213), .Y(n_1344) );
HB1xp67_ASAP7_75t_L g1345 ( .A(n_1312), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1315), .Y(n_1346) );
BUFx3_ASAP7_75t_L g1347 ( .A(n_1260), .Y(n_1347) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_1303), .Y(n_1348) );
INVx2_ASAP7_75t_SL g1349 ( .A(n_1185), .Y(n_1349) );
BUFx3_ASAP7_75t_L g1350 ( .A(n_1184), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1351 ( .A(n_1213), .B(n_1305), .Y(n_1351) );
AND2x4_ASAP7_75t_L g1352 ( .A(n_1249), .B(n_1223), .Y(n_1352) );
BUFx2_ASAP7_75t_L g1353 ( .A(n_1305), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1204), .B(n_1208), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1204), .B(n_1208), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1318), .Y(n_1356) );
BUFx6f_ASAP7_75t_L g1357 ( .A(n_1185), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1211), .B(n_1233), .Y(n_1358) );
INVxp67_ASAP7_75t_SL g1359 ( .A(n_1207), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1211), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1200), .B(n_1243), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1216), .B(n_1218), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1306), .B(n_1313), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1306), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1365 ( .A(n_1231), .Y(n_1365) );
HB1xp67_ASAP7_75t_L g1366 ( .A(n_1205), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1216), .B(n_1218), .Y(n_1367) );
CKINVDCx5p33_ASAP7_75t_R g1368 ( .A(n_1261), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1313), .Y(n_1369) );
AND2x4_ASAP7_75t_L g1370 ( .A(n_1251), .B(n_1265), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1316), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1190), .B(n_1257), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1212), .Y(n_1373) );
INVx2_ASAP7_75t_SL g1374 ( .A(n_1185), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1190), .B(n_1266), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_1236), .A2(n_1219), .B1(n_1202), .B2(n_1251), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1190), .B(n_1268), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1302), .B(n_1307), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1212), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1380 ( .A(n_1189), .Y(n_1380) );
BUFx2_ASAP7_75t_L g1381 ( .A(n_1189), .Y(n_1381) );
AND2x4_ASAP7_75t_L g1382 ( .A(n_1251), .B(n_1201), .Y(n_1382) );
BUFx2_ASAP7_75t_L g1383 ( .A(n_1227), .Y(n_1383) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_1201), .B(n_1302), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1281), .B(n_1246), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1275), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1205), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1302), .B(n_1307), .Y(n_1388) );
BUFx2_ASAP7_75t_L g1389 ( .A(n_1242), .Y(n_1389) );
INVx2_ASAP7_75t_SL g1390 ( .A(n_1185), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1205), .Y(n_1391) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_1242), .Y(n_1392) );
NOR2x1_ASAP7_75t_SL g1393 ( .A(n_1304), .B(n_1210), .Y(n_1393) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1186), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1297), .Y(n_1395) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_1304), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1307), .B(n_1201), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1297), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1281), .B(n_1297), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1400 ( .A(n_1217), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1240), .B(n_1282), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1276), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1240), .B(n_1282), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1404 ( .A(n_1192), .B(n_1214), .Y(n_1404) );
INVx1_ASAP7_75t_SL g1405 ( .A(n_1187), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1309), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1250), .B(n_1252), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1199), .B(n_1222), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1215), .B(n_1271), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1264), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1210), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1256), .Y(n_1412) );
AND2x4_ASAP7_75t_L g1413 ( .A(n_1217), .B(n_1308), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1273), .B(n_1300), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1299), .B(n_1308), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1314), .B(n_1295), .Y(n_1416) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1293), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_1217), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1358), .B(n_1224), .Y(n_1419) );
AND2x4_ASAP7_75t_SL g1420 ( .A(n_1335), .B(n_1239), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1332), .B(n_1295), .Y(n_1421) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1417), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1332), .B(n_1293), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1326), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1328), .Y(n_1425) );
BUFx2_ASAP7_75t_L g1426 ( .A(n_1319), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1336), .B(n_1230), .Y(n_1427) );
AND2x4_ASAP7_75t_SL g1428 ( .A(n_1335), .B(n_1194), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1358), .B(n_1363), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1336), .B(n_1230), .Y(n_1430) );
INVx4_ASAP7_75t_L g1431 ( .A(n_1319), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1339), .B(n_1230), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1338), .Y(n_1433) );
NAND4xp25_ASAP7_75t_L g1434 ( .A(n_1337), .B(n_1248), .C(n_1259), .D(n_1234), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1363), .B(n_1259), .Y(n_1435) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_1382), .B(n_1203), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1341), .Y(n_1437) );
INVx3_ASAP7_75t_L g1438 ( .A(n_1357), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1339), .B(n_1284), .Y(n_1439) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1394), .Y(n_1440) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_1382), .B(n_1317), .Y(n_1441) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1394), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1360), .B(n_1241), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1362), .B(n_1221), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1346), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1362), .B(n_1221), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1367), .B(n_1274), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1342), .B(n_1284), .Y(n_1448) );
CKINVDCx16_ASAP7_75t_R g1449 ( .A(n_1347), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1356), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1322), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1342), .B(n_1285), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1333), .Y(n_1453) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1327), .B(n_1232), .Y(n_1454) );
OAI22xp5_ASAP7_75t_L g1455 ( .A1(n_1376), .A2(n_1263), .B1(n_1277), .B2(n_1244), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1401), .B(n_1285), .Y(n_1456) );
INVx2_ASAP7_75t_SL g1457 ( .A(n_1347), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1401), .B(n_1291), .Y(n_1458) );
AND2x4_ASAP7_75t_L g1459 ( .A(n_1382), .B(n_1280), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1403), .B(n_1291), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1403), .B(n_1290), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1386), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1412), .Y(n_1463) );
OR2x2_ASAP7_75t_L g1464 ( .A(n_1367), .B(n_1278), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1410), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1407), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1320), .B(n_1235), .Y(n_1467) );
NOR2x1_ASAP7_75t_L g1468 ( .A(n_1350), .B(n_1280), .Y(n_1468) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_1409), .B(n_1261), .Y(n_1469) );
INVx2_ASAP7_75t_SL g1470 ( .A(n_1389), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1324), .B(n_1247), .Y(n_1471) );
INVx1_ASAP7_75t_SL g1472 ( .A(n_1405), .Y(n_1472) );
NOR2xp33_ASAP7_75t_L g1473 ( .A(n_1402), .B(n_1414), .Y(n_1473) );
AOI22xp5_ASAP7_75t_L g1474 ( .A1(n_1353), .A2(n_1289), .B1(n_1292), .B2(n_1255), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1409), .B(n_1286), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1324), .B(n_1283), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1364), .B(n_1253), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1321), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1329), .B(n_1283), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1369), .B(n_1253), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1329), .B(n_1286), .Y(n_1481) );
INVx2_ASAP7_75t_SL g1482 ( .A(n_1389), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1371), .B(n_1253), .Y(n_1483) );
OR2x2_ASAP7_75t_L g1484 ( .A(n_1323), .B(n_1267), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1330), .B(n_1288), .Y(n_1485) );
BUFx3_ASAP7_75t_L g1486 ( .A(n_1396), .Y(n_1486) );
INVx1_ASAP7_75t_SL g1487 ( .A(n_1361), .Y(n_1487) );
NOR4xp25_ASAP7_75t_SL g1488 ( .A(n_1353), .B(n_1348), .C(n_1334), .D(n_1368), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1489 ( .A(n_1392), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1424), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1432), .B(n_1372), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1492 ( .A(n_1429), .B(n_1331), .Y(n_1492) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1475), .B(n_1385), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1432), .B(n_1372), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1427), .B(n_1375), .Y(n_1495) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_1426), .Y(n_1496) );
INVx2_ASAP7_75t_L g1497 ( .A(n_1422), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1427), .B(n_1375), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1430), .B(n_1377), .Y(n_1499) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_1458), .B(n_1385), .Y(n_1500) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_1449), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1425), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1503 ( .A1(n_1434), .A2(n_1351), .B1(n_1392), .B2(n_1399), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1433), .Y(n_1504) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1437), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1473), .B(n_1354), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1507 ( .A(n_1473), .B(n_1355), .Y(n_1507) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1445), .Y(n_1508) );
NAND2x1p5_ASAP7_75t_L g1509 ( .A(n_1431), .B(n_1335), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1439), .B(n_1378), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1450), .Y(n_1511) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_1457), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1448), .B(n_1388), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1463), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1448), .B(n_1388), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1460), .B(n_1397), .Y(n_1516) );
INVx2_ASAP7_75t_SL g1517 ( .A(n_1457), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1462), .Y(n_1518) );
NAND2x2_ASAP7_75t_L g1519 ( .A(n_1435), .B(n_1351), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1419), .B(n_1355), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1440), .Y(n_1521) );
AOI32xp33_ASAP7_75t_L g1522 ( .A1(n_1454), .A2(n_1370), .A3(n_1404), .B1(n_1340), .B2(n_1343), .Y(n_1522) );
INVxp67_ASAP7_75t_L g1523 ( .A(n_1444), .Y(n_1523) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1466), .B(n_1408), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1460), .B(n_1384), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1421), .B(n_1384), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_1423), .B(n_1344), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1421), .B(n_1384), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1529 ( .A(n_1423), .B(n_1344), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1440), .Y(n_1530) );
NOR2xp33_ASAP7_75t_L g1531 ( .A(n_1487), .B(n_1368), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1485), .B(n_1416), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1485), .B(n_1467), .Y(n_1533) );
OR2x2_ASAP7_75t_L g1534 ( .A(n_1461), .B(n_1399), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1431), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1536 ( .A(n_1461), .B(n_1345), .Y(n_1536) );
NAND2x1p5_ASAP7_75t_L g1537 ( .A(n_1486), .B(n_1352), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1442), .Y(n_1538) );
NOR2xp67_ASAP7_75t_L g1539 ( .A(n_1454), .B(n_1325), .Y(n_1539) );
INVx1_ASAP7_75t_SL g1540 ( .A(n_1472), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1471), .B(n_1379), .Y(n_1541) );
INVxp67_ASAP7_75t_L g1542 ( .A(n_1446), .Y(n_1542) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1478), .B(n_1365), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1471), .B(n_1373), .Y(n_1544) );
NAND4xp25_ASAP7_75t_L g1545 ( .A(n_1522), .B(n_1455), .C(n_1474), .D(n_1443), .Y(n_1545) );
NAND2x1_ASAP7_75t_L g1546 ( .A(n_1539), .B(n_1468), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1547 ( .A(n_1500), .B(n_1476), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1490), .Y(n_1548) );
OR2x2_ASAP7_75t_L g1549 ( .A(n_1500), .B(n_1476), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1491), .B(n_1456), .Y(n_1550) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1490), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1511), .Y(n_1552) );
OAI21xp5_ASAP7_75t_L g1553 ( .A1(n_1503), .A2(n_1469), .B(n_1447), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1502), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1494), .B(n_1452), .Y(n_1555) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1504), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1505), .Y(n_1557) );
AOI21xp5_ASAP7_75t_L g1558 ( .A1(n_1535), .A2(n_1488), .B(n_1393), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1508), .Y(n_1559) );
NOR2xp33_ASAP7_75t_L g1560 ( .A(n_1540), .B(n_1464), .Y(n_1560) );
NAND3xp33_ASAP7_75t_L g1561 ( .A(n_1496), .B(n_1465), .C(n_1406), .Y(n_1561) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1514), .Y(n_1562) );
OAI21xp33_ASAP7_75t_SL g1563 ( .A1(n_1517), .A2(n_1470), .B(n_1489), .Y(n_1563) );
INVx1_ASAP7_75t_SL g1564 ( .A(n_1501), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1510), .B(n_1451), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1510), .B(n_1453), .Y(n_1566) );
OAI22xp5_ASAP7_75t_L g1567 ( .A1(n_1519), .A2(n_1428), .B1(n_1420), .B2(n_1370), .Y(n_1567) );
AND2x4_ASAP7_75t_L g1568 ( .A(n_1526), .B(n_1436), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1527), .B(n_1479), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1513), .B(n_1479), .Y(n_1570) );
INVx2_ASAP7_75t_SL g1571 ( .A(n_1517), .Y(n_1571) );
INVx1_ASAP7_75t_SL g1572 ( .A(n_1512), .Y(n_1572) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1497), .Y(n_1573) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1518), .Y(n_1574) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1527), .B(n_1481), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1529), .Y(n_1576) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1497), .Y(n_1577) );
INVxp67_ASAP7_75t_L g1578 ( .A(n_1543), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1529), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1494), .B(n_1452), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1495), .B(n_1481), .Y(n_1581) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1543), .Y(n_1582) );
NOR2xp67_ASAP7_75t_SL g1583 ( .A(n_1558), .B(n_1486), .Y(n_1583) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1548), .Y(n_1584) );
OAI22xp33_ASAP7_75t_L g1585 ( .A1(n_1545), .A2(n_1519), .B1(n_1509), .B2(n_1537), .Y(n_1585) );
INVx1_ASAP7_75t_SL g1586 ( .A(n_1564), .Y(n_1586) );
NAND2xp5_ASAP7_75t_SL g1587 ( .A(n_1563), .B(n_1509), .Y(n_1587) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1551), .Y(n_1588) );
OAI211xp5_ASAP7_75t_SL g1589 ( .A1(n_1553), .A2(n_1542), .B(n_1523), .C(n_1531), .Y(n_1589) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1552), .Y(n_1590) );
INVxp67_ASAP7_75t_L g1591 ( .A(n_1560), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1592 ( .A(n_1547), .B(n_1498), .Y(n_1592) );
INVx2_ASAP7_75t_L g1593 ( .A(n_1573), .Y(n_1593) );
OR2x2_ASAP7_75t_L g1594 ( .A(n_1549), .B(n_1498), .Y(n_1594) );
INVxp67_ASAP7_75t_SL g1595 ( .A(n_1561), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1596 ( .A(n_1569), .B(n_1499), .Y(n_1596) );
OAI32xp33_ASAP7_75t_L g1597 ( .A1(n_1572), .A2(n_1509), .A3(n_1537), .B1(n_1534), .B2(n_1536), .Y(n_1597) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1554), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1581), .B(n_1550), .Y(n_1599) );
BUFx3_ASAP7_75t_L g1600 ( .A(n_1571), .Y(n_1600) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1556), .Y(n_1601) );
AOI22xp5_ASAP7_75t_L g1602 ( .A1(n_1567), .A2(n_1526), .B1(n_1528), .B2(n_1520), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1603 ( .A(n_1578), .B(n_1513), .Y(n_1603) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1557), .Y(n_1604) );
OAI22xp33_ASAP7_75t_L g1605 ( .A1(n_1546), .A2(n_1537), .B1(n_1534), .B2(n_1536), .Y(n_1605) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1559), .Y(n_1606) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1562), .Y(n_1607) );
AOI222xp33_ASAP7_75t_L g1608 ( .A1(n_1595), .A2(n_1578), .B1(n_1560), .B2(n_1582), .C1(n_1579), .C2(n_1576), .Y(n_1608) );
OA22x2_ASAP7_75t_L g1609 ( .A1(n_1587), .A2(n_1428), .B1(n_1568), .B2(n_1420), .Y(n_1609) );
AOI211xp5_ASAP7_75t_L g1610 ( .A1(n_1585), .A2(n_1568), .B(n_1566), .C(n_1565), .Y(n_1610) );
OAI211xp5_ASAP7_75t_SL g1611 ( .A1(n_1585), .A2(n_1574), .B(n_1507), .C(n_1506), .Y(n_1611) );
INVxp67_ASAP7_75t_L g1612 ( .A(n_1586), .Y(n_1612) );
AOI211xp5_ASAP7_75t_L g1613 ( .A1(n_1587), .A2(n_1597), .B(n_1583), .C(n_1605), .Y(n_1613) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1584), .Y(n_1614) );
OAI22xp33_ASAP7_75t_L g1615 ( .A1(n_1602), .A2(n_1575), .B1(n_1570), .B2(n_1493), .Y(n_1615) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1588), .Y(n_1616) );
OAI21xp5_ASAP7_75t_L g1617 ( .A1(n_1589), .A2(n_1580), .B(n_1555), .Y(n_1617) );
AOI211xp5_ASAP7_75t_L g1618 ( .A1(n_1591), .A2(n_1528), .B(n_1370), .C(n_1525), .Y(n_1618) );
INVx1_ASAP7_75t_SL g1619 ( .A(n_1600), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_1599), .B(n_1515), .Y(n_1620) );
AOI221xp5_ASAP7_75t_L g1621 ( .A1(n_1598), .A2(n_1555), .B1(n_1525), .B2(n_1515), .C(n_1516), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1590), .Y(n_1622) );
AOI21xp33_ASAP7_75t_L g1623 ( .A1(n_1600), .A2(n_1414), .B(n_1387), .Y(n_1623) );
AOI21xp5_ASAP7_75t_L g1624 ( .A1(n_1613), .A2(n_1607), .B(n_1606), .Y(n_1624) );
AOI211xp5_ASAP7_75t_L g1625 ( .A1(n_1611), .A2(n_1603), .B(n_1604), .C(n_1601), .Y(n_1625) );
AOI22xp5_ASAP7_75t_L g1626 ( .A1(n_1608), .A2(n_1610), .B1(n_1609), .B2(n_1619), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1621), .B(n_1615), .Y(n_1627) );
NAND2xp33_ASAP7_75t_SL g1628 ( .A(n_1617), .B(n_1592), .Y(n_1628) );
OAI21xp33_ASAP7_75t_SL g1629 ( .A1(n_1619), .A2(n_1596), .B(n_1594), .Y(n_1629) );
NAND3xp33_ASAP7_75t_L g1630 ( .A(n_1612), .B(n_1593), .C(n_1411), .Y(n_1630) );
AOI211xp5_ASAP7_75t_SL g1631 ( .A1(n_1618), .A2(n_1359), .B(n_1352), .C(n_1343), .Y(n_1631) );
OAI211xp5_ASAP7_75t_SL g1632 ( .A1(n_1623), .A2(n_1492), .B(n_1391), .C(n_1524), .Y(n_1632) );
NAND2xp5_ASAP7_75t_SL g1633 ( .A(n_1629), .B(n_1614), .Y(n_1633) );
AOI21xp5_ASAP7_75t_L g1634 ( .A1(n_1628), .A2(n_1622), .B(n_1616), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1627), .B(n_1620), .Y(n_1635) );
NAND5xp2_ASAP7_75t_L g1636 ( .A(n_1626), .B(n_1383), .C(n_1398), .D(n_1395), .E(n_1279), .Y(n_1636) );
NAND3xp33_ASAP7_75t_SL g1637 ( .A(n_1631), .B(n_1381), .C(n_1380), .Y(n_1637) );
NOR5xp2_ASAP7_75t_L g1638 ( .A(n_1630), .B(n_1366), .C(n_1418), .D(n_1538), .E(n_1530), .Y(n_1638) );
AOI211xp5_ASAP7_75t_L g1639 ( .A1(n_1624), .A2(n_1343), .B(n_1352), .C(n_1441), .Y(n_1639) );
NOR5xp2_ASAP7_75t_L g1640 ( .A(n_1632), .B(n_1521), .C(n_1530), .D(n_1538), .E(n_1294), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1625), .B(n_1533), .Y(n_1641) );
NOR5xp2_ASAP7_75t_L g1642 ( .A(n_1640), .B(n_1436), .C(n_1482), .D(n_1349), .E(n_1390), .Y(n_1642) );
INVx2_ASAP7_75t_SL g1643 ( .A(n_1635), .Y(n_1643) );
NAND3xp33_ASAP7_75t_L g1644 ( .A(n_1633), .B(n_1577), .C(n_1573), .Y(n_1644) );
AND2x4_ASAP7_75t_L g1645 ( .A(n_1641), .B(n_1541), .Y(n_1645) );
OR5x1_ASAP7_75t_L g1646 ( .A(n_1637), .B(n_1400), .C(n_1482), .D(n_1413), .E(n_1415), .Y(n_1646) );
NAND4xp75_ASAP7_75t_L g1647 ( .A(n_1634), .B(n_1541), .C(n_1544), .D(n_1532), .Y(n_1647) );
XNOR2xp5_ASAP7_75t_L g1648 ( .A(n_1643), .B(n_1639), .Y(n_1648) );
OR4x1_ASAP7_75t_L g1649 ( .A(n_1646), .B(n_1636), .C(n_1638), .D(n_1349), .Y(n_1649) );
NAND3xp33_ASAP7_75t_L g1650 ( .A(n_1642), .B(n_1577), .C(n_1415), .Y(n_1650) );
INVx2_ASAP7_75t_L g1651 ( .A(n_1647), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1645), .B(n_1532), .Y(n_1652) );
INVx2_ASAP7_75t_L g1653 ( .A(n_1649), .Y(n_1653) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1651), .Y(n_1654) );
XNOR2xp5_ASAP7_75t_L g1655 ( .A(n_1648), .B(n_1644), .Y(n_1655) );
INVx2_ASAP7_75t_L g1656 ( .A(n_1650), .Y(n_1656) );
OA22x2_ASAP7_75t_L g1657 ( .A1(n_1654), .A2(n_1652), .B1(n_1650), .B2(n_1413), .Y(n_1657) );
BUFx2_ASAP7_75t_L g1658 ( .A(n_1653), .Y(n_1658) );
AO22x2_ASAP7_75t_L g1659 ( .A1(n_1656), .A2(n_1390), .B1(n_1374), .B2(n_1400), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1658), .B(n_1655), .Y(n_1660) );
AOI22xp5_ASAP7_75t_L g1661 ( .A1(n_1657), .A2(n_1459), .B1(n_1374), .B2(n_1255), .Y(n_1661) );
OAI21xp5_ASAP7_75t_SL g1662 ( .A1(n_1659), .A2(n_1459), .B(n_1484), .Y(n_1662) );
AOI222xp33_ASAP7_75t_L g1663 ( .A1(n_1660), .A2(n_1659), .B1(n_1438), .B2(n_1287), .C1(n_1483), .C2(n_1480), .Y(n_1663) );
NAND3xp33_ASAP7_75t_L g1664 ( .A(n_1661), .B(n_1662), .C(n_1357), .Y(n_1664) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1664), .Y(n_1665) );
AOI21xp5_ASAP7_75t_L g1666 ( .A1(n_1665), .A2(n_1663), .B(n_1477), .Y(n_1666) );
endmodule