module fake_jpeg_27478_n_295 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_270;
wire n_112;
wire n_199;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_37),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_29),
.B1(n_22),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_59),
.B1(n_71),
.B2(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_22),
.B2(n_23),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_30),
.B(n_26),
.C(n_27),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_68),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_38),
.C(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_20),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_73),
.B(n_83),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_30),
.B(n_27),
.C(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_36),
.B1(n_35),
.B2(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_77),
.B1(n_80),
.B2(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_31),
.B1(n_37),
.B2(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_48),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_18),
.B1(n_34),
.B2(n_3),
.Y(n_86)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_104),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_12),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_44),
.B1(n_43),
.B2(n_48),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_55),
.B1(n_69),
.B2(n_67),
.Y(n_123)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_17),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_115),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_74),
.B1(n_67),
.B2(n_56),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_116),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_54),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_54),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_95),
.B1(n_101),
.B2(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_47),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_150),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_48),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_133),
.B(n_136),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_47),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_47),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_97),
.B(n_111),
.C(n_93),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_1),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_53),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_136),
.B(n_126),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_56),
.B1(n_34),
.B2(n_4),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_94),
.B1(n_96),
.B2(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_1),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_162),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_123),
.B1(n_131),
.B2(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_126),
.B1(n_143),
.B2(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_167),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_92),
.C(n_106),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_130),
.C(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_90),
.B1(n_91),
.B2(n_116),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_142),
.B1(n_148),
.B2(n_134),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_92),
.B(n_88),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_89),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_117),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_104),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_149),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_124),
.B1(n_4),
.B2(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_127),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_98),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_130),
.B1(n_142),
.B2(n_148),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_193),
.B1(n_205),
.B2(n_157),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_205),
.B1(n_190),
.B2(n_200),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_16),
.C(n_15),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_202),
.C(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_166),
.C(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_205)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_181),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_215),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_161),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_222),
.B(n_162),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_223),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_165),
.B(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_153),
.B1(n_175),
.B2(n_154),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_185),
.B1(n_197),
.B2(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_224),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_222),
.B(n_185),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_202),
.C(n_191),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_158),
.C(n_168),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_196),
.B(n_200),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_229),
.B(n_178),
.C(n_158),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_252),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_186),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_195),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_194),
.C(n_201),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_230),
.C(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_265),
.C(n_270),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_238),
.B1(n_236),
.B2(n_211),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_254),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_211),
.B1(n_199),
.B2(n_235),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_251),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_250),
.B1(n_259),
.B2(n_233),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_156),
.B(n_233),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_257),
.C(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_264),
.C(n_275),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_269),
.B(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_271),
.B1(n_15),
.B2(n_13),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_7),
.B(n_8),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_280),
.C(n_283),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_289),
.A3(n_287),
.B1(n_290),
.B2(n_284),
.C1(n_10),
.C2(n_9),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_9),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_11),
.B(n_163),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_11),
.Y(n_295)
);


endmodule