module fake_jpeg_24682_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_42),
.C(n_36),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_54),
.B1(n_41),
.B2(n_39),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_60),
.B1(n_41),
.B2(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_27),
.B(n_30),
.C(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_16),
.B1(n_23),
.B2(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_32),
.B1(n_21),
.B2(n_22),
.Y(n_108)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_85),
.B1(n_53),
.B2(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_83),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_19),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_50),
.B1(n_40),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_92),
.B1(n_98),
.B2(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_40),
.B1(n_50),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_72),
.B2(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_55),
.B1(n_38),
.B2(n_25),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_25),
.C(n_38),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_101),
.C(n_75),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_38),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_67),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_80),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_38),
.B1(n_32),
.B2(n_21),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_68),
.B1(n_87),
.B2(n_70),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_38),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_80),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_97),
.B1(n_92),
.B2(n_89),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_117),
.B(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

OR2x4_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_118),
.B(n_122),
.Y(n_163)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_90),
.B1(n_102),
.B2(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_134),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_84),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_126),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_67),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_147),
.B1(n_124),
.B2(n_72),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_150),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_144),
.B(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_96),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_97),
.B1(n_91),
.B2(n_105),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_53),
.C(n_28),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_129),
.B(n_128),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_69),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_94),
.B(n_22),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_127),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_183),
.B(n_139),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_94),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_156),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_119),
.B1(n_131),
.B2(n_118),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_184),
.B1(n_139),
.B2(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_85),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_123),
.B1(n_114),
.B2(n_58),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_64),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_174),
.B(n_171),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_64),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_188),
.C(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_162),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_33),
.C(n_28),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_32),
.B(n_21),
.C(n_18),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_191),
.C(n_199),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_153),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_160),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_21),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_162),
.B1(n_150),
.B2(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_196),
.B1(n_206),
.B2(n_85),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_164),
.B1(n_159),
.B2(n_145),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_154),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_207),
.C(n_209),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_204),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_183),
.B(n_82),
.Y(n_216)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_163),
.B1(n_144),
.B2(n_143),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_157),
.C(n_103),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_23),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_123),
.C(n_114),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_170),
.B1(n_173),
.B2(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_184),
.B1(n_182),
.B2(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_215),
.B1(n_221),
.B2(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_209),
.B1(n_203),
.B2(n_197),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_172),
.B1(n_178),
.B2(n_176),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_172),
.B1(n_183),
.B2(n_188),
.Y(n_215)
);

OAI322xp33_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_207),
.A3(n_202),
.B1(n_192),
.B2(n_190),
.C1(n_200),
.C2(n_191),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_70),
.C(n_87),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_1),
.C(n_2),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_33),
.C(n_14),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_1),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_27),
.B1(n_20),
.B2(n_19),
.Y(n_222)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.C(n_29),
.Y(n_225)
);

OAI321xp33_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_9),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C(n_6),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_231),
.B1(n_222),
.B2(n_214),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_221),
.C(n_10),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_233),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.C(n_239),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_218),
.C(n_226),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.C(n_12),
.Y(n_248)
);

BUFx12f_ASAP7_75t_SL g239 ( 
.A(n_216),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_233),
.B(n_232),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_212),
.B1(n_213),
.B2(n_211),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_226),
.C(n_210),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_247),
.B(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_230),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_2),
.C(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_253),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_233),
.B1(n_232),
.B2(n_234),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_6),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_8),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_259),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_246),
.B(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_11),
.B(n_15),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_251),
.B1(n_15),
.B2(n_4),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_254),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_257),
.C(n_262),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_260),
.C(n_3),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_267),
.B(n_269),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_270),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_2),
.C(n_5),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_5),
.B(n_141),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_5),
.Y(n_276)
);


endmodule