module real_aes_7607_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g453 ( .A(n_1), .Y(n_453) );
INVx1_ASAP7_75t_L g181 ( .A(n_2), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_3), .A2(n_37), .B1(n_142), .B2(n_483), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g149 ( .A1(n_4), .A2(n_123), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_5), .B(n_116), .Y(n_466) );
AND2x6_ASAP7_75t_L g128 ( .A(n_6), .B(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_7), .A2(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_8), .B(n_38), .Y(n_105) );
INVx1_ASAP7_75t_L g156 ( .A(n_9), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_10), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g447 ( .A(n_12), .Y(n_447) );
INVx1_ASAP7_75t_L g237 ( .A(n_13), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_14), .B(n_164), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_15), .B(n_117), .Y(n_524) );
AO32x2_ASAP7_75t_L g496 ( .A1(n_16), .A2(n_116), .A3(n_161), .B1(n_475), .B2(n_497), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_17), .A2(n_99), .B1(n_738), .B2(n_747), .C1(n_756), .C2(n_762), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_17), .A2(n_107), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_17), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_18), .B(n_142), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_19), .B(n_137), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_20), .B(n_117), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_21), .A2(n_49), .B1(n_142), .B2(n_483), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_22), .B(n_123), .Y(n_193) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_23), .A2(n_74), .B1(n_142), .B2(n_164), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_24), .B(n_142), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_25), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_26), .A2(n_235), .B(n_236), .C(n_238), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_27), .Y(n_755) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_28), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_29), .B(n_158), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_30), .B(n_154), .Y(n_183) );
INVx1_ASAP7_75t_L g170 ( .A(n_31), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_32), .B(n_158), .Y(n_513) );
INVx2_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_34), .B(n_142), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_35), .B(n_158), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_36), .A2(n_128), .B(n_132), .C(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g168 ( .A(n_39), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_40), .B(n_154), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_41), .B(n_142), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_42), .A2(n_84), .B1(n_200), .B2(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_43), .B(n_142), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_44), .B(n_142), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_45), .Y(n_171) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_46), .A2(n_100), .B1(n_726), .B2(n_727), .C1(n_732), .C2(n_737), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_46), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_47), .B(n_452), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_48), .B(n_123), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_50), .A2(n_59), .B1(n_142), .B2(n_164), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_51), .A2(n_132), .B1(n_164), .B2(n_166), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_52), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_53), .B(n_142), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_54), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_55), .B(n_142), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_56), .A2(n_141), .B(n_153), .C(n_155), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_57), .Y(n_213) );
INVx1_ASAP7_75t_L g151 ( .A(n_58), .Y(n_151) );
INVx1_ASAP7_75t_L g129 ( .A(n_60), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_61), .B(n_142), .Y(n_454) );
INVx1_ASAP7_75t_L g120 ( .A(n_62), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_63), .Y(n_743) );
AO32x2_ASAP7_75t_L g480 ( .A1(n_64), .A2(n_116), .A3(n_217), .B1(n_475), .B2(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g473 ( .A(n_65), .Y(n_473) );
INVx1_ASAP7_75t_L g508 ( .A(n_66), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_67), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_SL g136 ( .A1(n_68), .A2(n_137), .B(n_138), .C(n_141), .Y(n_136) );
INVxp67_ASAP7_75t_L g139 ( .A(n_69), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_70), .B(n_164), .Y(n_509) );
INVx1_ASAP7_75t_L g742 ( .A(n_71), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_72), .Y(n_174) );
INVx1_ASAP7_75t_L g206 ( .A(n_73), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_75), .A2(n_128), .B(n_132), .C(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_76), .B(n_483), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_77), .B(n_164), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_78), .B(n_182), .Y(n_196) );
INVx2_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_80), .B(n_137), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_81), .B(n_164), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_82), .A2(n_128), .B(n_132), .C(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g102 ( .A(n_83), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g434 ( .A(n_83), .Y(n_434) );
OR2x2_ASAP7_75t_L g746 ( .A(n_83), .B(n_736), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_85), .A2(n_97), .B1(n_164), .B2(n_165), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_86), .B(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_87), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_88), .A2(n_128), .B(n_132), .C(n_220), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_89), .Y(n_227) );
INVx1_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_91), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_92), .B(n_182), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_93), .B(n_164), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_94), .B(n_116), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_95), .A2(n_123), .B(n_130), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_96), .B(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_106), .B1(n_432), .B2(n_435), .Y(n_100) );
INVx2_ASAP7_75t_L g729 ( .A(n_101), .Y(n_729) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x2_ASAP7_75t_L g433 ( .A(n_103), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g736 ( .A(n_103), .Y(n_736) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_107), .A2(n_728), .B1(n_730), .B2(n_731), .Y(n_727) );
INVx2_ASAP7_75t_L g751 ( .A(n_107), .Y(n_751) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND4x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_350), .C(n_397), .D(n_417), .Y(n_108) );
NOR3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_280), .C(n_305), .Y(n_109) );
OAI211xp5_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_188), .B(n_240), .C(n_270), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_159), .Y(n_112) );
INVx3_ASAP7_75t_SL g322 ( .A(n_113), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_113), .B(n_253), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_113), .B(n_175), .Y(n_403) );
AND2x2_ASAP7_75t_L g426 ( .A(n_113), .B(n_292), .Y(n_426) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_147), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g244 ( .A(n_115), .B(n_148), .Y(n_244) );
INVx3_ASAP7_75t_L g257 ( .A(n_115), .Y(n_257) );
AND2x2_ASAP7_75t_L g262 ( .A(n_115), .B(n_147), .Y(n_262) );
OR2x2_ASAP7_75t_L g313 ( .A(n_115), .B(n_254), .Y(n_313) );
BUFx2_ASAP7_75t_L g333 ( .A(n_115), .Y(n_333) );
AND2x2_ASAP7_75t_L g343 ( .A(n_115), .B(n_254), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_115), .B(n_160), .Y(n_349) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_122), .B(n_144), .Y(n_115) );
INVx4_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_116), .A2(n_459), .B(n_466), .Y(n_458) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_118), .B(n_119), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
BUFx2_ASAP7_75t_L g231 ( .A(n_123), .Y(n_231) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_124), .B(n_128), .Y(n_172) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx1_ASAP7_75t_L g452 ( .A(n_125), .Y(n_452) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
INVx1_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx1_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
INVx1_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
INVx3_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_127), .Y(n_167) );
INVx4_ASAP7_75t_SL g143 ( .A(n_128), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_128), .A2(n_446), .B(n_450), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_128), .A2(n_460), .B(n_463), .Y(n_459) );
BUFx3_ASAP7_75t_L g475 ( .A(n_128), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_128), .A2(n_488), .B(n_492), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_128), .A2(n_507), .B(n_510), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B(n_136), .C(n_143), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_131), .A2(n_143), .B(n_151), .C(n_152), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_131), .A2(n_143), .B(n_233), .C(n_234), .Y(n_232) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_133), .Y(n_142) );
BUFx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
INVx1_ASAP7_75t_L g483 ( .A(n_133), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_137), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_140), .B(n_156), .Y(n_155) );
INVx5_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_140), .A2(n_154), .B1(n_482), .B2(n_484), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_SL g507 ( .A1(n_141), .A2(n_182), .B(n_508), .C(n_509), .Y(n_507) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_163), .B1(n_171), .B2(n_172), .Y(n_162) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_145), .A2(n_149), .B(n_157), .Y(n_148) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_146), .B(n_203), .Y(n_202) );
AO21x1_ASAP7_75t_L g519 ( .A1(n_146), .A2(n_520), .B(n_523), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_146), .B(n_475), .C(n_520), .Y(n_538) );
INVx1_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_148), .B(n_254), .Y(n_268) );
INVx2_ASAP7_75t_L g278 ( .A(n_148), .Y(n_278) );
AND2x2_ASAP7_75t_L g291 ( .A(n_148), .B(n_257), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_148), .B(n_254), .Y(n_302) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_148), .B(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g360 ( .A(n_148), .Y(n_360) );
AND2x2_ASAP7_75t_L g406 ( .A(n_148), .B(n_160), .Y(n_406) );
O2A1O1Ixp5_ASAP7_75t_L g472 ( .A1(n_153), .A2(n_451), .B(n_473), .C(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_153), .A2(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx4_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_154), .A2(n_455), .B1(n_498), .B2(n_499), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_154), .A2(n_455), .B1(n_521), .B2(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx2_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_158), .A2(n_230), .B(n_239), .Y(n_229) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_158), .A2(n_487), .B(n_495), .Y(n_486) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_158), .A2(n_506), .B(n_513), .Y(n_505) );
INVx3_ASAP7_75t_SL g279 ( .A(n_159), .Y(n_279) );
OR2x2_ASAP7_75t_L g332 ( .A(n_159), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_175), .Y(n_159) );
INVx3_ASAP7_75t_L g254 ( .A(n_160), .Y(n_254) );
AND2x2_ASAP7_75t_L g321 ( .A(n_160), .B(n_176), .Y(n_321) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_160), .Y(n_389) );
AOI33xp33_ASAP7_75t_L g393 ( .A1(n_160), .A2(n_322), .A3(n_329), .B1(n_338), .B2(n_394), .B3(n_395), .Y(n_393) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_173), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_161), .B(n_174), .Y(n_173) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_161), .A2(n_177), .B(n_185), .Y(n_176) );
INVx2_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
INVx2_ASAP7_75t_L g184 ( .A(n_164), .Y(n_184) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_166) );
INVx2_ASAP7_75t_L g169 ( .A(n_167), .Y(n_169) );
INVx4_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_172), .A2(n_178), .B(n_179), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_172), .A2(n_206), .B(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_175), .B(n_257), .Y(n_256) );
NOR3xp33_ASAP7_75t_L g316 ( .A(n_175), .B(n_317), .C(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g342 ( .A(n_175), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_175), .B(n_349), .Y(n_352) );
AND2x2_ASAP7_75t_L g405 ( .A(n_175), .B(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
OR2x2_ASAP7_75t_L g355 ( .A(n_176), .B(n_254), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g455 ( .A(n_182), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_182), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_182), .A2(n_470), .B(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_184), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_187), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_187), .B(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_214), .Y(n_188) );
AOI32xp33_ASAP7_75t_L g306 ( .A1(n_189), .A2(n_307), .A3(n_309), .B1(n_311), .B2(n_314), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_189), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g409 ( .A(n_189), .Y(n_409) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g341 ( .A(n_190), .B(n_325), .Y(n_341) );
AND2x2_ASAP7_75t_L g361 ( .A(n_190), .B(n_287), .Y(n_361) );
AND2x2_ASAP7_75t_L g429 ( .A(n_190), .B(n_347), .Y(n_429) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_204), .Y(n_190) );
INVx3_ASAP7_75t_L g250 ( .A(n_191), .Y(n_250) );
AND2x2_ASAP7_75t_L g264 ( .A(n_191), .B(n_248), .Y(n_264) );
OR2x2_ASAP7_75t_L g269 ( .A(n_191), .B(n_247), .Y(n_269) );
INVx1_ASAP7_75t_L g276 ( .A(n_191), .Y(n_276) );
AND2x2_ASAP7_75t_L g284 ( .A(n_191), .B(n_258), .Y(n_284) );
AND2x2_ASAP7_75t_L g286 ( .A(n_191), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_191), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g339 ( .A(n_191), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_191), .B(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
AOI21xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B(n_201), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_198), .A2(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
INVx1_ASAP7_75t_L g211 ( .A(n_201), .Y(n_211) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_201), .A2(n_445), .B(n_456), .Y(n_444) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_201), .A2(n_468), .B(n_476), .Y(n_467) );
INVx2_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
AND2x2_ASAP7_75t_L g294 ( .A(n_204), .B(n_215), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_204), .B(n_229), .Y(n_304) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_204) );
INVx2_ASAP7_75t_L g424 ( .A(n_214), .Y(n_424) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_215), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g265 ( .A(n_215), .Y(n_265) );
AND2x2_ASAP7_75t_L g309 ( .A(n_215), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g325 ( .A(n_215), .B(n_288), .Y(n_325) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g273 ( .A(n_216), .Y(n_273) );
AND2x2_ASAP7_75t_L g287 ( .A(n_216), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g338 ( .A(n_216), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_216), .B(n_248), .Y(n_370) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_226), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_225), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_224), .Y(n_220) );
AND2x2_ASAP7_75t_L g249 ( .A(n_228), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g310 ( .A(n_228), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_228), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g347 ( .A(n_228), .Y(n_347) );
INVx1_ASAP7_75t_L g380 ( .A(n_228), .Y(n_380) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g258 ( .A(n_229), .B(n_248), .Y(n_258) );
INVx1_ASAP7_75t_L g288 ( .A(n_229), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_235), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g449 ( .A(n_235), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_235), .A2(n_511), .B(n_512), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .B1(n_251), .B2(n_258), .C(n_259), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_242), .B(n_262), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_242), .B(n_325), .Y(n_402) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_244), .B(n_292), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_244), .B(n_253), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_244), .B(n_267), .Y(n_396) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g318 ( .A(n_248), .Y(n_318) );
AND2x2_ASAP7_75t_L g293 ( .A(n_249), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g371 ( .A(n_249), .Y(n_371) );
AND2x2_ASAP7_75t_L g303 ( .A(n_250), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_250), .B(n_273), .Y(n_319) );
AND2x2_ASAP7_75t_L g383 ( .A(n_250), .B(n_309), .Y(n_383) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g292 ( .A(n_254), .B(n_261), .Y(n_292) );
AND2x2_ASAP7_75t_L g388 ( .A(n_255), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_257), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_258), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_258), .B(n_265), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_258), .B(n_273), .Y(n_373) );
AND2x2_ASAP7_75t_L g394 ( .A(n_258), .B(n_338), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .A3(n_265), .B1(n_266), .B2(n_269), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_SL g267 ( .A(n_261), .Y(n_267) );
NAND2x1_ASAP7_75t_L g308 ( .A(n_261), .B(n_291), .Y(n_308) );
OR2x2_ASAP7_75t_L g312 ( .A(n_261), .B(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_261), .B(n_360), .Y(n_413) );
INVx1_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_263), .A2(n_354), .B1(n_400), .B2(n_403), .C(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g271 ( .A(n_264), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g314 ( .A(n_264), .B(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_264), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_264), .B(n_325), .Y(n_392) );
INVxp67_ASAP7_75t_L g328 ( .A(n_265), .Y(n_328) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g398 ( .A(n_267), .B(n_385), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_267), .B(n_348), .Y(n_421) );
INVx1_ASAP7_75t_L g296 ( .A(n_269), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_269), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g414 ( .A(n_269), .B(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_274), .B(n_277), .Y(n_270) );
AND2x2_ASAP7_75t_L g283 ( .A(n_272), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g367 ( .A(n_276), .B(n_287), .Y(n_367) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g385 ( .A(n_278), .B(n_343), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_278), .B(n_342), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_279), .B(n_291), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_285), .C(n_295), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_281), .A2(n_316), .B1(n_320), .B2(n_323), .C(n_326), .Y(n_315) );
AOI31xp33_ASAP7_75t_L g410 ( .A1(n_281), .A2(n_411), .A3(n_412), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B1(n_291), .B2(n_293), .Y(n_285) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g411 ( .A(n_291), .Y(n_411) );
INVx1_ASAP7_75t_L g374 ( .A(n_292), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g417 ( .A1(n_294), .A2(n_418), .B(n_420), .C(n_422), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B1(n_299), .B2(n_303), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_300), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI221xp5_ASAP7_75t_SL g390 ( .A1(n_302), .A2(n_336), .B1(n_355), .B2(n_391), .C(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g386 ( .A(n_303), .Y(n_386) );
INVx1_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
NAND3xp33_ASAP7_75t_SL g305 ( .A(n_306), .B(n_315), .C(n_330), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_307), .A2(n_357), .B(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_309), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g416 ( .A(n_310), .Y(n_416) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_337), .Y(n_354) );
INVx1_ASAP7_75t_L g329 ( .A(n_318), .Y(n_329) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g327 ( .A(n_321), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_321), .B(n_359), .Y(n_358) );
NOR4xp25_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .C(n_328), .D(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_341), .B2(n_342), .C1(n_344), .C2(n_348), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx1_ASAP7_75t_L g428 ( .A(n_332), .Y(n_428) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_344), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_349), .A2(n_405), .B(n_407), .Y(n_404) );
NOR4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_362), .C(n_375), .D(n_390), .Y(n_350) );
OAI221xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_353), .B1(n_354), .B2(n_355), .C(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g431 ( .A(n_352), .Y(n_431) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_359), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OAI222xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_368), .B2(n_369), .C1(n_372), .C2(n_374), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_398), .B(n_399), .C(n_410), .Y(n_397) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OAI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_381), .B1(n_382), .B2(n_384), .C1(n_386), .C2(n_387), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_392), .A2(n_395), .B1(n_428), .B2(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI211xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_425), .B(n_427), .C(n_430), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx6_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g730 ( .A(n_433), .Y(n_730) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_434), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g731 ( .A(n_435), .Y(n_731) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_692), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_596), .C(n_680), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_539), .C(n_561), .D(n_577), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_477), .B1(n_500), .B2(n_518), .C(n_525), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_457), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_441), .B(n_518), .Y(n_551) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_441), .B(n_579), .C(n_592), .D(n_594), .Y(n_591) );
INVxp67_ASAP7_75t_L g708 ( .A(n_441), .Y(n_708) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g590 ( .A(n_442), .B(n_528), .Y(n_590) );
AND2x2_ASAP7_75t_L g614 ( .A(n_442), .B(n_457), .Y(n_614) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g581 ( .A(n_443), .B(n_517), .Y(n_581) );
AND2x2_ASAP7_75t_L g621 ( .A(n_443), .B(n_602), .Y(n_621) );
AND2x2_ASAP7_75t_L g638 ( .A(n_443), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_443), .B(n_458), .Y(n_662) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g516 ( .A(n_444), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g533 ( .A(n_444), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g545 ( .A(n_444), .B(n_458), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_444), .B(n_467), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B(n_454), .C(n_455), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_455), .A2(n_464), .B(n_465), .Y(n_463) );
AND2x2_ASAP7_75t_L g548 ( .A(n_457), .B(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_457), .A2(n_598), .B1(n_601), .B2(n_603), .C(n_607), .Y(n_597) );
AND2x2_ASAP7_75t_L g656 ( .A(n_457), .B(n_621), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_457), .B(n_638), .Y(n_690) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
INVx3_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
AND2x2_ASAP7_75t_L g565 ( .A(n_458), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g619 ( .A(n_458), .B(n_534), .Y(n_619) );
AND2x2_ASAP7_75t_L g677 ( .A(n_458), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g518 ( .A(n_467), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g534 ( .A(n_467), .Y(n_534) );
INVx1_ASAP7_75t_L g589 ( .A(n_467), .Y(n_589) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_467), .Y(n_595) );
AND2x2_ASAP7_75t_L g640 ( .A(n_467), .B(n_517), .Y(n_640) );
OR2x2_ASAP7_75t_L g679 ( .A(n_467), .B(n_519), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B(n_475), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_477), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
AND2x2_ASAP7_75t_L g675 ( .A(n_478), .B(n_672), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_478), .B(n_657), .Y(n_707) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g606 ( .A(n_479), .B(n_530), .Y(n_606) );
AND2x2_ASAP7_75t_L g655 ( .A(n_479), .B(n_503), .Y(n_655) );
INVx1_ASAP7_75t_L g701 ( .A(n_479), .Y(n_701) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_480), .Y(n_515) );
AND2x2_ASAP7_75t_L g556 ( .A(n_480), .B(n_530), .Y(n_556) );
INVx1_ASAP7_75t_L g573 ( .A(n_480), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_480), .B(n_496), .Y(n_579) );
AND2x2_ASAP7_75t_L g647 ( .A(n_485), .B(n_555), .Y(n_647) );
INVx2_ASAP7_75t_L g712 ( .A(n_485), .Y(n_712) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g529 ( .A(n_486), .B(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g542 ( .A(n_486), .B(n_504), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_486), .B(n_503), .Y(n_570) );
INVx1_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
INVx1_ASAP7_75t_L g593 ( .A(n_486), .Y(n_593) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_486), .Y(n_605) );
INVx2_ASAP7_75t_L g673 ( .A(n_486), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .Y(n_488) );
INVx2_ASAP7_75t_L g530 ( .A(n_496), .Y(n_530) );
BUFx2_ASAP7_75t_L g627 ( .A(n_496), .Y(n_627) );
AND2x2_ASAP7_75t_L g672 ( .A(n_496), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_514), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_502), .B(n_609), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_502), .A2(n_671), .B(n_685), .Y(n_695) );
AND2x2_ASAP7_75t_L g720 ( .A(n_502), .B(n_606), .Y(n_720) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g642 ( .A(n_504), .Y(n_642) );
AND2x2_ASAP7_75t_L g671 ( .A(n_504), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_505), .Y(n_555) );
INVx2_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_505), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g528 ( .A(n_515), .Y(n_528) );
OR2x2_ASAP7_75t_L g541 ( .A(n_515), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g609 ( .A(n_515), .B(n_605), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_515), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g710 ( .A(n_515), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_515), .B(n_647), .Y(n_722) );
AND2x2_ASAP7_75t_L g601 ( .A(n_516), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g624 ( .A(n_516), .B(n_518), .Y(n_624) );
INVx2_ASAP7_75t_L g536 ( .A(n_517), .Y(n_536) );
AND2x2_ASAP7_75t_L g564 ( .A(n_517), .B(n_537), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_517), .B(n_589), .Y(n_645) );
AND2x2_ASAP7_75t_L g559 ( .A(n_518), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g706 ( .A(n_518), .Y(n_706) );
AND2x2_ASAP7_75t_L g718 ( .A(n_518), .B(n_581), .Y(n_718) );
AND2x2_ASAP7_75t_L g544 ( .A(n_519), .B(n_534), .Y(n_544) );
INVx1_ASAP7_75t_L g639 ( .A(n_519), .Y(n_639) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g537 ( .A(n_524), .B(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_528), .B(n_575), .Y(n_584) );
OR2x2_ASAP7_75t_L g716 ( .A(n_528), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g633 ( .A(n_529), .B(n_574), .Y(n_633) );
AND2x2_ASAP7_75t_L g641 ( .A(n_529), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g700 ( .A(n_529), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g724 ( .A(n_529), .B(n_571), .Y(n_724) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_530), .B(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g711 ( .A(n_530), .B(n_574), .Y(n_711) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g563 ( .A(n_533), .B(n_564), .Y(n_563) );
INVxp67_ASAP7_75t_L g725 ( .A(n_533), .Y(n_725) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g560 ( .A(n_536), .Y(n_560) );
AND2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_544), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_536), .B(n_679), .Y(n_705) );
INVx2_ASAP7_75t_L g550 ( .A(n_537), .Y(n_550) );
INVx3_ASAP7_75t_L g602 ( .A(n_537), .Y(n_602) );
OR2x2_ASAP7_75t_L g630 ( .A(n_537), .B(n_631), .Y(n_630) );
AOI311xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .A3(n_545), .B(n_546), .C(n_557), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g577 ( .A1(n_540), .A2(n_578), .B(n_580), .C(n_582), .Y(n_577) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g562 ( .A(n_542), .Y(n_562) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g580 ( .A(n_544), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_544), .B(n_560), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_544), .B(n_545), .Y(n_713) );
AND2x2_ASAP7_75t_L g635 ( .A(n_545), .B(n_549), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_551), .B(n_552), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g693 ( .A(n_549), .B(n_581), .Y(n_693) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_550), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g587 ( .A(n_550), .Y(n_587) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g578 ( .A(n_554), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g623 ( .A(n_556), .Y(n_623) );
AND2x4_ASAP7_75t_L g685 ( .A(n_556), .B(n_654), .Y(n_685) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_559), .A2(n_625), .B1(n_637), .B2(n_641), .C1(n_643), .C2(n_647), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_565), .C(n_568), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_562), .B(n_606), .Y(n_629) );
INVx1_ASAP7_75t_L g651 ( .A(n_564), .Y(n_651) );
INVx1_ASAP7_75t_L g585 ( .A(n_566), .Y(n_585) );
OR2x2_ASAP7_75t_L g650 ( .A(n_567), .B(n_651), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_571), .B(n_575), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_569), .B(n_587), .C(n_588), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_569), .A2(n_606), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_573), .Y(n_626) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_574), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g683 ( .A(n_574), .Y(n_683) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_574), .Y(n_699) );
INVx2_ASAP7_75t_L g657 ( .A(n_575), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_579), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g631 ( .A(n_581), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B1(n_586), .B2(n_590), .C(n_591), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_585), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g719 ( .A(n_585), .Y(n_719) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g600 ( .A(n_592), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_592), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g658 ( .A(n_592), .B(n_606), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_592), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g691 ( .A(n_592), .B(n_626), .Y(n_691) );
BUFx3_ASAP7_75t_L g654 ( .A(n_593), .Y(n_654) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND5xp2_ASAP7_75t_L g596 ( .A(n_597), .B(n_615), .C(n_636), .D(n_648), .E(n_663), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI32xp33_ASAP7_75t_L g688 ( .A1(n_600), .A2(n_627), .A3(n_643), .B1(n_689), .B2(n_691), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_602), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g612 ( .A(n_606), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_624), .B2(n_625), .C(n_628), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g687 ( .A(n_619), .B(n_638), .Y(n_687) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_624), .A2(n_685), .B1(n_703), .B2(n_708), .C(n_709), .Y(n_702) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_L g668 ( .A(n_627), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_632), .B2(n_634), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g646 ( .A(n_638), .Y(n_646) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B1(n_656), .B2(n_657), .C1(n_658), .C2(n_659), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_657), .A2(n_704), .B1(n_706), .B2(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_669), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_674), .B(n_676), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g717 ( .A(n_672), .Y(n_717) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_686), .C(n_688), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_696), .C(n_721), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_693), .Y(n_697) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_702), .C(n_714), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B(n_713), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_744), .Y(n_739) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_SL g761 ( .A(n_741), .Y(n_761) );
INVx1_ASAP7_75t_L g760 ( .A(n_743), .Y(n_760) );
OA21x2_ASAP7_75t_L g763 ( .A1(n_743), .A2(n_752), .B(n_761), .Y(n_763) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g752 ( .A(n_746), .Y(n_752) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_746), .Y(n_754) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_753), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g753 ( .A(n_754), .B(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
CKINVDCx6p67_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
endmodule