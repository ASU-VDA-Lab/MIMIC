module fake_jpeg_30469_n_452 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_452);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_349;
wire n_21;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_20),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_82),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_79),
.Y(n_103)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_20),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_80),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_32),
.B(n_0),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_89),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_29),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_102),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_40),
.CON(n_97),
.SN(n_97)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_97),
.B(n_74),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_137),
.Y(n_146)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_56),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_45),
.B(n_43),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_75),
.Y(n_149)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_52),
.C(n_50),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_40),
.C(n_41),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_22),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_151),
.Y(n_179)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_168),
.B(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_22),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_40),
.B1(n_79),
.B2(n_42),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_174),
.B1(n_176),
.B2(n_49),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_92),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_177),
.B1(n_40),
.B2(n_57),
.Y(n_184)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_39),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_161),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_172),
.Y(n_196)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_128),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_97),
.B(n_39),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_58),
.B(n_53),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_39),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_91),
.Y(n_191)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_66),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_124),
.Y(n_180)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_118),
.A2(n_70),
.B1(n_62),
.B2(n_65),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_118),
.B1(n_105),
.B2(n_113),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_199),
.B1(n_175),
.B2(n_173),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_182),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_121),
.B1(n_127),
.B2(n_113),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_139),
.B1(n_119),
.B2(n_42),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_197),
.B(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_119),
.B1(n_42),
.B2(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_144),
.A2(n_105),
.B1(n_127),
.B2(n_121),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_123),
.B1(n_96),
.B2(n_81),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_72),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_165),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_228),
.B1(n_199),
.B2(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_146),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_145),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_143),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_142),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_180),
.C(n_182),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_196),
.C(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_174),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

BUFx4f_ASAP7_75t_SL g229 ( 
.A(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_184),
.B1(n_224),
.B2(n_214),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_186),
.B(n_192),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_250),
.B(n_229),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_196),
.C(n_197),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_190),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_181),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_191),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_190),
.B(n_200),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_222),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_166),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_203),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_211),
.B1(n_207),
.B2(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_203),
.B1(n_185),
.B2(n_170),
.Y(n_276)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_220),
.B1(n_203),
.B2(n_228),
.Y(n_256)
);

AO22x2_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_243),
.B1(n_231),
.B2(n_249),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_215),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_258),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_276),
.B1(n_232),
.B2(n_247),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_226),
.B1(n_218),
.B2(n_217),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_274),
.B1(n_275),
.B2(n_254),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_278),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_236),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_200),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_265),
.B(n_268),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_236),
.B(n_238),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_229),
.B(n_212),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_253),
.B(n_231),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_230),
.B1(n_221),
.B2(n_229),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_254),
.B1(n_232),
.B2(n_253),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_244),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_221),
.B1(n_227),
.B2(n_185),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_213),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_260),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_246),
.C(n_234),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.C(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_206),
.B1(n_150),
.B2(n_153),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_289),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_246),
.C(n_237),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_237),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_303),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_290),
.A2(n_294),
.B1(n_194),
.B2(n_266),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_231),
.B1(n_247),
.B2(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_243),
.C(n_244),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_110),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_270),
.B(n_43),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_304),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_201),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_260),
.B(n_248),
.CI(n_245),
.CON(n_304),
.SN(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_201),
.C(n_194),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_262),
.C(n_278),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_280),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_306),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_245),
.B1(n_248),
.B2(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_263),
.B1(n_255),
.B2(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_283),
.C(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_321),
.C(n_332),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_267),
.B(n_269),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_276),
.C(n_281),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_SL g322 ( 
.A(n_295),
.B(n_266),
.C(n_271),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_322),
.B(n_304),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_308),
.B1(n_316),
.B2(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_223),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_288),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_328),
.A2(n_330),
.B1(n_336),
.B2(n_293),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_297),
.A2(n_206),
.B1(n_110),
.B2(n_136),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_58),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_198),
.C(n_148),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_53),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_297),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_198),
.C(n_167),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_335),
.C(n_332),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_156),
.C(n_160),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_153),
.B1(n_96),
.B2(n_123),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_107),
.B1(n_91),
.B2(n_76),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_323),
.B(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_344),
.Y(n_372)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_345),
.A2(n_356),
.B1(n_340),
.B2(n_355),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_304),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_351),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_321),
.A2(n_307),
.B(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_348),
.B(n_346),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_350),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_313),
.A2(n_308),
.B1(n_306),
.B2(n_296),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_307),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_282),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_361),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_296),
.B1(n_301),
.B2(n_293),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_324),
.A2(n_171),
.B1(n_172),
.B2(n_176),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_333),
.A2(n_141),
.B1(n_155),
.B2(n_101),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_162),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_356),
.B(n_359),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_36),
.B1(n_159),
.B2(n_33),
.Y(n_358)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_358),
.A2(n_29),
.A3(n_36),
.B1(n_107),
.B2(n_68),
.C1(n_21),
.C2(n_30),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_311),
.C(n_314),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_377),
.C(n_339),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_311),
.C(n_329),
.Y(n_363)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

OAI22x1_ASAP7_75t_SL g364 ( 
.A1(n_347),
.A2(n_336),
.B1(n_334),
.B2(n_331),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_370),
.B1(n_380),
.B2(n_125),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_360),
.A2(n_130),
.B(n_106),
.Y(n_365)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_132),
.A3(n_135),
.B1(n_140),
.B2(n_130),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_378),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_354),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_376),
.B(n_379),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_59),
.C(n_84),
.Y(n_377)
);

BUFx12_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_125),
.B(n_120),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_375),
.B(n_369),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_382),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_384),
.B(n_391),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_373),
.B(n_352),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_387),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_371),
.C(n_372),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_351),
.C(n_342),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_339),
.C(n_83),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_55),
.C(n_69),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_395),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_21),
.C(n_33),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_397),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_30),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_377),
.B(n_36),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_399),
.Y(n_407)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_402),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_393),
.A2(n_364),
.B(n_381),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_401),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_394),
.Y(n_402)
);

AOI31xp33_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_378),
.A3(n_382),
.B(n_368),
.Y(n_404)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_406),
.C(n_28),
.Y(n_423)
);

AOI21x1_ASAP7_75t_SL g406 ( 
.A1(n_398),
.A2(n_382),
.B(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_408),
.B(n_411),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_29),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_384),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_414),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_389),
.C(n_392),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_409),
.A2(n_390),
.B1(n_383),
.B2(n_21),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_420),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_403),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_27),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g417 ( 
.A1(n_406),
.A2(n_29),
.B(n_2),
.C(n_3),
.Y(n_417)
);

AOI31xp67_ASAP7_75t_L g432 ( 
.A1(n_417),
.A2(n_1),
.A3(n_3),
.B(n_4),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_405),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_41),
.C(n_28),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_1),
.B(n_2),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_411),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_26),
.Y(n_429)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_423),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_418),
.A2(n_27),
.B(n_2),
.Y(n_425)
);

O2A1O1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_425),
.A2(n_431),
.B(n_432),
.C(n_417),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_429),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_27),
.C(n_60),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_428),
.B(n_430),
.Y(n_436)
);

AOI211x1_ASAP7_75t_L g434 ( 
.A1(n_419),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_434)
);

XNOR2x2_ASAP7_75t_SL g441 ( 
.A(n_434),
.B(n_428),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_424),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g445 ( 
.A(n_435),
.B(n_439),
.CI(n_440),
.CON(n_445),
.SN(n_445)
);

AOI332xp33_ASAP7_75t_L g444 ( 
.A1(n_438),
.A2(n_441),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.B3(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_417),
.B(n_6),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_26),
.C(n_7),
.Y(n_440)
);

AOI322xp5_ASAP7_75t_L g442 ( 
.A1(n_436),
.A2(n_26),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_5),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_443),
.Y(n_448)
);

AOI322xp5_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_26),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_12),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_11),
.C(n_13),
.Y(n_447)
);

AOI321xp33_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_26),
.C(n_418),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_SL g449 ( 
.A(n_446),
.B(n_447),
.C(n_14),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_448),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_14),
.Y(n_452)
);


endmodule