module fake_jpeg_27511_n_30 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_4),
.B1(n_10),
.B2(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AOI21x1_ASAP7_75t_SL g25 ( 
.A1(n_24),
.A2(n_18),
.B(n_17),
.Y(n_25)
);

OAI322xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_24),
.A3(n_22),
.B1(n_17),
.B2(n_14),
.C1(n_1),
.C2(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_26),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_0),
.B(n_11),
.Y(n_30)
);


endmodule