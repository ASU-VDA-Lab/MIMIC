module fake_netlist_1_6909_n_886 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_886);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_886;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_163;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_59), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_52), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_64), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_38), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_99), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_10), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_49), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_29), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_46), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_83), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_1), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_71), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_54), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_44), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_65), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_57), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_19), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_40), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_101), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_33), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_37), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_1), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_21), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_24), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_2), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_17), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_19), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_105), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_70), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_86), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_109), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_43), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_45), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_68), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_45), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_123), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_123), .B(n_0), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_134), .B(n_0), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_134), .B(n_3), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_154), .B(n_3), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_143), .B(n_4), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
NOR2xp67_ASAP7_75t_L g170 ( .A(n_118), .B(n_50), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_114), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_120), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_159), .A2(n_133), .B1(n_116), .B2(n_143), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_171), .B(n_144), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_156), .B(n_118), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_159), .A2(n_133), .B1(n_144), .B2(n_154), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g184 ( .A1(n_176), .A2(n_142), .B1(n_127), .B2(n_152), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_176), .A2(n_137), .B1(n_122), .B2(n_151), .Y(n_185) );
OAI22xp33_ASAP7_75t_SL g186 ( .A1(n_171), .A2(n_138), .B1(n_124), .B2(n_125), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
OA22x2_ASAP7_75t_L g188 ( .A1(n_156), .A2(n_154), .B1(n_130), .B2(n_139), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_171), .B(n_141), .Y(n_189) );
AO22x2_ASAP7_75t_L g190 ( .A1(n_158), .A2(n_115), .B1(n_117), .B2(n_119), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_171), .B(n_145), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_159), .A2(n_146), .B1(n_119), .B2(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
AO22x2_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_164), .B1(n_161), .B2(n_172), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_156), .B(n_111), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_158), .B(n_117), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_161), .B(n_112), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g200 ( .A1(n_160), .A2(n_135), .B1(n_140), .B2(n_153), .Y(n_200) );
NAND2xp33_ASAP7_75t_SL g201 ( .A(n_158), .B(n_140), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_164), .A2(n_150), .B1(n_149), .B2(n_148), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_164), .A2(n_147), .B1(n_136), .B2(n_131), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_164), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_160), .A2(n_129), .B1(n_128), .B2(n_126), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_155), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_161), .B(n_113), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_155), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_161), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_172), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_214) );
OR2x6_ASAP7_75t_L g215 ( .A(n_165), .B(n_11), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_161), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_216) );
AOI22x1_ASAP7_75t_SL g217 ( .A1(n_172), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_165), .B(n_15), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_170), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_174), .B(n_18), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_170), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_162), .B(n_20), .Y(n_226) );
OAI22xp33_ASAP7_75t_SL g227 ( .A1(n_174), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_227) );
AO22x2_ASAP7_75t_L g228 ( .A1(n_174), .A2(n_23), .B1(n_25), .B2(n_26), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_180), .B(n_170), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
INVx4_ASAP7_75t_SL g232 ( .A(n_226), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_180), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_194), .B(n_162), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_200), .B(n_205), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_198), .B(n_162), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_180), .B(n_25), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_197), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_184), .Y(n_246) );
XNOR2xp5_ASAP7_75t_L g247 ( .A(n_179), .B(n_26), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_181), .B(n_166), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_198), .B(n_166), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_185), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_190), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_190), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_193), .B(n_27), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_220), .B(n_166), .Y(n_256) );
XNOR2xp5_ASAP7_75t_L g257 ( .A(n_179), .B(n_27), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_195), .B(n_166), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_182), .B(n_28), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_199), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_189), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_181), .B(n_166), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_207), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_215), .B(n_28), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_191), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_213), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_202), .B(n_51), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_213), .Y(n_270) );
XOR2xp5_ASAP7_75t_L g271 ( .A(n_182), .B(n_29), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_215), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_203), .B(n_53), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_213), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_225), .B(n_55), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_208), .A2(n_174), .B(n_173), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_215), .B(n_30), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_216), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_188), .B(n_30), .Y(n_279) );
INVxp67_ASAP7_75t_SL g280 ( .A(n_200), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_192), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_216), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_188), .B(n_31), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_183), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_204), .Y(n_285) );
XNOR2x2_ASAP7_75t_L g286 ( .A(n_228), .B(n_174), .Y(n_286) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_205), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_223), .B(n_173), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_183), .Y(n_291) );
XOR2x2_ASAP7_75t_L g292 ( .A(n_186), .B(n_31), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
AND3x1_ASAP7_75t_SL g295 ( .A(n_292), .B(n_217), .C(n_204), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_261), .B(n_201), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_234), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_261), .B(n_201), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_280), .B(n_212), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_238), .B(n_212), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_238), .B(n_214), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_234), .B(n_204), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_239), .B(n_218), .Y(n_305) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_242), .A2(n_227), .B(n_221), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_290), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_243), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_230), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_287), .B(n_221), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_236), .B(n_183), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_243), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_239), .B(n_228), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_250), .B(n_32), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_231), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_266), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_231), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_230), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_262), .A2(n_173), .B(n_228), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_236), .B(n_224), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_237), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_262), .B(n_173), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_265), .A2(n_173), .B(n_224), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_265), .B(n_173), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_266), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_235), .B(n_32), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_255), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_250), .B(n_34), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_229), .B(n_34), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_241), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_235), .B(n_35), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_237), .B(n_173), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_229), .B(n_35), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_251), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_241), .A2(n_224), .B(n_178), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_241), .A2(n_224), .B(n_178), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_251), .B(n_36), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_245), .B(n_178), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_36), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_253), .B(n_178), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_254), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_255), .B(n_178), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_254), .B(n_37), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_240), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_245), .B(n_178), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_318), .B(n_277), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_311), .B(n_293), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_297), .B(n_318), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_327), .B(n_277), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_327), .B(n_255), .Y(n_354) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_297), .B(n_268), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_338), .Y(n_357) );
NOR2xp33_ASAP7_75t_SL g358 ( .A(n_297), .B(n_268), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_297), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_309), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_311), .B(n_293), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_303), .B(n_263), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_297), .B(n_255), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_344), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_303), .B(n_294), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_328), .B(n_294), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_297), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_302), .B(n_270), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_305), .B(n_285), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_305), .B(n_240), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_348), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_329), .B(n_232), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_302), .B(n_270), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_305), .B(n_260), .Y(n_378) );
AND2x6_ASAP7_75t_L g379 ( .A(n_328), .B(n_274), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_309), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_329), .B(n_232), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_374), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_365), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_365), .B(n_338), .Y(n_386) );
INVx4_ASAP7_75t_L g387 ( .A(n_379), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_365), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_368), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_365), .B(n_321), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_363), .A2(n_295), .B1(n_271), .B2(n_304), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
BUFx2_ASAP7_75t_R g394 ( .A(n_374), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_365), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_365), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_368), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_363), .A2(n_304), .B1(n_271), .B2(n_260), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_363), .A2(n_295), .B1(n_304), .B2(n_314), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_360), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_365), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_360), .Y(n_406) );
BUFx12f_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
CKINVDCx11_ASAP7_75t_R g408 ( .A(n_375), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_368), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_378), .B(n_301), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_365), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_403), .Y(n_414) );
INVx6_ASAP7_75t_L g415 ( .A(n_407), .Y(n_415) );
BUFx10_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_392), .A2(n_378), .B1(n_292), .B2(n_229), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_384), .Y(n_419) );
INVx6_ASAP7_75t_L g420 ( .A(n_407), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_384), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_396), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_392), .A2(n_378), .B1(n_229), .B2(n_373), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_402), .B(n_378), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_396), .Y(n_425) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_408), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_392), .A2(n_378), .B1(n_373), .B2(n_272), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_399), .A2(n_321), .B1(n_354), .B2(n_373), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_396), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_412), .B(n_366), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_394), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_394), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_400), .A2(n_355), .B1(n_358), .B2(n_354), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_397), .A2(n_367), .B1(n_379), .B2(n_286), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_394), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_397), .A2(n_367), .B1(n_379), .B2(n_286), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_391), .A2(n_301), .B(n_306), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_407), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_400), .A2(n_399), .B1(n_412), .B2(n_373), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_404), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_400), .A2(n_373), .B1(n_372), .B2(n_367), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_412), .B(n_366), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_387), .A2(n_348), .B1(n_299), .B2(n_358), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_397), .A2(n_372), .B1(n_367), .B2(n_247), .Y(n_456) );
INVx8_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_407), .A2(n_367), .B1(n_379), .B2(n_354), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_411), .B(n_366), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_458), .A2(n_257), .B(n_247), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_417), .A2(n_314), .B1(n_372), .B2(n_387), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_439), .B(n_413), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_444), .A2(n_387), .B1(n_389), .B2(n_409), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_423), .A2(n_314), .B1(n_372), .B2(n_387), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_457), .A2(n_387), .B1(n_398), .B2(n_409), .Y(n_465) );
OAI21xp5_ASAP7_75t_SL g466 ( .A1(n_438), .A2(n_383), .B(n_375), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_437), .A2(n_372), .B1(n_387), .B2(n_367), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_439), .B(n_404), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_416), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_439), .B(n_410), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_424), .B(n_351), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_437), .A2(n_367), .B1(n_379), .B2(n_408), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_449), .A2(n_367), .B1(n_379), .B2(n_409), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_428), .A2(n_367), .B1(n_379), .B2(n_409), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_442), .B(n_410), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_428), .A2(n_367), .B1(n_379), .B2(n_389), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_427), .A2(n_367), .B1(n_379), .B2(n_389), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_443), .A2(n_306), .B(n_332), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_447), .A2(n_367), .B1(n_379), .B2(n_398), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_438), .A2(n_367), .B1(n_379), .B2(n_398), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_442), .B(n_410), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_424), .B(n_351), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_441), .A2(n_383), .B(n_375), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_419), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_442), .B(n_410), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_456), .A2(n_354), .B1(n_328), .B2(n_389), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_441), .A2(n_383), .B(n_375), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_430), .B(n_351), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g492 ( .A1(n_444), .A2(n_246), .B1(n_281), .B2(n_267), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_414), .A2(n_283), .B(n_279), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_434), .Y(n_494) );
OAI22x1_ASAP7_75t_SL g495 ( .A1(n_431), .A2(n_252), .B1(n_398), .B2(n_411), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_414), .A2(n_283), .B(n_279), .Y(n_496) );
OAI22xp33_ASAP7_75t_SL g497 ( .A1(n_415), .A2(n_386), .B1(n_410), .B2(n_395), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_457), .A2(n_367), .B1(n_379), .B2(n_336), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_416), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_457), .A2(n_367), .B1(n_379), .B2(n_336), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_421), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_457), .A2(n_379), .B1(n_332), .B2(n_353), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_415), .A2(n_328), .B1(n_353), .B2(n_350), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_416), .Y(n_505) );
INVx5_ASAP7_75t_SL g506 ( .A(n_435), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_434), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_457), .A2(n_379), .B1(n_328), .B2(n_353), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_415), .A2(n_328), .B1(n_353), .B2(n_350), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_454), .A2(n_383), .B(n_375), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_436), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_415), .A2(n_350), .B1(n_353), .B2(n_352), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_415), .A2(n_350), .B1(n_352), .B2(n_386), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_430), .B(n_362), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g515 ( .A1(n_426), .A2(n_298), .B1(n_350), .B2(n_331), .C1(n_316), .C2(n_362), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_457), .A2(n_358), .B1(n_355), .B2(n_299), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_426), .A2(n_379), .B1(n_368), .B2(n_352), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_426), .A2(n_355), .B1(n_370), .B2(n_368), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_416), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_420), .A2(n_352), .B1(n_386), .B2(n_364), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_418), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_448), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_418), .B(n_405), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_436), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_448), .B(n_385), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_420), .A2(n_401), .B1(n_390), .B2(n_386), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_420), .A2(n_370), .B1(n_368), .B2(n_359), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_420), .A2(n_352), .B1(n_369), .B2(n_375), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_453), .B(n_362), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_448), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_432), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_420), .A2(n_352), .B1(n_386), .B2(n_364), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_452), .B(n_385), .Y(n_533) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_453), .A2(n_383), .B(n_375), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g535 ( .A1(n_492), .A2(n_440), .B1(n_446), .B2(n_450), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_521), .B(n_446), .Y(n_536) );
AOI21xp5_ASAP7_75t_SL g537 ( .A1(n_500), .A2(n_459), .B(n_450), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_534), .A2(n_459), .B1(n_386), .B2(n_452), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_515), .A2(n_383), .B1(n_352), .B2(n_289), .Y(n_539) );
OAI222xp33_ASAP7_75t_L g540 ( .A1(n_513), .A2(n_455), .B1(n_445), .B2(n_425), .C1(n_422), .C2(n_452), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_467), .A2(n_383), .B1(n_289), .B2(n_369), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_500), .A2(n_445), .B1(n_455), .B2(n_425), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_472), .A2(n_289), .B1(n_369), .B2(n_364), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_460), .B(n_435), .C(n_393), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_512), .A2(n_369), .B1(n_364), .B2(n_341), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_476), .A2(n_369), .B1(n_364), .B2(n_341), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_534), .A2(n_422), .B1(n_388), .B2(n_405), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_478), .A2(n_341), .B1(n_343), .B2(n_347), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_489), .A2(n_347), .B1(n_343), .B2(n_334), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_483), .A2(n_347), .B1(n_343), .B2(n_334), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_492), .A2(n_405), .B1(n_388), .B2(n_393), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_482), .A2(n_334), .B1(n_391), .B2(n_370), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_479), .A2(n_370), .B1(n_435), .B2(n_371), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_508), .A2(n_435), .B1(n_371), .B2(n_376), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_473), .B(n_475), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_504), .A2(n_435), .B1(n_371), .B2(n_376), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_497), .B(n_388), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_509), .A2(n_435), .B1(n_376), .B2(n_359), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_466), .A2(n_388), .B1(n_405), .B2(n_393), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_475), .B(n_451), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_461), .A2(n_359), .B1(n_401), .B2(n_390), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_519), .A2(n_390), .B1(n_401), .B2(n_451), .Y(n_564) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_520), .A2(n_451), .B1(n_395), .B2(n_385), .C1(n_390), .C2(n_401), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_474), .A2(n_401), .B1(n_390), .B2(n_451), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_460), .A2(n_269), .B1(n_273), .B2(n_298), .C(n_316), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_464), .A2(n_331), .B1(n_382), .B2(n_381), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_382), .B1(n_381), .B2(n_357), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_495), .A2(n_300), .B1(n_337), .B2(n_326), .C(n_324), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_532), .A2(n_382), .B1(n_381), .B2(n_357), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_486), .A2(n_490), .B1(n_510), .B2(n_469), .Y(n_572) );
OAI222xp33_ASAP7_75t_L g573 ( .A1(n_469), .A2(n_385), .B1(n_395), .B2(n_278), .C1(n_282), .C2(n_288), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_481), .A2(n_382), .B1(n_381), .B2(n_357), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_499), .A2(n_382), .B1(n_357), .B2(n_274), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_501), .A2(n_382), .B1(n_395), .B2(n_385), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_526), .B(n_490), .C(n_486), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_494), .B(n_385), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_517), .A2(n_382), .B1(n_395), .B2(n_393), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_510), .A2(n_395), .B(n_380), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_465), .A2(n_405), .B1(n_393), .B2(n_388), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_494), .B(n_388), .Y(n_582) );
AOI221xp5_ASAP7_75t_SL g583 ( .A1(n_497), .A2(n_337), .B1(n_377), .B2(n_356), .C(n_300), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_528), .A2(n_405), .B1(n_393), .B2(n_388), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_527), .A2(n_382), .B1(n_393), .B2(n_388), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_493), .A2(n_405), .B1(n_393), .B2(n_319), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_493), .A2(n_405), .B1(n_393), .B2(n_319), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_496), .A2(n_405), .B1(n_393), .B2(n_319), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_496), .A2(n_405), .B1(n_319), .B2(n_345), .Y(n_590) );
OAI22xp33_ASAP7_75t_SL g591 ( .A1(n_505), .A2(n_346), .B1(n_361), .B2(n_380), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_471), .A2(n_345), .B1(n_346), .B2(n_356), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g593 ( .A1(n_505), .A2(n_380), .B1(n_361), .B2(n_377), .C1(n_356), .C2(n_349), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_485), .A2(n_345), .B1(n_377), .B2(n_296), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_505), .A2(n_365), .B(n_361), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_518), .A2(n_308), .B1(n_313), .B2(n_296), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_516), .A2(n_308), .B1(n_313), .B2(n_296), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_463), .A2(n_380), .B1(n_361), .B2(n_349), .C1(n_342), .C2(n_323), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_491), .A2(n_308), .B1(n_313), .B2(n_232), .Y(n_599) );
NAND2xp33_ASAP7_75t_R g600 ( .A(n_502), .B(n_38), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_514), .A2(n_232), .B1(n_317), .B2(n_380), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_495), .A2(n_317), .B1(n_323), .B2(n_320), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_529), .A2(n_232), .B1(n_317), .B2(n_342), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_507), .B(n_39), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_511), .B(n_39), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_511), .A2(n_323), .B1(n_259), .B2(n_275), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_524), .B(n_157), .C(n_163), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_524), .A2(n_259), .B1(n_324), .B2(n_326), .Y(n_608) );
AOI222xp33_ASAP7_75t_L g609 ( .A1(n_487), .A2(n_40), .B1(n_41), .B2(n_42), .C1(n_44), .C2(n_46), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_480), .A2(n_259), .B1(n_333), .B2(n_309), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_480), .A2(n_259), .B1(n_333), .B2(n_310), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_468), .B(n_41), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_462), .B(n_157), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g615 ( .A1(n_487), .A2(n_42), .B1(n_47), .B2(n_48), .C1(n_310), .C2(n_320), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_523), .A2(n_344), .B1(n_333), .B2(n_310), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_498), .A2(n_310), .B1(n_320), .B2(n_333), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_498), .A2(n_320), .B1(n_344), .B2(n_312), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_468), .B(n_47), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_506), .A2(n_344), .B1(n_264), .B2(n_325), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_502), .A2(n_344), .B1(n_335), .B2(n_325), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_525), .A2(n_312), .B1(n_322), .B2(n_167), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_462), .B(n_169), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_506), .A2(n_177), .B1(n_163), .B2(n_167), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_523), .B(n_157), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_530), .A2(n_335), .B1(n_248), .B2(n_322), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_525), .A2(n_157), .B1(n_163), .B2(n_167), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_533), .A2(n_157), .B1(n_163), .B2(n_167), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_470), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_531), .A2(n_178), .B1(n_163), .B2(n_167), .C1(n_168), .C2(n_169), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_530), .A2(n_340), .B1(n_339), .B2(n_249), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_533), .A2(n_157), .B1(n_163), .B2(n_167), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_477), .B(n_276), .C(n_249), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_477), .A2(n_157), .B1(n_163), .B2(n_178), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_583), .B(n_488), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_629), .B(n_488), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_577), .A2(n_484), .B(n_178), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_535), .B(n_484), .C(n_340), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_536), .B(n_506), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_554), .B(n_506), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_577), .A2(n_177), .B1(n_163), .B2(n_167), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_572), .A2(n_175), .B(n_163), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_535), .A2(n_177), .B1(n_163), .B2(n_167), .C(n_168), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_602), .A2(n_175), .B(n_163), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_600), .B(n_56), .Y(n_645) );
NOR3xp33_ASAP7_75t_SL g646 ( .A(n_570), .B(n_258), .C(n_339), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_551), .B(n_58), .C(n_61), .Y(n_647) );
OA21x2_ASAP7_75t_L g648 ( .A1(n_583), .A2(n_244), .B(n_284), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_604), .B(n_244), .C(n_256), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_602), .A2(n_175), .B1(n_163), .B2(n_167), .C(n_168), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_609), .A2(n_177), .B1(n_167), .B2(n_168), .C(n_169), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_595), .A2(n_169), .B(n_167), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_544), .A2(n_175), .B1(n_167), .B2(n_168), .Y(n_653) );
OAI22xp33_ASAP7_75t_SL g654 ( .A1(n_538), .A2(n_62), .B1(n_63), .B2(n_66), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_609), .A2(n_177), .B1(n_168), .B2(n_169), .C(n_175), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_538), .B(n_177), .Y(n_656) );
AOI221xp5_ASAP7_75t_SL g657 ( .A1(n_551), .A2(n_177), .B1(n_175), .B2(n_169), .C(n_168), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_595), .B(n_556), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_630), .B(n_177), .C(n_168), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_614), .B(n_177), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_611), .B(n_177), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_584), .B(n_175), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_591), .B(n_175), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_591), .B(n_175), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_544), .A2(n_157), .B1(n_168), .B2(n_169), .C(n_175), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_615), .A2(n_175), .B(n_169), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_580), .A2(n_169), .B(n_168), .Y(n_667) );
OAI221xp5_ASAP7_75t_SL g668 ( .A1(n_580), .A2(n_169), .B1(n_168), .B2(n_157), .C(n_74), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_584), .B(n_623), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_547), .B(n_168), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_562), .B(n_157), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_557), .B(n_67), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_630), .B(n_157), .C(n_307), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_547), .B(n_69), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_561), .B(n_72), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_561), .B(n_75), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_562), .B(n_77), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_582), .B(n_78), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_582), .B(n_79), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_605), .A2(n_80), .B(n_81), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_559), .B(n_85), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_539), .A2(n_330), .B1(n_307), .B2(n_88), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_578), .B(n_87), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_537), .A2(n_330), .B(n_307), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_581), .B(n_89), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_581), .B(n_90), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_537), .B(n_307), .C(n_330), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_585), .B(n_92), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_585), .B(n_564), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_613), .B(n_93), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_542), .B(n_94), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_555), .A2(n_330), .B1(n_307), .B2(n_97), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_619), .Y(n_693) );
AND4x1_ASAP7_75t_L g694 ( .A(n_596), .B(n_95), .C(n_96), .D(n_98), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_567), .B(n_100), .Y(n_695) );
AOI21xp5_ASAP7_75t_SL g696 ( .A1(n_616), .A2(n_330), .B(n_307), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_616), .B(n_102), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_558), .B(n_103), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_597), .B(n_104), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_543), .A2(n_330), .B1(n_290), .B2(n_284), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_560), .B(n_571), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_607), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_625), .B(n_586), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_607), .B(n_290), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_579), .B(n_290), .C(n_291), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_627), .B(n_106), .C(n_107), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_617), .B(n_108), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_540), .A2(n_110), .B1(n_593), .B2(n_594), .C(n_568), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_566), .B(n_563), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_574), .B(n_545), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_598), .B(n_621), .C(n_626), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_576), .B(n_552), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_628), .B(n_632), .C(n_624), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_634), .B(n_633), .C(n_610), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_573), .B(n_565), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_626), .B(n_620), .C(n_631), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_541), .B(n_589), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_549), .B(n_553), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_612), .B(n_588), .C(n_587), .Y(n_719) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_569), .A2(n_546), .B1(n_550), .B2(n_575), .C(n_548), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_592), .B(n_590), .Y(n_721) );
NAND2xp33_ASAP7_75t_SL g722 ( .A(n_599), .B(n_618), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_601), .B(n_603), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_608), .A2(n_606), .B(n_622), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_631), .B(n_630), .C(n_609), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_630), .B(n_609), .C(n_583), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_577), .A2(n_572), .B1(n_544), .B2(n_539), .Y(n_727) );
AOI21xp5_ASAP7_75t_SL g728 ( .A1(n_538), .A2(n_580), .B(n_577), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_629), .B(n_554), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_629), .B(n_536), .Y(n_730) );
NAND4xp75_ASAP7_75t_L g731 ( .A(n_708), .B(n_657), .C(n_647), .D(n_691), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_727), .B(n_728), .C(n_726), .Y(n_732) );
NAND4xp75_ASAP7_75t_L g733 ( .A(n_691), .B(n_663), .C(n_664), .D(n_715), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_662), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_669), .B(n_689), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_725), .A2(n_722), .B1(n_711), .B2(n_709), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_693), .B(n_730), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_645), .A2(n_689), .B1(n_687), .B2(n_654), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_716), .B(n_637), .C(n_642), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_652), .B(n_722), .C(n_641), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_636), .B(n_656), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_635), .B(n_644), .C(n_719), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_635), .B(n_714), .C(n_638), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_656), .B(n_658), .Y(n_744) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_649), .B(n_665), .C(n_695), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_670), .B(n_640), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_643), .B(n_655), .C(n_651), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_709), .B(n_717), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_671), .Y(n_749) );
NAND2xp33_ASAP7_75t_L g750 ( .A(n_684), .B(n_697), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_670), .B(n_674), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_718), .B(n_720), .Y(n_752) );
INVx1_ASAP7_75t_SL g753 ( .A(n_639), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_662), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_685), .B(n_686), .Y(n_755) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_704), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_712), .A2(n_710), .B1(n_666), .B2(n_723), .Y(n_757) );
CKINVDCx14_ASAP7_75t_R g758 ( .A(n_697), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_667), .B(n_724), .C(n_659), .Y(n_759) );
AOI211xp5_ASAP7_75t_L g760 ( .A1(n_696), .A2(n_673), .B(n_712), .C(n_668), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_710), .A2(n_721), .B1(n_713), .B2(n_701), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_650), .B(n_680), .C(n_690), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_702), .B(n_676), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_685), .A2(n_686), .B1(n_703), .B2(n_676), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_675), .B(n_702), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_661), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_660), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_677), .B(n_681), .Y(n_768) );
NAND4xp75_ASAP7_75t_L g769 ( .A(n_648), .B(n_681), .C(n_688), .D(n_646), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_653), .B(n_688), .C(n_704), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_678), .Y(n_771) );
INVxp33_ASAP7_75t_L g772 ( .A(n_672), .Y(n_772) );
INVxp67_ASAP7_75t_L g773 ( .A(n_678), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_679), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_694), .B(n_679), .C(n_698), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_683), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_683), .B(n_698), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_705), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_700), .B(n_699), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_706), .B(n_692), .C(n_682), .Y(n_780) );
INVxp33_ASAP7_75t_L g781 ( .A(n_699), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_707), .B(n_726), .C(n_708), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_669), .B(n_729), .Y(n_783) );
OA211x2_ASAP7_75t_L g784 ( .A1(n_727), .A2(n_684), .B(n_580), .C(n_664), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_669), .B(n_729), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_725), .A2(n_577), .B1(n_726), .B2(n_572), .Y(n_786) );
INVx3_ASAP7_75t_SL g787 ( .A(n_691), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_730), .B(n_636), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_669), .B(n_729), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_727), .A2(n_572), .B1(n_577), .B2(n_535), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_693), .B(n_531), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_726), .B(n_708), .C(n_642), .Y(n_792) );
INVx2_ASAP7_75t_SL g793 ( .A(n_734), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_748), .B(n_735), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_788), .Y(n_795) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_787), .B(n_732), .Y(n_796) );
INVx1_ASAP7_75t_SL g797 ( .A(n_753), .Y(n_797) );
NAND4xp75_ASAP7_75t_L g798 ( .A(n_790), .B(n_784), .C(n_736), .D(n_752), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_788), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_783), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_734), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_786), .B(n_743), .C(n_761), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_759), .B(n_742), .C(n_792), .Y(n_803) );
NAND4xp75_ASAP7_75t_L g804 ( .A(n_765), .B(n_755), .C(n_791), .D(n_779), .Y(n_804) );
NAND4xp75_ASAP7_75t_L g805 ( .A(n_779), .B(n_744), .C(n_738), .D(n_787), .Y(n_805) );
NOR4xp25_ASAP7_75t_L g806 ( .A(n_757), .B(n_739), .C(n_740), .D(n_737), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_785), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_778), .B(n_756), .Y(n_808) );
NAND4xp75_ASAP7_75t_L g809 ( .A(n_777), .B(n_763), .C(n_776), .D(n_768), .Y(n_809) );
NAND4xp75_ASAP7_75t_SL g810 ( .A(n_733), .B(n_763), .C(n_731), .D(n_751), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_789), .Y(n_811) );
XNOR2x2_ASAP7_75t_L g812 ( .A(n_733), .B(n_769), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_741), .B(n_749), .Y(n_813) );
NOR2xp33_ASAP7_75t_SL g814 ( .A(n_775), .B(n_731), .Y(n_814) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_769), .B(n_778), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_754), .Y(n_816) );
XOR2x2_ASAP7_75t_L g817 ( .A(n_782), .B(n_764), .Y(n_817) );
XNOR2x2_ASAP7_75t_L g818 ( .A(n_770), .B(n_745), .Y(n_818) );
XOR2x2_ASAP7_75t_L g819 ( .A(n_758), .B(n_760), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_772), .B(n_781), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_746), .Y(n_821) );
INVx2_ASAP7_75t_SL g822 ( .A(n_793), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_800), .Y(n_823) );
AO22x2_ASAP7_75t_L g824 ( .A1(n_798), .A2(n_774), .B1(n_771), .B2(n_773), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_816), .B(n_766), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_797), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_807), .Y(n_827) );
XOR2xp5_ASAP7_75t_L g828 ( .A(n_798), .B(n_772), .Y(n_828) );
XOR2x2_ASAP7_75t_L g829 ( .A(n_819), .B(n_747), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_811), .Y(n_830) );
XOR2x2_ASAP7_75t_L g831 ( .A(n_817), .B(n_780), .Y(n_831) );
INVx1_ASAP7_75t_SL g832 ( .A(n_801), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_813), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_795), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_814), .A2(n_750), .B1(n_781), .B2(n_762), .Y(n_835) );
XOR2xp5_ASAP7_75t_L g836 ( .A(n_810), .B(n_767), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_799), .Y(n_837) );
INVxp67_ASAP7_75t_L g838 ( .A(n_802), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_825), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_833), .Y(n_840) );
OA22x2_ASAP7_75t_L g841 ( .A1(n_828), .A2(n_820), .B1(n_818), .B2(n_808), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_834), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_825), .Y(n_843) );
XNOR2xp5_ASAP7_75t_L g844 ( .A(n_829), .B(n_796), .Y(n_844) );
CKINVDCx16_ASAP7_75t_R g845 ( .A(n_826), .Y(n_845) );
AO22x1_ASAP7_75t_L g846 ( .A1(n_838), .A2(n_803), .B1(n_815), .B2(n_818), .Y(n_846) );
AOI22x1_ASAP7_75t_L g847 ( .A1(n_828), .A2(n_796), .B1(n_806), .B2(n_812), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_822), .Y(n_848) );
AO22x2_ASAP7_75t_L g849 ( .A1(n_832), .A2(n_805), .B1(n_808), .B2(n_804), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_837), .Y(n_850) );
AO22x2_ASAP7_75t_L g851 ( .A1(n_822), .A2(n_804), .B1(n_809), .B2(n_821), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_835), .B(n_794), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_840), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_845), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_848), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_842), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_850), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_839), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_839), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_843), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_843), .Y(n_861) );
AOI311xp33_ASAP7_75t_L g862 ( .A1(n_855), .A2(n_841), .A3(n_831), .B(n_844), .C(n_829), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_854), .Y(n_863) );
AOI22x1_ASAP7_75t_L g864 ( .A1(n_854), .A2(n_844), .B1(n_849), .B2(n_851), .Y(n_864) );
OA22x2_ASAP7_75t_L g865 ( .A1(n_853), .A2(n_847), .B1(n_841), .B2(n_846), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_858), .Y(n_866) );
OAI22xp5_ASAP7_75t_SL g867 ( .A1(n_863), .A2(n_836), .B1(n_841), .B2(n_847), .Y(n_867) );
AO22x1_ASAP7_75t_L g868 ( .A1(n_865), .A2(n_846), .B1(n_853), .B2(n_856), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_864), .Y(n_869) );
BUFx2_ASAP7_75t_L g870 ( .A(n_869), .Y(n_870) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_868), .B(n_866), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_867), .A2(n_865), .B1(n_831), .B2(n_849), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_872), .A2(n_849), .B1(n_851), .B2(n_824), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_870), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_874), .Y(n_875) );
AOI22xp5_ASAP7_75t_SL g876 ( .A1(n_873), .A2(n_862), .B1(n_864), .B2(n_836), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_876), .B(n_871), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_875), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_878), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_879), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_880), .A2(n_877), .B1(n_852), .B2(n_866), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_881), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_861), .B1(n_860), .B2(n_859), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_883), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_884), .A2(n_857), .B1(n_849), .B2(n_851), .C(n_824), .Y(n_885) );
AOI211xp5_ASAP7_75t_L g886 ( .A1(n_885), .A2(n_823), .B(n_827), .C(n_830), .Y(n_886) );
endmodule