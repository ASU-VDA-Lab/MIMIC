module fake_jpeg_11740_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVxp67_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.C(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_48),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

XNOR2x1_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_2),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_47),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.C(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_30),
.B(n_4),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_3),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_78),
.B1(n_79),
.B2(n_76),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_5),
.B(n_6),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_5),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_70),
.B1(n_77),
.B2(n_73),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.C(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_80),
.B(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_16),
.C(n_7),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_18),
.C(n_12),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_19),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_22),
.B(n_13),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_23),
.C(n_14),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_15),
.Y(n_91)
);


endmodule