module real_aes_11834_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_730;
wire n_1023;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_1710;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_0), .Y(n_1384) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_2), .Y(n_1214) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_3), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_4), .A2(n_284), .B1(n_1038), .B2(n_1358), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_4), .A2(n_284), .B1(n_1177), .B2(n_1183), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_5), .A2(n_259), .B1(n_566), .B2(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g587 ( .A(n_5), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_6), .A2(n_248), .B1(n_1268), .B2(n_1270), .Y(n_1267) );
INVx1_ASAP7_75t_L g1303 ( .A(n_6), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_7), .A2(n_75), .B1(n_568), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g786 ( .A(n_7), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g1400 ( .A(n_8), .Y(n_1400) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_9), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_9), .B(n_225), .Y(n_349) );
INVx1_ASAP7_75t_L g379 ( .A(n_9), .Y(n_379) );
AND2x2_ASAP7_75t_L g383 ( .A(n_9), .B(n_378), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g1335 ( .A(n_10), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_11), .A2(n_180), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
INVx1_ASAP7_75t_L g1203 ( .A(n_11), .Y(n_1203) );
INVx1_ASAP7_75t_L g957 ( .A(n_12), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_12), .A2(n_163), .B1(n_992), .B2(n_995), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_13), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_14), .Y(n_1399) );
INVx1_ASAP7_75t_L g514 ( .A(n_15), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_15), .A2(n_80), .B1(n_580), .B2(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g1546 ( .A(n_16), .Y(n_1546) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_17), .Y(n_880) );
CKINVDCx16_ASAP7_75t_R g1472 ( .A(n_18), .Y(n_1472) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_19), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_19), .A2(n_271), .B1(n_980), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1078 ( .A(n_20), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_20), .A2(n_223), .B1(n_570), .B2(n_887), .Y(n_1096) );
AO221x2_ASAP7_75t_L g1451 ( .A1(n_21), .A2(n_64), .B1(n_1423), .B2(n_1430), .C(n_1452), .Y(n_1451) );
XNOR2xp5_ASAP7_75t_L g1666 ( .A(n_21), .B(n_1667), .Y(n_1666) );
AOI22xp33_ASAP7_75t_L g1706 ( .A1(n_21), .A2(n_1707), .B1(n_1711), .B2(n_1716), .Y(n_1706) );
INVx1_ASAP7_75t_L g1441 ( .A(n_22), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_23), .A2(n_53), .B1(n_1020), .B2(n_1022), .Y(n_1279) );
INVx1_ASAP7_75t_L g1315 ( .A(n_23), .Y(n_1315) );
INVx2_ASAP7_75t_L g335 ( .A(n_24), .Y(n_335) );
OR2x2_ASAP7_75t_L g453 ( .A(n_24), .B(n_333), .Y(n_453) );
INVx1_ASAP7_75t_L g1453 ( .A(n_25), .Y(n_1453) );
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_26), .A2(n_89), .B1(n_966), .B2(n_971), .Y(n_970) );
INVxp33_ASAP7_75t_L g1000 ( .A(n_26), .Y(n_1000) );
INVx1_ASAP7_75t_L g1227 ( .A(n_27), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_27), .A2(n_197), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_28), .A2(n_117), .B1(n_537), .B2(n_539), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_28), .A2(n_117), .B1(n_559), .B2(n_561), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_29), .A2(n_96), .B1(n_374), .B2(n_861), .C(n_862), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_29), .A2(n_172), .B1(n_457), .B2(n_870), .Y(n_928) );
BUFx2_ASAP7_75t_L g329 ( .A(n_30), .Y(n_329) );
BUFx2_ASAP7_75t_L g344 ( .A(n_30), .Y(n_344) );
INVx1_ASAP7_75t_L g454 ( .A(n_30), .Y(n_454) );
OR2x2_ASAP7_75t_L g750 ( .A(n_30), .B(n_349), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_31), .A2(n_219), .B1(n_542), .B2(n_1036), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_31), .A2(n_219), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_32), .Y(n_1172) );
INVx1_ASAP7_75t_L g1216 ( .A(n_33), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_33), .A2(n_168), .B1(n_571), .B2(n_1043), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_34), .Y(n_743) );
INVx1_ASAP7_75t_L g952 ( .A(n_35), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_35), .A2(n_71), .B1(n_434), .B2(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g1544 ( .A(n_36), .Y(n_1544) );
INVx1_ASAP7_75t_L g1678 ( .A(n_37), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1684 ( .A1(n_37), .A2(n_220), .B1(n_966), .B2(n_1036), .Y(n_1684) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_38), .A2(n_122), .B1(n_673), .B2(n_1066), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1394 ( .A1(n_38), .A2(n_122), .B1(n_404), .B2(n_406), .C(n_762), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_39), .A2(n_111), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g794 ( .A(n_39), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g1027 ( .A1(n_40), .A2(n_67), .B1(n_311), .B2(n_596), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_40), .A2(n_195), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
INVx1_ASAP7_75t_L g894 ( .A(n_41), .Y(n_894) );
OAI211xp5_ASAP7_75t_SL g916 ( .A1(n_41), .A2(n_612), .B(n_917), .C(n_924), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_42), .Y(n_1131) );
CKINVDCx16_ASAP7_75t_R g1431 ( .A(n_43), .Y(n_1431) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_44), .Y(n_1385) );
INVx1_ASAP7_75t_L g1540 ( .A(n_45), .Y(n_1540) );
INVx1_ASAP7_75t_L g655 ( .A(n_46), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_46), .A2(n_61), .B1(n_673), .B2(n_675), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g1681 ( .A1(n_47), .A2(n_249), .B1(n_673), .B2(n_1363), .Y(n_1681) );
AOI22xp33_ASAP7_75t_SL g1688 ( .A1(n_47), .A2(n_249), .B1(n_861), .B2(n_1352), .Y(n_1688) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_48), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g1382 ( .A1(n_49), .A2(n_55), .B1(n_468), .B2(n_684), .Y(n_1382) );
INVx1_ASAP7_75t_L g1390 ( .A(n_49), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_50), .A2(n_292), .B1(n_542), .B2(n_543), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_50), .A2(n_292), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
INVx1_ASAP7_75t_L g526 ( .A(n_51), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_51), .A2(n_270), .B1(n_547), .B2(n_550), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_52), .A2(n_87), .B1(n_966), .B2(n_968), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g979 ( .A1(n_52), .A2(n_87), .B1(n_684), .B2(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g1274 ( .A(n_53), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_54), .Y(n_1289) );
INVx1_ASAP7_75t_L g1389 ( .A(n_55), .Y(n_1389) );
INVx1_ASAP7_75t_L g1060 ( .A(n_56), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_56), .A2(n_170), .B1(n_547), .B2(n_550), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1712 ( .A1(n_57), .A2(n_1713), .B1(n_1714), .B2(n_1715), .Y(n_1712) );
CKINVDCx5p33_ASAP7_75t_R g1713 ( .A(n_57), .Y(n_1713) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_58), .A2(n_255), .B1(n_995), .B2(n_1069), .Y(n_1672) );
OAI22xp33_ASAP7_75t_L g1696 ( .A1(n_58), .A2(n_255), .B1(n_956), .B2(n_1076), .Y(n_1696) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_59), .A2(n_79), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_59), .A2(n_79), .B1(n_434), .B2(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g644 ( .A(n_60), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_60), .A2(n_188), .B1(n_667), .B2(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g652 ( .A(n_61), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_62), .A2(n_100), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g764 ( .A(n_62), .Y(n_764) );
INVx1_ASAP7_75t_L g1168 ( .A(n_63), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_63), .A2(n_65), .B1(n_374), .B2(n_1194), .C(n_1195), .Y(n_1193) );
INVx1_ASAP7_75t_L g1166 ( .A(n_65), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_66), .A2(n_104), .B1(n_861), .B2(n_974), .Y(n_973) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_66), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_67), .A2(n_247), .B1(n_1020), .B2(n_1022), .Y(n_1019) );
INVx1_ASAP7_75t_L g1065 ( .A(n_68), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_68), .A2(n_140), .B1(n_953), .B2(n_1088), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_69), .Y(n_837) );
AO22x2_ASAP7_75t_L g492 ( .A1(n_70), .A2(n_493), .B1(n_598), .B2(n_599), .Y(n_492) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_70), .Y(n_598) );
INVxp33_ASAP7_75t_L g948 ( .A(n_71), .Y(n_948) );
INVx1_ASAP7_75t_L g1464 ( .A(n_72), .Y(n_1464) );
CKINVDCx16_ASAP7_75t_R g1469 ( .A(n_73), .Y(n_1469) );
AO221x1_ASAP7_75t_L g1397 ( .A1(n_74), .A2(n_97), .B1(n_538), .B2(n_863), .C(n_975), .Y(n_1397) );
INVx1_ASAP7_75t_L g1408 ( .A(n_74), .Y(n_1408) );
INVx1_ASAP7_75t_L g795 ( .A(n_75), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_76), .A2(n_538), .B(n_863), .Y(n_1237) );
INVx1_ASAP7_75t_L g1240 ( .A(n_76), .Y(n_1240) );
INVx1_ASAP7_75t_L g1099 ( .A(n_77), .Y(n_1099) );
INVx1_ASAP7_75t_L g1342 ( .A(n_78), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_78), .A2(n_156), .B1(n_980), .B2(n_1183), .Y(n_1368) );
INVx1_ASAP7_75t_L g519 ( .A(n_80), .Y(n_519) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_81), .B(n_806), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_82), .A2(n_130), .B1(n_472), .B2(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g865 ( .A(n_82), .Y(n_865) );
INVx1_ASAP7_75t_L g1344 ( .A(n_83), .Y(n_1344) );
AOI22xp33_ASAP7_75t_SL g1366 ( .A1(n_83), .A2(n_230), .B1(n_1363), .B2(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1117 ( .A(n_84), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_84), .A2(n_114), .B1(n_566), .B2(n_568), .Y(n_1151) );
INVx1_ASAP7_75t_L g1488 ( .A(n_85), .Y(n_1488) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_86), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_88), .A2(n_293), .B1(n_570), .B2(n_887), .Y(n_886) );
INVxp67_ASAP7_75t_SL g914 ( .A(n_88), .Y(n_914) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_89), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_90), .A2(n_164), .B1(n_708), .B2(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g755 ( .A(n_90), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_91), .A2(n_146), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_91), .A2(n_146), .B1(n_1036), .B2(n_1038), .Y(n_1037) );
XNOR2x2_ASAP7_75t_L g1055 ( .A(n_92), .B(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1338 ( .A(n_93), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_93), .A2(n_149), .B1(n_966), .B2(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1014 ( .A(n_94), .Y(n_1014) );
OAI222xp33_ASAP7_75t_L g1025 ( .A1(n_94), .A2(n_195), .B1(n_209), .B2(n_582), .C1(n_850), .C2(n_1026), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_95), .A2(n_187), .B1(n_667), .B2(n_1183), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_95), .A2(n_187), .B1(n_609), .B2(n_610), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_96), .A2(n_148), .B1(n_872), .B2(n_874), .Y(n_929) );
INVx1_ASAP7_75t_L g1410 ( .A(n_97), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_98), .A2(n_119), .B1(n_367), .B2(n_369), .C(n_374), .Y(n_366) );
INVx1_ASAP7_75t_L g455 ( .A(n_98), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_99), .Y(n_1297) );
INVx1_ASAP7_75t_L g760 ( .A(n_100), .Y(n_760) );
AO22x2_ASAP7_75t_L g1324 ( .A1(n_101), .A2(n_1325), .B1(n_1326), .B2(n_1369), .Y(n_1324) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_101), .Y(n_1325) );
INVx1_ASAP7_75t_L g333 ( .A(n_102), .Y(n_333) );
INVx1_ASAP7_75t_L g424 ( .A(n_102), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_103), .Y(n_714) );
INVxp33_ASAP7_75t_L g997 ( .A(n_104), .Y(n_997) );
OAI222xp33_ASAP7_75t_L g1329 ( .A1(n_105), .A2(n_205), .B1(n_242), .B2(n_992), .C1(n_995), .C2(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1345 ( .A(n_105), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_106), .A2(n_127), .B1(n_1194), .B2(n_1195), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_106), .A2(n_127), .B1(n_673), .B2(n_1363), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_107), .A2(n_282), .B1(n_901), .B2(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g926 ( .A(n_107), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_108), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_109), .A2(n_184), .B1(n_1363), .B2(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1701 ( .A(n_109), .Y(n_1701) );
AOI22xp33_ASAP7_75t_SL g1682 ( .A1(n_110), .A2(n_159), .B1(n_667), .B2(n_1178), .Y(n_1682) );
AOI22xp33_ASAP7_75t_L g1687 ( .A1(n_110), .A2(n_159), .B1(n_920), .B2(n_1038), .Y(n_1687) );
INVx1_ASAP7_75t_L g788 ( .A(n_111), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_112), .A2(n_157), .B1(n_861), .B2(n_862), .C(n_863), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_112), .A2(n_192), .B1(n_872), .B2(n_874), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g1444 ( .A1(n_113), .A2(n_167), .B1(n_1445), .B2(n_1448), .Y(n_1444) );
INVx1_ASAP7_75t_L g1122 ( .A(n_114), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_115), .A2(n_264), .B1(n_1038), .B2(n_1234), .C(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1241 ( .A(n_115), .Y(n_1241) );
AOI22x1_ASAP7_75t_L g1371 ( .A1(n_116), .A2(n_1372), .B1(n_1373), .B2(n_1411), .Y(n_1371) );
INVxp67_ASAP7_75t_SL g1411 ( .A(n_116), .Y(n_1411) );
CKINVDCx5p33_ASAP7_75t_R g1295 ( .A(n_118), .Y(n_1295) );
INVx1_ASAP7_75t_L g463 ( .A(n_119), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_120), .A2(n_229), .B1(n_896), .B2(n_898), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_120), .A2(n_229), .B1(n_906), .B2(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g1334 ( .A(n_121), .Y(n_1334) );
AOI22xp33_ASAP7_75t_SL g1351 ( .A1(n_121), .A2(n_242), .B1(n_1195), .B2(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1438 ( .A(n_123), .Y(n_1438) );
INVx1_ASAP7_75t_L g1121 ( .A(n_124), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_124), .A2(n_252), .B1(n_426), .B2(n_1147), .C(n_1149), .Y(n_1146) );
INVx1_ASAP7_75t_L g877 ( .A(n_125), .Y(n_877) );
INVx1_ASAP7_75t_L g395 ( .A(n_126), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_126), .A2(n_261), .B1(n_426), .B2(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_128), .A2(n_243), .B1(n_356), .B2(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_128), .A2(n_243), .B1(n_426), .B2(n_429), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_129), .Y(n_633) );
INVx1_ASAP7_75t_L g866 ( .A(n_130), .Y(n_866) );
XOR2x2_ASAP7_75t_L g605 ( .A(n_131), .B(n_606), .Y(n_605) );
AO221x2_ASAP7_75t_L g1485 ( .A1(n_131), .A2(n_208), .B1(n_1430), .B2(n_1471), .C(n_1486), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_132), .A2(n_291), .B1(n_861), .B2(n_862), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_132), .A2(n_291), .B1(n_513), .B2(n_673), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_133), .B(n_1018), .Y(n_1278) );
INVx1_ASAP7_75t_L g1313 ( .A(n_133), .Y(n_1313) );
INVx1_ASAP7_75t_L g1670 ( .A(n_134), .Y(n_1670) );
AOI22xp33_ASAP7_75t_L g1685 ( .A1(n_134), .A2(n_218), .B1(n_405), .B2(n_861), .Y(n_1685) );
CKINVDCx5p33_ASAP7_75t_R g1173 ( .A(n_135), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_136), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_137), .A2(n_237), .B1(n_1183), .B2(n_1377), .Y(n_1376) );
AOI22xp33_ASAP7_75t_SL g1392 ( .A1(n_137), .A2(n_237), .B1(n_545), .B2(n_1393), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_138), .A2(n_266), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_138), .A2(n_266), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_139), .A2(n_206), .B1(n_1363), .B2(n_1380), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_139), .A2(n_612), .B1(n_1397), .B2(n_1398), .C(n_1401), .Y(n_1396) );
INVx1_ASAP7_75t_L g1059 ( .A(n_140), .Y(n_1059) );
INVx1_ASAP7_75t_L g302 ( .A(n_141), .Y(n_302) );
OA22x2_ASAP7_75t_L g1263 ( .A1(n_142), .A2(n_1264), .B1(n_1319), .B2(n_1320), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_142), .Y(n_1320) );
CKINVDCx5p33_ASAP7_75t_R g1232 ( .A(n_143), .Y(n_1232) );
CKINVDCx5p33_ASAP7_75t_R g1675 ( .A(n_144), .Y(n_1675) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_145), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g1223 ( .A1(n_147), .A2(n_404), .B(n_406), .Y(n_1223) );
INVx1_ASAP7_75t_L g1250 ( .A(n_147), .Y(n_1250) );
INVx1_ASAP7_75t_L g918 ( .A(n_148), .Y(n_918) );
INVx1_ASAP7_75t_L g1337 ( .A(n_149), .Y(n_1337) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_150), .Y(n_1130) );
XNOR2xp5_ASAP7_75t_L g1159 ( .A(n_151), .B(n_1160), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1450 ( .A1(n_151), .A2(n_201), .B1(n_1423), .B2(n_1430), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_152), .A2(n_245), .B1(n_356), .B2(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g466 ( .A(n_152), .Y(n_466) );
INVx1_ASAP7_75t_L g1074 ( .A(n_153), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_153), .A2(n_227), .B1(n_568), .B2(n_1011), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_154), .A2(n_272), .B1(n_561), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g594 ( .A(n_154), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_155), .Y(n_1213) );
INVx1_ASAP7_75t_L g1341 ( .A(n_156), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_157), .A2(n_222), .B1(n_457), .B2(n_870), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g1126 ( .A(n_158), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_160), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_161), .Y(n_631) );
INVx1_ASAP7_75t_L g1454 ( .A(n_162), .Y(n_1454) );
INVxp67_ASAP7_75t_SL g954 ( .A(n_163), .Y(n_954) );
INVx1_ASAP7_75t_L g767 ( .A(n_164), .Y(n_767) );
INVx1_ASAP7_75t_L g892 ( .A(n_165), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_165), .A2(n_639), .B1(n_909), .B2(n_912), .C(n_915), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_166), .A2(n_240), .B1(n_386), .B2(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g485 ( .A(n_166), .Y(n_485) );
INVx1_ASAP7_75t_L g1217 ( .A(n_168), .Y(n_1217) );
INVx1_ASAP7_75t_L g1104 ( .A(n_169), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_169), .A2(n_277), .B1(n_445), .B2(n_724), .Y(n_1141) );
INVx1_ASAP7_75t_L g1063 ( .A(n_170), .Y(n_1063) );
INVx1_ASAP7_75t_L g490 ( .A(n_171), .Y(n_490) );
INVx1_ASAP7_75t_L g922 ( .A(n_172), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_173), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1692 ( .A1(n_174), .A2(n_256), .B1(n_1183), .B2(n_1377), .Y(n_1692) );
INVx1_ASAP7_75t_L g1698 ( .A(n_174), .Y(n_1698) );
INVx1_ASAP7_75t_L g1029 ( .A(n_175), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_175), .A2(n_178), .B1(n_570), .B2(n_887), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_176), .A2(n_238), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_176), .A2(n_238), .B1(n_681), .B2(n_684), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_177), .A2(n_204), .B1(n_537), .B2(n_539), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1094 ( .A1(n_177), .A2(n_204), .B1(n_559), .B2(n_1011), .Y(n_1094) );
INVx1_ASAP7_75t_L g1030 ( .A(n_178), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_179), .Y(n_629) );
INVx1_ASAP7_75t_L g1204 ( .A(n_180), .Y(n_1204) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_181), .A2(n_190), .B1(n_1445), .B2(n_1448), .Y(n_1479) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_182), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_183), .A2(n_236), .B1(n_434), .B2(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1200 ( .A(n_183), .Y(n_1200) );
INVx1_ASAP7_75t_L g1695 ( .A(n_184), .Y(n_1695) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_185), .Y(n_1128) );
AOI22x1_ASAP7_75t_SL g1005 ( .A1(n_186), .A2(n_1006), .B1(n_1050), .B2(n_1051), .Y(n_1005) );
INVx1_ASAP7_75t_L g1050 ( .A(n_186), .Y(n_1050) );
INVx1_ASAP7_75t_L g648 ( .A(n_188), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_189), .Y(n_1169) );
INVx1_ASAP7_75t_L g695 ( .A(n_191), .Y(n_695) );
INVx1_ASAP7_75t_L g855 ( .A(n_192), .Y(n_855) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_193), .Y(n_304) );
AND3x2_ASAP7_75t_L g1424 ( .A(n_193), .B(n_302), .C(n_1425), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_193), .B(n_302), .Y(n_1435) );
INVx1_ASAP7_75t_L g1010 ( .A(n_194), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_194), .A2(n_247), .B1(n_537), .B2(n_1033), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g1480 ( .A1(n_196), .A2(n_233), .B1(n_1471), .B2(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1221 ( .A(n_197), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_198), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_199), .Y(n_1236) );
INVx2_ASAP7_75t_L g315 ( .A(n_200), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_202), .A2(n_411), .B1(n_639), .B2(n_640), .C(n_649), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_202), .A2(n_260), .B1(n_675), .B2(n_678), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_203), .Y(n_1229) );
INVx1_ASAP7_75t_L g1346 ( .A(n_205), .Y(n_1346) );
INVx1_ASAP7_75t_L g1395 ( .A(n_206), .Y(n_1395) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_207), .A2(n_216), .B1(n_1423), .B2(n_1430), .Y(n_1475) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_209), .Y(n_1013) );
INVx1_ASAP7_75t_L g1067 ( .A(n_210), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_210), .A2(n_239), .B1(n_580), .B2(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1425 ( .A(n_211), .Y(n_1425) );
INVx1_ASAP7_75t_L g885 ( .A(n_212), .Y(n_885) );
INVx1_ASAP7_75t_L g830 ( .A(n_213), .Y(n_830) );
OAI211xp5_ASAP7_75t_SL g852 ( .A1(n_213), .A2(n_612), .B(n_853), .C(n_864), .Y(n_852) );
CKINVDCx16_ASAP7_75t_R g937 ( .A(n_214), .Y(n_937) );
INVx1_ASAP7_75t_L g1185 ( .A(n_215), .Y(n_1185) );
INVx1_ASAP7_75t_L g1542 ( .A(n_217), .Y(n_1542) );
INVx1_ASAP7_75t_L g1674 ( .A(n_218), .Y(n_1674) );
INVx1_ASAP7_75t_L g1677 ( .A(n_220), .Y(n_1677) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_221), .A2(n_267), .B1(n_404), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_221), .A2(n_267), .B1(n_568), .B2(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g859 ( .A(n_222), .Y(n_859) );
INVx1_ASAP7_75t_L g1079 ( .A(n_223), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_224), .A2(n_231), .B1(n_770), .B2(n_774), .C(n_1112), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_224), .A2(n_231), .B1(n_719), .B2(n_1137), .C(n_1139), .Y(n_1136) );
INVx1_ASAP7_75t_L g317 ( .A(n_225), .Y(n_317) );
INVx2_ASAP7_75t_L g378 ( .A(n_225), .Y(n_378) );
INVx1_ASAP7_75t_L g826 ( .A(n_226), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_226), .A2(n_411), .B1(n_639), .B2(n_841), .C(n_849), .Y(n_840) );
INVx1_ASAP7_75t_L g1081 ( .A(n_227), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_228), .A2(n_295), .B1(n_570), .B2(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g844 ( .A(n_228), .Y(n_844) );
INVx1_ASAP7_75t_L g1348 ( .A(n_230), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g1474 ( .A1(n_232), .A2(n_262), .B1(n_1445), .B2(n_1448), .Y(n_1474) );
AO22x2_ASAP7_75t_L g1207 ( .A1(n_233), .A2(n_1208), .B1(n_1257), .B2(n_1258), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_233), .Y(n_1257) );
CKINVDCx5p33_ASAP7_75t_R g1266 ( .A(n_234), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_235), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g1201 ( .A(n_236), .Y(n_1201) );
INVx1_ASAP7_75t_L g1070 ( .A(n_239), .Y(n_1070) );
INVx1_ASAP7_75t_L g478 ( .A(n_240), .Y(n_478) );
INVx1_ASAP7_75t_L g522 ( .A(n_241), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_241), .A2(n_250), .B1(n_537), .B2(n_539), .Y(n_551) );
INVx1_ASAP7_75t_L g659 ( .A(n_244), .Y(n_659) );
INVx1_ASAP7_75t_L g449 ( .A(n_245), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_246), .A2(n_276), .B1(n_716), .B2(n_719), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_246), .A2(n_276), .B1(n_770), .B2(n_774), .C(n_777), .Y(n_769) );
INVx1_ASAP7_75t_L g1304 ( .A(n_248), .Y(n_1304) );
INVx1_ASAP7_75t_L g511 ( .A(n_250), .Y(n_511) );
INVx1_ASAP7_75t_L g949 ( .A(n_251), .Y(n_949) );
INVx1_ASAP7_75t_L g1119 ( .A(n_252), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g1280 ( .A1(n_253), .A2(n_1015), .B(n_1281), .C(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1317 ( .A(n_253), .Y(n_1317) );
INVx1_ASAP7_75t_L g1465 ( .A(n_254), .Y(n_1465) );
INVx1_ASAP7_75t_L g1699 ( .A(n_256), .Y(n_1699) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_257), .Y(n_814) );
INVx1_ASAP7_75t_L g1428 ( .A(n_258), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_258), .B(n_1437), .Y(n_1440) );
INVx1_ASAP7_75t_L g591 ( .A(n_259), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_260), .A2(n_612), .B1(n_613), .B2(n_624), .C(n_632), .Y(n_611) );
INVx1_ASAP7_75t_L g399 ( .A(n_261), .Y(n_399) );
INVx1_ASAP7_75t_L g746 ( .A(n_263), .Y(n_746) );
INVx1_ASAP7_75t_L g1243 ( .A(n_264), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_265), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g1165 ( .A(n_268), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g1271 ( .A1(n_269), .A2(n_946), .B(n_1118), .C(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1301 ( .A(n_269), .Y(n_1301) );
INVx1_ASAP7_75t_L g505 ( .A(n_270), .Y(n_505) );
INVx1_ASAP7_75t_L g943 ( .A(n_271), .Y(n_943) );
INVx1_ASAP7_75t_L g575 ( .A(n_272), .Y(n_575) );
INVx1_ASAP7_75t_L g1108 ( .A(n_273), .Y(n_1108) );
AOI21xp33_ASAP7_75t_L g1142 ( .A1(n_273), .A2(n_1143), .B(n_1144), .Y(n_1142) );
INVx2_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_275), .Y(n_739) );
INVx1_ASAP7_75t_L g1109 ( .A(n_277), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_278), .A2(n_279), .B1(n_678), .B2(n_1180), .Y(n_1181) );
OAI211xp5_ASAP7_75t_SL g1187 ( .A1(n_278), .A2(n_612), .B(n_1188), .C(n_1197), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1198 ( .A1(n_279), .A2(n_639), .B1(n_915), .B2(n_1199), .C(n_1202), .Y(n_1198) );
INVx1_ASAP7_75t_L g384 ( .A(n_280), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_280), .A2(n_294), .B1(n_440), .B2(n_442), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_281), .A2(n_286), .B1(n_566), .B2(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_281), .A2(n_286), .B1(n_609), .B2(n_610), .Y(n_839) );
INVx1_ASAP7_75t_L g925 ( .A(n_282), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g1133 ( .A(n_283), .Y(n_1133) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_285), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_287), .Y(n_636) );
BUFx3_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
INVx1_ASAP7_75t_L g432 ( .A(n_288), .Y(n_432) );
BUFx3_ASAP7_75t_L g340 ( .A(n_289), .Y(n_340) );
INVx1_ASAP7_75t_L g428 ( .A(n_289), .Y(n_428) );
INVx1_ASAP7_75t_L g884 ( .A(n_290), .Y(n_884) );
INVxp33_ASAP7_75t_SL g913 ( .A(n_293), .Y(n_913) );
INVx1_ASAP7_75t_L g402 ( .A(n_294), .Y(n_402) );
INVx1_ASAP7_75t_L g848 ( .A(n_295), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_296), .Y(n_1284) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_318), .B(n_1413), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
AND2x4_ASAP7_75t_L g1705 ( .A(n_300), .B(n_306), .Y(n_1705) );
NOR2xp33_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_SL g1710 ( .A(n_301), .Y(n_1710) );
NAND2xp5_ASAP7_75t_L g1721 ( .A(n_301), .B(n_303), .Y(n_1721) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_303), .B(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_311), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g597 ( .A(n_308), .B(n_329), .Y(n_597) );
OR2x6_ASAP7_75t_L g940 ( .A(n_308), .B(n_329), .Y(n_940) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g535 ( .A(n_309), .B(n_317), .Y(n_535) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g406 ( .A(n_310), .B(n_407), .Y(n_406) );
INVx8_ASAP7_75t_L g593 ( .A(n_311), .Y(n_593) );
OR2x6_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
OR2x6_ASAP7_75t_L g596 ( .A(n_312), .B(n_586), .Y(n_596) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_312), .Y(n_621) );
OR2x2_ASAP7_75t_L g749 ( .A(n_312), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g785 ( .A(n_312), .Y(n_785) );
INVx2_ASAP7_75t_SL g800 ( .A(n_312), .Y(n_800) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_312), .Y(n_1116) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_315), .Y(n_352) );
INVx2_ASAP7_75t_L g358 ( .A(n_314), .Y(n_358) );
AND2x4_ASAP7_75t_L g364 ( .A(n_314), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g373 ( .A(n_314), .Y(n_373) );
INVx1_ASAP7_75t_L g415 ( .A(n_314), .Y(n_415) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
INVx2_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
INVx1_ASAP7_75t_L g389 ( .A(n_315), .Y(n_389) );
INVx1_ASAP7_75t_L g414 ( .A(n_315), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_315), .B(n_358), .Y(n_628) );
AND2x4_ASAP7_75t_L g581 ( .A(n_316), .B(n_389), .Y(n_581) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g582 ( .A(n_317), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_317), .B(n_583), .Y(n_1076) );
XNOR2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_931), .Y(n_318) );
OA22x2_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_601), .B1(n_602), .B2(n_930), .Y(n_319) );
INVx1_ASAP7_75t_L g930 ( .A(n_320), .Y(n_930) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI21x1_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_491), .B(n_600), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g600 ( .A(n_323), .B(n_492), .Y(n_600) );
XOR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_490), .Y(n_323) );
NOR3xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_353), .C(n_418), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_327), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_327), .B(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_327), .B(n_880), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_327), .B(n_1185), .Y(n_1184) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_341), .Y(n_327) );
INVx2_ASAP7_75t_L g751 ( .A(n_328), .Y(n_751) );
AOI222xp33_ASAP7_75t_L g1407 ( .A1(n_328), .A2(n_450), .B1(n_464), .B2(n_1399), .C1(n_1402), .C2(n_1408), .Y(n_1407) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g446 ( .A(n_329), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g572 ( .A(n_329), .B(n_447), .Y(n_572) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_336), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_331), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g717 ( .A(n_331), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g720 ( .A(n_331), .B(n_474), .Y(n_720) );
INVx1_ASAP7_75t_L g737 ( .A(n_331), .Y(n_737) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_331), .B(n_718), .Y(n_1138) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g447 ( .A(n_334), .B(n_424), .Y(n_447) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g423 ( .A(n_335), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g499 ( .A(n_335), .Y(n_499) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_335), .Y(n_504) );
INVx1_ASAP7_75t_L g508 ( .A(n_335), .Y(n_508) );
BUFx2_ASAP7_75t_L g434 ( .A(n_336), .Y(n_434) );
INVx2_ASAP7_75t_L g441 ( .A(n_336), .Y(n_441) );
AND2x4_ASAP7_75t_L g502 ( .A(n_336), .B(n_503), .Y(n_502) );
INVx6_ASAP7_75t_L g525 ( .A(n_336), .Y(n_525) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g475 ( .A(n_337), .Y(n_475) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g427 ( .A(n_338), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g438 ( .A(n_338), .B(n_340), .Y(n_438) );
INVx1_ASAP7_75t_L g483 ( .A(n_339), .Y(n_483) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g431 ( .A(n_340), .B(n_432), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx2_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g421 ( .A(n_343), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g534 ( .A(n_343), .B(n_535), .Y(n_534) );
OR2x6_ASAP7_75t_L g556 ( .A(n_343), .B(n_557), .Y(n_556) );
OAI31xp33_ASAP7_75t_L g607 ( .A1(n_343), .A2(n_608), .A3(n_611), .B(n_638), .Y(n_607) );
BUFx2_ASAP7_75t_L g867 ( .A(n_343), .Y(n_867) );
AND2x4_ASAP7_75t_L g963 ( .A(n_343), .B(n_535), .Y(n_963) );
OR2x2_ASAP7_75t_L g978 ( .A(n_343), .B(n_557), .Y(n_978) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g530 ( .A(n_344), .Y(n_530) );
OR2x6_ASAP7_75t_L g782 ( .A(n_344), .B(n_406), .Y(n_782) );
INVx1_ASAP7_75t_L g1212 ( .A(n_345), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
AND2x2_ASAP7_75t_L g634 ( .A(n_346), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_347), .B(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g411 ( .A(n_347), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g915 ( .A(n_347), .B(n_412), .Y(n_915) );
INVx1_ASAP7_75t_L g1405 ( .A(n_347), .Y(n_1405) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g861 ( .A(n_350), .Y(n_861) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g538 ( .A(n_351), .Y(n_538) );
INVx2_ASAP7_75t_SL g766 ( .A(n_351), .Y(n_766) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_352), .Y(n_368) );
AOI31xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_393), .A3(n_400), .B(n_416), .Y(n_353) );
AOI221xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_366), .B1(n_380), .B2(n_384), .C(n_385), .Y(n_354) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_383), .Y(n_394) );
BUFx2_ASAP7_75t_L g542 ( .A(n_357), .Y(n_542) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_357), .Y(n_549) );
AND2x4_ASAP7_75t_L g585 ( .A(n_357), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g967 ( .A(n_357), .Y(n_967) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_357), .Y(n_1038) );
BUFx6f_ASAP7_75t_L g1393 ( .A(n_357), .Y(n_1393) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g847 ( .A(n_362), .Y(n_847) );
INVx2_ASAP7_75t_L g969 ( .A(n_362), .Y(n_969) );
INVx2_ASAP7_75t_L g972 ( .A(n_362), .Y(n_972) );
INVx2_ASAP7_75t_L g1355 ( .A(n_362), .Y(n_1355) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_363), .Y(n_647) );
INVx3_ASAP7_75t_L g758 ( .A(n_363), .Y(n_758) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g398 ( .A(n_364), .Y(n_398) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_364), .Y(n_545) );
INVx1_ASAP7_75t_L g590 ( .A(n_364), .Y(n_590) );
AND2x4_ASAP7_75t_L g372 ( .A(n_365), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g401 ( .A(n_368), .B(n_383), .Y(n_401) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
INVx3_ASAP7_75t_L g1196 ( .A(n_368), .Y(n_1196) );
AOI211xp5_ASAP7_75t_L g574 ( .A1(n_369), .A2(n_575), .B(n_576), .C(n_579), .Y(n_574) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g1194 ( .A(n_370), .Y(n_1194) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g380 ( .A(n_371), .B(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_372), .Y(n_405) );
AND2x4_ASAP7_75t_L g576 ( .A(n_372), .B(n_577), .Y(n_576) );
BUFx3_ASAP7_75t_L g762 ( .A(n_372), .Y(n_762) );
BUFx6f_ASAP7_75t_L g975 ( .A(n_372), .Y(n_975) );
INVx1_ASAP7_75t_L g623 ( .A(n_374), .Y(n_623) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x6_ASAP7_75t_L g553 ( .A(n_376), .B(n_477), .Y(n_553) );
BUFx2_ASAP7_75t_L g863 ( .A(n_376), .Y(n_863) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g578 ( .A(n_377), .Y(n_578) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
INVx8_ASAP7_75t_L g612 ( .A(n_380), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g1210 ( .A1(n_380), .A2(n_401), .B1(n_1211), .B2(n_1212), .C1(n_1213), .C2(n_1214), .Y(n_1210) );
AND2x4_ASAP7_75t_L g396 ( .A(n_381), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g759 ( .A(n_383), .B(n_454), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
NAND2x1_ASAP7_75t_SL g772 ( .A(n_387), .B(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g1404 ( .A1(n_387), .A2(n_959), .B1(n_1384), .B2(n_1385), .Y(n_1404) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_389), .Y(n_635) );
CKINVDCx11_ASAP7_75t_R g637 ( .A(n_391), .Y(n_637) );
INVx1_ASAP7_75t_L g776 ( .A(n_392), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_396), .B2(n_399), .Y(n_393) );
INVx3_ASAP7_75t_L g609 ( .A(n_394), .Y(n_609) );
INVx3_ASAP7_75t_L g906 ( .A(n_394), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_394), .A2(n_396), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_394), .A2(n_396), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
INVx3_ASAP7_75t_L g610 ( .A(n_396), .Y(n_610) );
INVx3_ASAP7_75t_L g907 ( .A(n_396), .Y(n_907) );
INVx1_ASAP7_75t_L g921 ( .A(n_397), .Y(n_921) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g409 ( .A(n_398), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_403), .B2(n_408), .C(n_410), .Y(n_400) );
CKINVDCx6p67_ASAP7_75t_R g639 ( .A(n_401), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g1391 ( .A1(n_401), .A2(n_1392), .B1(n_1394), .B2(n_1395), .Y(n_1391) );
INVx1_ASAP7_75t_L g1089 ( .A(n_404), .Y(n_1089) );
INVx2_ASAP7_75t_SL g540 ( .A(n_405), .Y(n_540) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_405), .Y(n_862) );
INVx1_ASAP7_75t_L g586 ( .A(n_407), .Y(n_586) );
INVx1_ASAP7_75t_L g858 ( .A(n_409), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g1218 ( .A(n_410), .B(n_1219), .C(n_1233), .Y(n_1218) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g651 ( .A(n_412), .Y(n_651) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g850 ( .A(n_413), .Y(n_850) );
BUFx2_ASAP7_75t_L g911 ( .A(n_413), .Y(n_911) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_414), .B(n_415), .Y(n_617) );
INVx1_ASAP7_75t_L g583 ( .A(n_415), .Y(n_583) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI31xp33_ASAP7_75t_L g904 ( .A1(n_417), .A2(n_905), .A3(n_908), .B(n_916), .Y(n_904) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_419), .B(n_448), .C(n_462), .D(n_470), .Y(n_418) );
AOI33xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_425), .A3(n_433), .B1(n_439), .B2(n_444), .B3(n_446), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g1361 ( .A(n_420), .B(n_1362), .C(n_1364), .Y(n_1361) );
NAND3xp33_ASAP7_75t_L g1680 ( .A(n_420), .B(n_1681), .C(n_1682), .Y(n_1680) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g557 ( .A(n_423), .Y(n_557) );
INVx2_ASAP7_75t_SL g729 ( .A(n_423), .Y(n_729) );
BUFx3_ASAP7_75t_L g1150 ( .A(n_423), .Y(n_1150) );
INVx1_ASAP7_75t_L g529 ( .A(n_424), .Y(n_529) );
BUFx3_ASAP7_75t_L g565 ( .A(n_426), .Y(n_565) );
INVx2_ASAP7_75t_SL g709 ( .A(n_426), .Y(n_709) );
AND2x4_ASAP7_75t_L g712 ( .A(n_426), .B(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_SL g469 ( .A(n_427), .Y(n_469) );
AND2x6_ASAP7_75t_L g527 ( .A(n_427), .B(n_498), .Y(n_527) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_427), .Y(n_571) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_427), .Y(n_683) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_427), .Y(n_724) );
BUFx3_ASAP7_75t_L g897 ( .A(n_427), .Y(n_897) );
BUFx2_ASAP7_75t_L g980 ( .A(n_427), .Y(n_980) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_427), .Y(n_1177) );
INVx1_ASAP7_75t_L g461 ( .A(n_428), .Y(n_461) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x6_ASAP7_75t_L g451 ( .A(n_430), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g870 ( .A(n_430), .B(n_452), .Y(n_870) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_431), .Y(n_445) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_431), .Y(n_509) );
INVx2_ASAP7_75t_L g671 ( .A(n_431), .Y(n_671) );
INVx1_ASAP7_75t_L g888 ( .A(n_431), .Y(n_888) );
INVx1_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g1363 ( .A(n_436), .Y(n_1363) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
AND2x4_ASAP7_75t_L g496 ( .A(n_437), .B(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_437), .Y(n_513) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_437), .Y(n_563) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_438), .Y(n_443) );
AND2x2_ASAP7_75t_L g464 ( .A(n_440), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g568 ( .A(n_441), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_442), .B(n_489), .Y(n_689) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_442), .Y(n_1254) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g676 ( .A(n_443), .Y(n_676) );
AND2x4_ASAP7_75t_L g733 ( .A(n_443), .B(n_713), .Y(n_733) );
INVx1_ASAP7_75t_L g984 ( .A(n_443), .Y(n_984) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_443), .Y(n_1045) );
BUFx4f_ASAP7_75t_L g1066 ( .A(n_443), .Y(n_1066) );
INVx1_ASAP7_75t_L g1246 ( .A(n_443), .Y(n_1246) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_445), .Y(n_566) );
BUFx3_ASAP7_75t_L g731 ( .A(n_445), .Y(n_731) );
INVx1_ASAP7_75t_L g821 ( .A(n_445), .Y(n_821) );
INVx1_ASAP7_75t_L g686 ( .A(n_446), .Y(n_686) );
AOI33xp33_ASAP7_75t_L g976 ( .A1(n_446), .A2(n_977), .A3(n_979), .B1(n_981), .B2(n_982), .B3(n_985), .Y(n_976) );
AOI33xp33_ASAP7_75t_L g1174 ( .A1(n_446), .A2(n_1175), .A3(n_1176), .B1(n_1179), .B2(n_1181), .B3(n_1182), .Y(n_1174) );
AOI33xp33_ASAP7_75t_L g1375 ( .A1(n_446), .A2(n_977), .A3(n_1376), .B1(n_1378), .B2(n_1379), .B3(n_1382), .Y(n_1375) );
NAND3xp33_ASAP7_75t_L g1689 ( .A(n_446), .B(n_1690), .C(n_1692), .Y(n_1689) );
INVx2_ASAP7_75t_L g706 ( .A(n_447), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_447), .Y(n_1144) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_455), .B2(n_456), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_450), .A2(n_456), .B1(n_618), .B2(n_631), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_450), .A2(n_456), .B1(n_1165), .B2(n_1166), .Y(n_1164) );
CKINVDCx6p67_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g457 ( .A(n_452), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
OR2x2_ASAP7_75t_L g872 ( .A(n_452), .B(n_873), .Y(n_872) );
OR2x2_ASAP7_75t_L g874 ( .A(n_452), .B(n_875), .Y(n_874) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g713 ( .A(n_453), .Y(n_713) );
OR2x2_ASAP7_75t_L g741 ( .A(n_453), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g745 ( .A(n_453), .B(n_671), .Y(n_745) );
INVx1_ASAP7_75t_L g477 ( .A(n_454), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g1409 ( .A1(n_456), .A2(n_467), .B1(n_1400), .B2(n_1410), .Y(n_1409) );
CKINVDCx6p67_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g1300 ( .A(n_458), .Y(n_1300) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx4f_ASAP7_75t_L g818 ( .A(n_459), .Y(n_818) );
INVx1_ASAP7_75t_L g829 ( .A(n_459), .Y(n_829) );
INVx1_ASAP7_75t_L g1332 ( .A(n_459), .Y(n_1332) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OR2x2_ASAP7_75t_L g742 ( .A(n_460), .B(n_461), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_466), .B2(n_467), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_464), .A2(n_467), .B1(n_622), .B2(n_629), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_464), .A2(n_467), .B1(n_1168), .B2(n_1169), .Y(n_1167) );
AND2x2_ASAP7_75t_L g467 ( .A(n_465), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_469), .A2(n_1303), .B1(n_1304), .B2(n_1305), .Y(n_1302) );
INVx1_ASAP7_75t_L g1377 ( .A(n_469), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_478), .B1(n_479), .B2(n_485), .C(n_486), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_471), .A2(n_633), .B1(n_636), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_471), .A2(n_902), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_471), .A2(n_479), .B1(n_486), .B2(n_1384), .C(n_1385), .Y(n_1383) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
OR2x2_ASAP7_75t_L g903 ( .A(n_473), .B(n_476), .Y(n_903) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g520 ( .A(n_475), .B(n_499), .Y(n_520) );
INVx2_ASAP7_75t_SL g484 ( .A(n_476), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_476), .Y(n_489) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g663 ( .A(n_480), .Y(n_663) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_480), .Y(n_835) );
INVx1_ASAP7_75t_L g902 ( .A(n_480), .Y(n_902) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g718 ( .A(n_482), .Y(n_718) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g518 ( .A(n_483), .Y(n_518) );
BUFx2_ASAP7_75t_L g808 ( .A(n_486), .Y(n_808) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g703 ( .A(n_488), .Y(n_703) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
AOI211x1_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_528), .B(n_531), .C(n_573), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .C(n_510), .D(n_521), .Y(n_494) );
NAND4xp25_ASAP7_75t_SL g1057 ( .A(n_495), .B(n_1058), .C(n_1061), .D(n_1064), .Y(n_1057) );
BUFx2_ASAP7_75t_L g1247 ( .A(n_495), .Y(n_1247) );
INVx5_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI211xp5_ASAP7_75t_L g988 ( .A1(n_496), .A2(n_989), .B(n_990), .C(n_991), .Y(n_988) );
CKINVDCx8_ASAP7_75t_R g1015 ( .A(n_496), .Y(n_1015) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_496), .B(n_1329), .Y(n_1328) );
AOI211xp5_ASAP7_75t_L g1669 ( .A1(n_496), .A2(n_1670), .B(n_1671), .C(n_1672), .Y(n_1669) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g990 ( .A(n_498), .B(n_513), .Y(n_990) );
INVx1_ASAP7_75t_L g1021 ( .A(n_498), .Y(n_1021) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_505), .B2(n_506), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_501), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_502), .A2(n_949), .B1(n_997), .B2(n_998), .Y(n_996) );
INVx4_ASAP7_75t_L g1022 ( .A(n_502), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_502), .A2(n_506), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_502), .A2(n_506), .B1(n_1211), .B2(n_1243), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_502), .A2(n_523), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1673 ( .A1(n_502), .A2(n_523), .B1(n_1674), .B2(n_1675), .Y(n_1673) );
AND2x4_ASAP7_75t_L g516 ( .A(n_503), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_SL g1285 ( .A(n_503), .B(n_517), .Y(n_1285) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_506), .A2(n_527), .B1(n_1000), .B2(n_1001), .Y(n_999) );
INVx4_ASAP7_75t_L g1018 ( .A(n_506), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_506), .A2(n_527), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1676 ( .A1(n_506), .A2(n_527), .B1(n_1677), .B2(n_1678), .Y(n_1676) );
AND2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g523 ( .A(n_507), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g998 ( .A(n_507), .B(n_524), .Y(n_998) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g993 ( .A(n_508), .B(n_994), .Y(n_993) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_509), .Y(n_684) );
INVx2_ASAP7_75t_L g899 ( .A(n_509), .Y(n_899) );
BUFx6f_ASAP7_75t_L g986 ( .A(n_509), .Y(n_986) );
INVx1_ASAP7_75t_L g1305 ( .A(n_509), .Y(n_1305) );
AOI222xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_514), .B2(n_515), .C1(n_519), .C2(n_520), .Y(n_510) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g1671 ( .A(n_513), .Y(n_1671) );
AOI222xp33_ASAP7_75t_L g1244 ( .A1(n_515), .A2(n_520), .B1(n_1231), .B2(n_1232), .C1(n_1236), .C2(n_1245), .Y(n_1244) );
BUFx4f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_516), .A2(n_520), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
INVx1_ASAP7_75t_L g1069 ( .A(n_516), .Y(n_1069) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g994 ( .A(n_518), .Y(n_994) );
INVx3_ASAP7_75t_L g995 ( .A(n_520), .Y(n_995) );
AOI222xp33_ASAP7_75t_L g1064 ( .A1(n_520), .A2(n_1065), .B1(n_1066), .B2(n_1067), .C1(n_1068), .C2(n_1070), .Y(n_1064) );
AOI322xp5_ASAP7_75t_L g1282 ( .A1(n_520), .A2(n_683), .A3(n_1275), .B1(n_1276), .B2(n_1283), .C1(n_1284), .C2(n_1285), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_526), .B2(n_527), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_523), .A2(n_527), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_523), .A2(n_527), .B1(n_1240), .B2(n_1241), .Y(n_1239) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g560 ( .A(n_525), .Y(n_560) );
INVx2_ASAP7_75t_L g674 ( .A(n_525), .Y(n_674) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_525), .Y(n_679) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_525), .Y(n_1143) );
INVx1_ASAP7_75t_L g1367 ( .A(n_525), .Y(n_1367) );
CKINVDCx6p67_ASAP7_75t_R g1017 ( .A(n_527), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_528), .Y(n_1071) );
AO211x2_ASAP7_75t_L g1667 ( .A1(n_528), .A2(n_1668), .B(n_1679), .C(n_1693), .Y(n_1667) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_529), .B(n_530), .Y(n_1003) );
INVx2_ASAP7_75t_L g699 ( .A(n_530), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_554), .Y(n_531) );
AOI33xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .A3(n_541), .B1(n_546), .B2(n_551), .B3(n_552), .Y(n_532) );
AOI33xp33_ASAP7_75t_L g1083 ( .A1(n_533), .A2(n_552), .A3(n_1084), .B1(n_1085), .B2(n_1086), .B3(n_1087), .Y(n_1083) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g1686 ( .A(n_534), .B(n_1687), .C(n_1688), .Y(n_1686) );
INVx1_ASAP7_75t_L g657 ( .A(n_535), .Y(n_657) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI211xp5_ASAP7_75t_L g1694 ( .A1(n_539), .A2(n_576), .B(n_1695), .C(n_1696), .Y(n_1694) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g953 ( .A(n_540), .Y(n_953) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_544), .A2(n_714), .B1(n_743), .B2(n_790), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_544), .A2(n_626), .B1(n_913), .B2(n_914), .Y(n_912) );
INVx2_ASAP7_75t_L g1234 ( .A(n_544), .Y(n_1234) );
INVx4_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g550 ( .A(n_545), .Y(n_550) );
INVx2_ASAP7_75t_SL g630 ( .A(n_545), .Y(n_630) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g768 ( .A(n_549), .B(n_759), .Y(n_768) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_549), .B(n_759), .Y(n_1110) );
INVx1_ASAP7_75t_L g1127 ( .A(n_550), .Y(n_1127) );
AOI33xp33_ASAP7_75t_L g962 ( .A1(n_552), .A2(n_963), .A3(n_964), .B1(n_965), .B2(n_970), .B3(n_973), .Y(n_962) );
AOI33xp33_ASAP7_75t_L g1031 ( .A1(n_552), .A2(n_963), .A3(n_1032), .B1(n_1035), .B2(n_1037), .B3(n_1039), .Y(n_1031) );
INVx2_ASAP7_75t_L g1318 ( .A(n_552), .Y(n_1318) );
INVx6_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx5_ASAP7_75t_L g803 ( .A(n_553), .Y(n_803) );
AOI33xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .A3(n_564), .B1(n_567), .B2(n_569), .B3(n_572), .Y(n_554) );
AOI33xp33_ASAP7_75t_L g1040 ( .A1(n_555), .A2(n_572), .A3(n_1041), .B1(n_1044), .B2(n_1046), .B3(n_1049), .Y(n_1040) );
AOI33xp33_ASAP7_75t_L g1090 ( .A1(n_555), .A2(n_1091), .A3(n_1094), .B1(n_1095), .B2(n_1096), .B3(n_1097), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_556), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g809 ( .A1(n_556), .A2(n_810), .B1(n_822), .B2(n_823), .Y(n_809) );
OAI22xp5_ASAP7_75t_SL g882 ( .A1(n_556), .A2(n_883), .B1(n_889), .B2(n_891), .Y(n_882) );
INVx2_ASAP7_75t_L g1175 ( .A(n_556), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_556), .A2(n_889), .B1(n_1249), .B2(n_1255), .Y(n_1248) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_560), .Y(n_1047) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g726 ( .A(n_563), .Y(n_726) );
AND2x4_ASAP7_75t_L g735 ( .A(n_563), .B(n_736), .Y(n_735) );
BUFx6f_ASAP7_75t_L g1048 ( .A(n_563), .Y(n_1048) );
INVx1_ASAP7_75t_L g1148 ( .A(n_563), .Y(n_1148) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx4f_ASAP7_75t_L g667 ( .A(n_571), .Y(n_667) );
INVx1_ASAP7_75t_L g875 ( .A(n_571), .Y(n_875) );
INVx4_ASAP7_75t_L g822 ( .A(n_572), .Y(n_822) );
BUFx4f_ASAP7_75t_L g890 ( .A(n_572), .Y(n_890) );
BUFx4f_ASAP7_75t_L g1097 ( .A(n_572), .Y(n_1097) );
AOI31xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_584), .A3(n_592), .B(n_597), .Y(n_573) );
CKINVDCx11_ASAP7_75t_R g946 ( .A(n_576), .Y(n_946) );
NOR3xp33_ASAP7_75t_L g1024 ( .A(n_576), .B(n_1025), .C(n_1027), .Y(n_1024) );
AOI211xp5_ASAP7_75t_L g1073 ( .A1(n_576), .A2(n_1033), .B(n_1074), .C(n_1075), .Y(n_1073) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVxp67_ASAP7_75t_L g960 ( .A(n_578), .Y(n_960) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g956 ( .A(n_581), .Y(n_956) );
INVx2_ASAP7_75t_L g1026 ( .A(n_581), .Y(n_1026) );
AOI322xp5_ASAP7_75t_L g1272 ( .A1(n_581), .A2(n_958), .A3(n_1269), .B1(n_1273), .B2(n_1274), .C1(n_1275), .C2(n_1276), .Y(n_1272) );
INVx1_ASAP7_75t_L g959 ( .A(n_583), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_588), .B2(n_591), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_585), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_585), .A2(n_588), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_585), .A2(n_945), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_585), .A2(n_945), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
AOI22xp33_ASAP7_75t_SL g1697 ( .A1(n_585), .A2(n_588), .B1(n_1698), .B2(n_1699), .Y(n_1697) );
AND2x4_ASAP7_75t_L g588 ( .A(n_586), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g945 ( .A(n_586), .B(n_589), .Y(n_945) );
INVx1_ASAP7_75t_L g1269 ( .A(n_586), .Y(n_1269) );
INVx5_ASAP7_75t_SL g1270 ( .A(n_588), .Y(n_1270) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_590), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_593), .A2(n_948), .B1(n_949), .B2(n_950), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_593), .A2(n_950), .B1(n_1062), .B2(n_1081), .Y(n_1080) );
AOI211xp5_ASAP7_75t_L g1265 ( .A1(n_593), .A2(n_1266), .B(n_1267), .C(n_1271), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_593), .A2(n_595), .B1(n_1335), .B2(n_1348), .Y(n_1347) );
AOI22xp33_ASAP7_75t_SL g1700 ( .A1(n_593), .A2(n_595), .B1(n_1675), .B2(n_1701), .Y(n_1700) );
INVx5_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx4_ASAP7_75t_L g950 ( .A(n_596), .Y(n_950) );
OAI211xp5_ASAP7_75t_L g1264 ( .A1(n_597), .A2(n_1265), .B(n_1277), .C(n_1286), .Y(n_1264) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
XNOR2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_804), .Y(n_602) );
AOI22x1_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_693), .B2(n_694), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_658), .C(n_660), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_618), .B1(n_619), .B2(n_622), .C(n_623), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g787 ( .A(n_615), .Y(n_787) );
INVx2_ASAP7_75t_L g1316 ( .A(n_615), .Y(n_1316) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx3_ASAP7_75t_L g801 ( .A(n_616), .Y(n_801) );
BUFx3_ASAP7_75t_L g1222 ( .A(n_616), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_616), .B(n_1404), .Y(n_1403) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_619), .A2(n_656), .B1(n_884), .B2(n_885), .C(n_910), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g1199 ( .A1(n_619), .A2(n_656), .B1(n_1118), .B2(n_1200), .C(n_1201), .Y(n_1199) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g654 ( .A(n_621), .Y(n_654) );
BUFx2_ASAP7_75t_L g851 ( .A(n_621), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g1307 ( .A1(n_621), .A2(n_650), .B1(n_1295), .B2(n_1297), .Y(n_1307) );
OAI22xp33_ASAP7_75t_L g1314 ( .A1(n_621), .A2(n_1315), .B1(n_1316), .B2(n_1317), .Y(n_1314) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_626), .A2(n_1203), .B1(n_1204), .B2(n_1205), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_626), .A2(n_969), .B1(n_1399), .B2(n_1400), .Y(n_1398) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g1190 ( .A(n_627), .Y(n_1190) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g643 ( .A(n_628), .Y(n_643) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_628), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_630), .A2(n_790), .B1(n_794), .B2(n_795), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_634), .A2(n_637), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_634), .A2(n_637), .B1(n_925), .B2(n_926), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_634), .A2(n_637), .B1(n_1172), .B2(n_1173), .Y(n_1197) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_634), .A2(n_637), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B1(n_645), .B2(n_648), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g843 ( .A(n_642), .Y(n_843) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx3_ASAP7_75t_L g793 ( .A(n_643), .Y(n_793) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_SL g1124 ( .A(n_647), .Y(n_1124) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_653), .B2(n_655), .C(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_656), .A2(n_814), .B1(n_815), .B2(n_850), .C(n_851), .Y(n_849) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g660 ( .A(n_661), .B(n_690), .Y(n_660) );
NAND3xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_664), .C(n_687), .Y(n_661) );
AOI33xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .A3(n_672), .B1(n_677), .B2(n_680), .B3(n_685), .Y(n_664) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g1178 ( .A(n_669), .Y(n_1178) );
INVx1_ASAP7_75t_L g1183 ( .A(n_669), .Y(n_1183) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g711 ( .A(n_670), .Y(n_711) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g1293 ( .A(n_671), .Y(n_1293) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g1011 ( .A(n_676), .Y(n_1011) );
INVx1_ASAP7_75t_L g1180 ( .A(n_676), .Y(n_1180) );
INVx4_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g704 ( .A(n_679), .Y(n_704) );
INVx2_ASAP7_75t_L g1691 ( .A(n_679), .Y(n_1691) );
INVx1_ASAP7_75t_L g1290 ( .A(n_681), .Y(n_1290) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g1253 ( .A(n_682), .Y(n_1253) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g1365 ( .A(n_685), .B(n_1366), .C(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_687), .B(n_1171), .C(n_1174), .Y(n_1170) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
XNOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_752), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_746), .B2(n_747), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx8_ASAP7_75t_SL g1406 ( .A(n_699), .Y(n_1406) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_721), .C(n_738), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_707), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_701) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g1042 ( .A(n_709), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_712), .A2(n_1126), .B(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_730), .B1(n_732), .B2(n_734), .C(n_735), .Y(n_721) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g833 ( .A(n_724), .Y(n_833) );
BUFx3_ASAP7_75t_L g1092 ( .A(n_724), .Y(n_1092) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_732), .A2(n_735), .B1(n_1131), .B2(n_1146), .C(n_1151), .Y(n_1145) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_734), .A2(n_739), .B1(n_798), .B2(n_801), .Y(n_797) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_740), .A2(n_744), .B1(n_1128), .B2(n_1130), .Y(n_1152) );
INVx6_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g813 ( .A(n_742), .Y(n_813) );
INVx2_ASAP7_75t_L g825 ( .A(n_742), .Y(n_825) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_742), .B(n_1021), .Y(n_1020) );
INVx4_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g1132 ( .A1(n_747), .A2(n_1133), .B(n_1134), .Y(n_1132) );
INVx5_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx3_ASAP7_75t_L g773 ( .A(n_750), .Y(n_773) );
NOR3xp33_ASAP7_75t_SL g752 ( .A(n_753), .B(n_769), .C(n_779), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_763), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_760), .B2(n_761), .Y(n_754) );
BUFx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_757), .Y(n_1105) );
AND2x4_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g1228 ( .A(n_758), .Y(n_1228) );
INVx2_ASAP7_75t_L g1359 ( .A(n_758), .Y(n_1359) );
AND2x6_ASAP7_75t_L g761 ( .A(n_759), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g765 ( .A(n_759), .B(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_761), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
NAND2x1p5_ASAP7_75t_L g778 ( .A(n_762), .B(n_773), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_765), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1107) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_773), .B(n_776), .Y(n_775) );
BUFx4f_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_778), .Y(n_1112) );
OAI33xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .A3(n_789), .B1(n_796), .B2(n_797), .B3(n_802), .Y(n_779) );
OAI33xp33_ASAP7_75t_L g1113 ( .A1(n_780), .A2(n_802), .A3(n_1114), .B1(n_1120), .B2(n_1125), .B3(n_1129), .Y(n_1113) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI33xp33_ASAP7_75t_L g1306 ( .A1(n_782), .A2(n_1307), .A3(n_1308), .B1(n_1311), .B2(n_1314), .B3(n_1318), .Y(n_1306) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_SL g1312 ( .A(n_793), .Y(n_1312) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
CKINVDCx8_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g1350 ( .A(n_803), .B(n_1351), .C(n_1353), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1683 ( .A(n_803), .B(n_1684), .C(n_1685), .Y(n_1683) );
XOR2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_876), .Y(n_804) );
AND4x1_ASAP7_75t_L g806 ( .A(n_807), .B(n_836), .C(n_838), .D(n_868), .Y(n_806) );
NOR3xp33_ASAP7_75t_SL g807 ( .A(n_808), .B(n_809), .C(n_834), .Y(n_807) );
NOR3xp33_ASAP7_75t_SL g881 ( .A(n_808), .B(n_882), .C(n_900), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_814), .B1(n_815), .B2(n_816), .C(n_819), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_811), .A2(n_816), .B1(n_884), .B2(n_885), .C(n_886), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_811), .A2(n_1229), .B1(n_1250), .B2(n_1251), .C(n_1252), .Y(n_1249) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_812), .A2(n_827), .B1(n_1213), .B2(n_1214), .C(n_1256), .Y(n_1255) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g893 ( .A(n_818), .Y(n_893) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_818), .Y(n_1140) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OAI33xp33_ASAP7_75t_L g1287 ( .A1(n_822), .A2(n_978), .A3(n_1288), .B1(n_1294), .B2(n_1299), .B3(n_1302), .Y(n_1287) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_826), .B1(n_827), .B2(n_830), .C(n_831), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_824), .A2(n_892), .B1(n_893), .B2(n_894), .C(n_895), .Y(n_891) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g873 ( .A(n_825), .Y(n_873) );
INVx2_ASAP7_75t_L g1296 ( .A(n_825), .Y(n_1296) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
BUFx2_ASAP7_75t_L g1298 ( .A(n_829), .Y(n_1298) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
OAI31xp33_ASAP7_75t_SL g838 ( .A1(n_839), .A2(n_840), .A3(n_852), .B(n_867), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B1(n_845), .B2(n_848), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_842), .A2(n_1121), .B1(n_1122), .B2(n_1123), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_842), .A2(n_1126), .B1(n_1127), .B2(n_1128), .Y(n_1125) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g854 ( .A(n_843), .Y(n_854) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI21xp5_ASAP7_75t_SL g1235 ( .A1(n_850), .A2(n_1236), .B(n_1237), .Y(n_1235) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_851), .A2(n_1118), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_856), .B2(n_859), .C(n_860), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_854), .A2(n_918), .B1(n_919), .B2(n_922), .C(n_923), .Y(n_917) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
CKINVDCx8_ASAP7_75t_R g1154 ( .A(n_867), .Y(n_1154) );
AOI221x1_ASAP7_75t_SL g1208 ( .A1(n_867), .A2(n_1071), .B1(n_1209), .B2(n_1238), .C(n_1248), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .Y(n_868) );
XNOR2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
AND4x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .C(n_904), .D(n_927), .Y(n_878) );
INVx1_ASAP7_75t_L g1251 ( .A(n_887), .Y(n_1251) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g1043 ( .A(n_888), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
BUFx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1093 ( .A(n_899), .Y(n_1093) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g1118 ( .A(n_911), .Y(n_1118) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g1192 ( .A(n_921), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_921), .A2(n_1289), .B1(n_1291), .B2(n_1309), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
XNOR2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_1156), .Y(n_931) );
OA22x2_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_1053), .B1(n_1054), .B2(n_1155), .Y(n_932) );
INVx1_ASAP7_75t_L g1155 ( .A(n_933), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B1(n_1004), .B2(n_1052), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
XNOR2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g1421 ( .A1(n_937), .A2(n_1422), .B1(n_1429), .B2(n_1431), .Y(n_1421) );
AOI211xp5_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_941), .B(n_961), .C(n_987), .Y(n_938) );
AOI221x1_ASAP7_75t_L g1326 ( .A1(n_939), .A2(n_1071), .B1(n_1327), .B2(n_1339), .C(n_1349), .Y(n_1326) );
CKINVDCx16_ASAP7_75t_R g939 ( .A(n_940), .Y(n_939) );
AO21x1_ASAP7_75t_SL g1023 ( .A1(n_940), .A2(n_1024), .B(n_1028), .Y(n_1023) );
AOI31xp33_ASAP7_75t_L g1072 ( .A1(n_940), .A2(n_1073), .A3(n_1077), .B(n_1080), .Y(n_1072) );
AOI31xp33_ASAP7_75t_L g1693 ( .A1(n_940), .A2(n_1694), .A3(n_1697), .B(n_1700), .Y(n_1693) );
NAND4xp25_ASAP7_75t_SL g941 ( .A(n_942), .B(n_946), .C(n_947), .D(n_951), .Y(n_941) );
NAND4xp25_ASAP7_75t_SL g1339 ( .A(n_946), .B(n_1340), .C(n_1343), .D(n_1347), .Y(n_1339) );
AOI222xp33_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B1(n_954), .B2(n_955), .C1(n_957), .C2(n_958), .Y(n_951) );
AOI222xp33_ASAP7_75t_L g1343 ( .A1(n_953), .A2(n_955), .B1(n_958), .B2(n_1344), .C1(n_1345), .C2(n_1346), .Y(n_1343) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
AND2x4_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
NAND2xp5_ASAP7_75t_SL g961 ( .A(n_962), .B(n_976), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g1356 ( .A(n_963), .B(n_1357), .C(n_1360), .Y(n_1356) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g1036 ( .A(n_969), .Y(n_1036) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
BUFx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_975), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1352 ( .A(n_975), .Y(n_1352) );
INVx1_ASAP7_75t_SL g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AOI31xp33_ASAP7_75t_SL g987 ( .A1(n_988), .A2(n_996), .A3(n_999), .B(n_1002), .Y(n_987) );
INVx1_ASAP7_75t_L g1281 ( .A(n_990), .Y(n_1281) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_1003), .Y(n_1002) );
OAI31xp33_ASAP7_75t_L g1007 ( .A1(n_1003), .A2(n_1008), .A3(n_1016), .B(n_1019), .Y(n_1007) );
OAI31xp33_ASAP7_75t_SL g1277 ( .A1(n_1003), .A2(n_1278), .A3(n_1279), .B(n_1280), .Y(n_1277) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1004), .Y(n_1052) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
AND4x1_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1023), .C(n_1031), .D(n_1040), .Y(n_1006) );
NAND4xp25_ASAP7_75t_L g1051 ( .A(n_1007), .B(n_1023), .C(n_1031), .D(n_1040), .Y(n_1051) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .C(n_1015), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1021), .Y(n_1283) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
XNOR2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1098), .Y(n_1054) );
AOI211x1_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1071), .B(n_1072), .C(n_1082), .Y(n_1056) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1090), .Y(n_1082) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
XNOR2x1_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1100), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1132), .Y(n_1100) );
NOR3xp33_ASAP7_75t_SL g1101 ( .A(n_1102), .B(n_1111), .C(n_1113), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .Y(n_1102) );
OAI211xp5_ASAP7_75t_L g1139 ( .A1(n_1106), .A2(n_1140), .B(n_1141), .C(n_1142), .Y(n_1139) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_1115), .A2(n_1117), .B1(n_1118), .B2(n_1119), .Y(n_1114) );
INVx3_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1123), .A2(n_1284), .B1(n_1312), .B2(n_1313), .Y(n_1311) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI31xp33_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1145), .A3(n_1152), .B(n_1153), .Y(n_1134) );
INVx1_ASAP7_75t_SL g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1143), .Y(n_1381) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
OAI31xp33_ASAP7_75t_L g1186 ( .A1(n_1153), .A2(n_1187), .A3(n_1198), .B(n_1206), .Y(n_1186) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
XOR2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1261), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1207), .B1(n_1259), .B2(n_1260), .Y(n_1158) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1159), .Y(n_1259) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1184), .C(n_1186), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1170), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1167), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1188 ( .A1(n_1165), .A2(n_1169), .B1(n_1189), .B2(n_1191), .C(n_1193), .Y(n_1188) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
A2O1A1Ixp33_ASAP7_75t_L g1401 ( .A1(n_1195), .A2(n_1402), .B(n_1403), .C(n_1405), .Y(n_1401) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1196), .Y(n_1273) );
INVx2_ASAP7_75t_SL g1260 ( .A(n_1207), .Y(n_1260) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1208), .Y(n_1258) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1215), .C(n_1218), .Y(n_1209) );
OAI21xp5_ASAP7_75t_SL g1219 ( .A1(n_1220), .A2(n_1224), .B(n_1230), .Y(n_1219) );
OAI21xp5_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1222), .B(n_1223), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1227), .B1(n_1228), .B2(n_1229), .Y(n_1224) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1226), .B(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1226), .Y(n_1310) );
NAND4xp25_ASAP7_75t_SL g1238 ( .A(n_1239), .B(n_1242), .C(n_1244), .D(n_1247), .Y(n_1238) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1321), .B1(n_1322), .B2(n_1412), .Y(n_1261) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1262), .Y(n_1412) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1264), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g1299 ( .A1(n_1266), .A2(n_1296), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1306), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1290), .B1(n_1291), .B2(n_1292), .Y(n_1288) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
OAI22xp33_ASAP7_75t_SL g1294 ( .A1(n_1295), .A2(n_1296), .B1(n_1297), .B2(n_1298), .Y(n_1294) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
OAI22x1_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1324), .B1(n_1370), .B2(n_1371), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1326), .Y(n_1369) );
NAND3xp33_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1333), .C(n_1336), .Y(n_1327) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NAND4xp25_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1356), .C(n_1361), .D(n_1365), .Y(n_1349) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_1371), .Y(n_1370) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
NAND4xp75_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1386), .C(n_1407), .D(n_1409), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1383), .Y(n_1374) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
OAI21xp5_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1396), .B(n_1406), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .Y(n_1387) );
OAI221xp5_ASAP7_75t_L g1413 ( .A1(n_1414), .A2(n_1662), .B1(n_1664), .B2(n_1702), .C(n_1706), .Y(n_1413) );
AOI211xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1570), .B(n_1612), .C(n_1644), .Y(n_1414) );
NAND5xp2_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1512), .C(n_1530), .D(n_1559), .E(n_1562), .Y(n_1415) );
AOI321xp33_ASAP7_75t_L g1416 ( .A1(n_1417), .A2(n_1459), .A3(n_1476), .B1(n_1483), .B2(n_1491), .C(n_1502), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1455), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1442), .Y(n_1419) );
CKINVDCx6p67_ASAP7_75t_R g1458 ( .A(n_1420), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1420), .B(n_1457), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1420), .B(n_1505), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1521 ( .A(n_1420), .B(n_1457), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1420), .B(n_1528), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1420), .B(n_1555), .Y(n_1565) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1420), .B(n_1506), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1420), .B(n_1443), .Y(n_1599) );
A2O1A1Ixp33_ASAP7_75t_SL g1648 ( .A1(n_1420), .A2(n_1649), .B(n_1653), .C(n_1655), .Y(n_1648) );
OR2x6_ASAP7_75t_SL g1420 ( .A(n_1421), .B(n_1432), .Y(n_1420) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1426), .Y(n_1423) );
AND2x4_ASAP7_75t_L g1430 ( .A(n_1424), .B(n_1427), .Y(n_1430) );
AND2x4_ASAP7_75t_L g1471 ( .A(n_1424), .B(n_1426), .Y(n_1471) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1425), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g1720 ( .A(n_1426), .Y(n_1720) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1428), .B(n_1437), .Y(n_1436) );
OAI22xp5_ASAP7_75t_L g1468 ( .A1(n_1429), .A2(n_1469), .B1(n_1470), .B2(n_1472), .Y(n_1468) );
INVx1_ASAP7_75t_SL g1429 ( .A(n_1430), .Y(n_1429) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1430), .Y(n_1482) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_1433), .A2(n_1438), .B1(n_1439), .B2(n_1441), .Y(n_1432) );
OAI22xp33_ASAP7_75t_L g1463 ( .A1(n_1433), .A2(n_1464), .B1(n_1465), .B2(n_1466), .Y(n_1463) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_1433), .A2(n_1439), .B1(n_1487), .B2(n_1488), .Y(n_1486) );
BUFx3_ASAP7_75t_L g1545 ( .A(n_1433), .Y(n_1545) );
BUFx6f_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_1434), .A2(n_1439), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1436), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_1435), .B(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1435), .Y(n_1447) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1436), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g1719 ( .A(n_1437), .Y(n_1719) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1439), .Y(n_1467) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1440), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1442), .B(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1442), .Y(n_1507) );
OAI32xp33_ASAP7_75t_L g1574 ( .A1(n_1442), .A2(n_1473), .A3(n_1513), .B1(n_1575), .B2(n_1577), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1442), .B(n_1458), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1442), .B(n_1517), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1451), .Y(n_1442) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1443), .Y(n_1457) );
OR2x2_ASAP7_75t_L g1506 ( .A(n_1443), .B(n_1451), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1443), .B(n_1529), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1450), .Y(n_1443) );
AND2x4_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
AND2x4_ASAP7_75t_L g1448 ( .A(n_1447), .B(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1451), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1451), .B(n_1458), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1451), .B(n_1457), .Y(n_1555) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_1455), .A2(n_1490), .B1(n_1532), .B2(n_1534), .C(n_1537), .Y(n_1531) );
O2A1O1Ixp33_ASAP7_75t_L g1593 ( .A1(n_1455), .A2(n_1557), .B(n_1594), .C(n_1595), .Y(n_1593) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
A2O1A1Ixp33_ASAP7_75t_L g1608 ( .A1(n_1456), .A2(n_1477), .B(n_1566), .C(n_1609), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1457), .B(n_1458), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1458), .B(n_1478), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1458), .B(n_1555), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1458), .B(n_1528), .Y(n_1561) );
NOR2xp33_ASAP7_75t_L g1576 ( .A(n_1458), .B(n_1478), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1458), .B(n_1529), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1458), .B(n_1500), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1458), .B(n_1529), .Y(n_1620) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1459), .B(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
OAI22xp5_ASAP7_75t_SL g1617 ( .A1(n_1460), .A2(n_1526), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1473), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1461), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1461), .Y(n_1496) );
INVx3_ASAP7_75t_L g1558 ( .A(n_1461), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1461), .B(n_1553), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1461), .B(n_1523), .Y(n_1604) );
AOI221xp5_ASAP7_75t_L g1621 ( .A1(n_1461), .A2(n_1622), .B1(n_1623), .B2(n_1625), .C(n_1629), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1461), .B(n_1473), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1461), .B(n_1511), .Y(n_1655) );
INVx3_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1462), .B(n_1498), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1462), .B(n_1473), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1468), .Y(n_1462) );
HB1xp67_ASAP7_75t_L g1547 ( .A(n_1466), .Y(n_1547) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1471), .Y(n_1541) );
BUFx3_ASAP7_75t_L g1663 ( .A(n_1471), .Y(n_1663) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1473), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1473), .B(n_1485), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1473), .B(n_1485), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1473), .B(n_1520), .Y(n_1519) );
OR2x2_ASAP7_75t_L g1525 ( .A(n_1473), .B(n_1523), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1473), .B(n_1523), .Y(n_1533) );
AND2x4_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1475), .Y(n_1473) );
NOR2x1_ASAP7_75t_L g1578 ( .A(n_1476), .B(n_1579), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1476), .B(n_1493), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1476), .B(n_1565), .Y(n_1584) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1476), .B(n_1525), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1476), .B(n_1583), .Y(n_1618) );
INVx2_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1477), .B(n_1536), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1477), .B(n_1552), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1564 ( .A(n_1477), .B(n_1565), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_1477), .B(n_1658), .Y(n_1657) );
INVx2_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx4_ASAP7_75t_L g1501 ( .A(n_1478), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1478), .B(n_1523), .Y(n_1522) );
OR2x2_ASAP7_75t_L g1573 ( .A(n_1478), .B(n_1506), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1478), .B(n_1553), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1640 ( .A(n_1478), .B(n_1552), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1478), .B(n_1527), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1654 ( .A(n_1478), .B(n_1569), .Y(n_1654) );
AND2x6_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1480), .Y(n_1478) );
INVx2_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_1482), .A2(n_1540), .B1(n_1541), .B2(n_1542), .Y(n_1539) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1483), .Y(n_1622) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1489), .Y(n_1483) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1484), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1484), .B(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1484), .Y(n_1626) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1484), .Y(n_1643) );
HB1xp67_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx2_ASAP7_75t_SL g1523 ( .A(n_1485), .Y(n_1523) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1490), .Y(n_1514) );
OAI22xp5_ASAP7_75t_L g1491 ( .A1(n_1492), .A2(n_1494), .B1(n_1496), .B2(n_1499), .Y(n_1491) );
INVxp67_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1493), .B(n_1501), .Y(n_1591) );
INVxp67_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1497), .Y(n_1495) );
AOI21xp5_ASAP7_75t_L g1607 ( .A1(n_1496), .A2(n_1515), .B(n_1537), .Y(n_1607) );
AOI22xp5_ASAP7_75t_L g1633 ( .A1(n_1496), .A2(n_1634), .B1(n_1637), .B2(n_1641), .Y(n_1633) );
OAI211xp5_ASAP7_75t_L g1570 ( .A1(n_1497), .A2(n_1571), .B(n_1582), .C(n_1596), .Y(n_1570) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVxp67_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1501), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1501), .B(n_1533), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1501), .B(n_1561), .Y(n_1560) );
AOI21xp5_ASAP7_75t_L g1502 ( .A1(n_1503), .A2(n_1507), .B(n_1508), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1503), .B(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
OAI31xp33_ASAP7_75t_L g1656 ( .A1(n_1504), .A2(n_1535), .A3(n_1657), .B(n_1659), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1505), .B(n_1517), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1505), .B(n_1576), .Y(n_1628) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1511), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1510), .B(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1510), .B(n_1528), .Y(n_1609) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1511), .Y(n_1611) );
AOI211xp5_ASAP7_75t_SL g1512 ( .A1(n_1513), .A2(n_1515), .B(n_1518), .C(n_1524), .Y(n_1512) );
OAI22xp5_ASAP7_75t_L g1597 ( .A1(n_1513), .A2(n_1598), .B1(n_1600), .B2(n_1601), .Y(n_1597) );
AOI21xp5_ASAP7_75t_L g1613 ( .A1(n_1513), .A2(n_1614), .B(n_1617), .Y(n_1613) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1515), .B(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1516), .B(n_1643), .Y(n_1642) );
INVxp67_ASAP7_75t_SL g1518 ( .A(n_1519), .Y(n_1518) );
INVxp33_ASAP7_75t_L g1630 ( .A(n_1520), .Y(n_1630) );
NOR2xp33_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1522), .Y(n_1520) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1521), .Y(n_1658) );
INVx2_ASAP7_75t_SL g1553 ( .A(n_1523), .Y(n_1553) );
NOR2xp33_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1526), .Y(n_1524) );
INVx2_ASAP7_75t_L g1583 ( .A(n_1525), .Y(n_1583) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
OAI21xp33_ASAP7_75t_SL g1590 ( .A1(n_1527), .A2(n_1591), .B(n_1592), .Y(n_1590) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1528), .Y(n_1651) );
OAI21xp5_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1548), .B(n_1556), .Y(n_1530) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1533), .Y(n_1600) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVxp67_ASAP7_75t_L g1601 ( .A(n_1536), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1537), .B(n_1557), .Y(n_1556) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_1538), .Y(n_1537) );
OR2x6_ASAP7_75t_SL g1538 ( .A(n_1539), .B(n_1543), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_1544), .A2(n_1545), .B1(n_1546), .B2(n_1547), .Y(n_1543) );
INVxp67_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1554), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
AOI221xp5_ASAP7_75t_L g1571 ( .A1(n_1553), .A2(n_1558), .B1(n_1572), .B2(n_1574), .C(n_1580), .Y(n_1571) );
NOR2xp33_ASAP7_75t_L g1580 ( .A(n_1553), .B(n_1581), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1553), .B(n_1573), .Y(n_1589) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1553), .Y(n_1661) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1555), .Y(n_1652) );
AOI211xp5_ASAP7_75t_L g1596 ( .A1(n_1557), .A2(n_1597), .B(n_1602), .C(n_1610), .Y(n_1596) );
NOR2xp33_ASAP7_75t_L g1639 ( .A(n_1557), .B(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_SL g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1561), .Y(n_1636) );
AOI21xp5_ASAP7_75t_L g1562 ( .A1(n_1563), .A2(n_1566), .B(n_1567), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
NOR2xp33_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1568), .Y(n_1592) );
NOR2xp33_ASAP7_75t_L g1610 ( .A(n_1569), .B(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
AOI211xp5_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1584), .B(n_1585), .C(n_1593), .Y(n_1582) );
OAI21xp33_ASAP7_75t_L g1585 ( .A1(n_1586), .A2(n_1588), .B(n_1590), .Y(n_1585) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVxp67_ASAP7_75t_SL g1588 ( .A(n_1589), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1595), .B(n_1638), .Y(n_1637) );
OAI211xp5_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1605), .B(n_1607), .C(n_1608), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
AOI21xp33_ASAP7_75t_SL g1629 ( .A1(n_1605), .A2(n_1630), .B(n_1631), .Y(n_1629) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
NAND3xp33_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1621), .C(n_1633), .Y(n_1612) );
INVxp67_ASAP7_75t_SL g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
INVxp67_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
INVxp67_ASAP7_75t_SL g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
OAI211xp5_ASAP7_75t_L g1644 ( .A1(n_1645), .A2(n_1647), .B(n_1648), .C(n_1656), .Y(n_1644) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1646), .B(n_1661), .Y(n_1660) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1652), .Y(n_1650) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
HB1xp67_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
HB1xp67_ASAP7_75t_L g1715 ( .A(n_1667), .Y(n_1715) );
NAND3xp33_ASAP7_75t_L g1668 ( .A(n_1669), .B(n_1673), .C(n_1676), .Y(n_1668) );
NAND4xp25_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1683), .C(n_1686), .D(n_1689), .Y(n_1679) );
INVx4_ASAP7_75t_SL g1702 ( .A(n_1703), .Y(n_1702) );
BUFx3_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
BUFx2_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
CKINVDCx5p33_ASAP7_75t_R g1708 ( .A(n_1709), .Y(n_1708) );
A2O1A1Ixp33_ASAP7_75t_L g1717 ( .A1(n_1710), .A2(n_1718), .B(n_1720), .C(n_1721), .Y(n_1717) );
INVxp33_ASAP7_75t_SL g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
HB1xp67_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
endmodule