module fake_ibex_579_n_2975 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_2975);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_2975;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2697;
wire n_2224;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_874;
wire n_1505;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2667;
wire n_2218;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2864;
wire n_1632;
wire n_2406;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2931;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_783;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_1365;
wire n_1472;
wire n_2802;
wire n_2443;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

INVx1_ASAP7_75t_L g632 ( 
.A(n_249),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_462),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_82),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_425),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_514),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_416),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_112),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_625),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_235),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_89),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_202),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_363),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_447),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_572),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_223),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_610),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_365),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_76),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_426),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_7),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_257),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_617),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_305),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_166),
.B(n_518),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_99),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_397),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_25),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_448),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_545),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_152),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_414),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_88),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_420),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_343),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_164),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_15),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_396),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_347),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_322),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_336),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_496),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_270),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_450),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_393),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_624),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_573),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_7),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_437),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_250),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_296),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_216),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_188),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_489),
.Y(n_686)
);

CKINVDCx16_ASAP7_75t_R g687 ( 
.A(n_83),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_200),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_60),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_114),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_41),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_125),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_613),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_592),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_512),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_124),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_502),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_142),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_37),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_300),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_281),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_11),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_79),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_259),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_331),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_216),
.B(n_265),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_590),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_292),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_147),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_485),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_373),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_448),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_587),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_327),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_93),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_508),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_236),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_419),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_128),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_110),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_518),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_278),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_612),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_402),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_567),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_470),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_103),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_534),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_84),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_129),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_66),
.Y(n_731)
);

BUFx5_ASAP7_75t_L g732 ( 
.A(n_407),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_444),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_283),
.Y(n_734)
);

BUFx5_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_469),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_437),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_124),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_505),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_42),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_349),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_556),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_474),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_609),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_166),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_251),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_9),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_21),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_474),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_505),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_267),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_72),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_312),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_45),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_196),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_280),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_430),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_605),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_421),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_524),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_628),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_606),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_619),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_473),
.Y(n_764)
);

XOR2xp5_ASAP7_75t_L g765 ( 
.A(n_467),
.B(n_489),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_446),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_472),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_279),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_167),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_615),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_153),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_78),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_571),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_210),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_475),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_557),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_542),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_31),
.B(n_95),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_33),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_339),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_334),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_318),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_435),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_59),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_507),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_620),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_321),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_500),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_598),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_333),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_468),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_136),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_285),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_52),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_135),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_158),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_86),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_6),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_600),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_183),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_436),
.Y(n_802)
);

BUFx5_ASAP7_75t_L g803 ( 
.A(n_404),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_348),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_284),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_589),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_597),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_137),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_386),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_447),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_577),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_149),
.Y(n_812)
);

BUFx8_ASAP7_75t_SL g813 ( 
.A(n_232),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_281),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_345),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_546),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_171),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_287),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_130),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_328),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_25),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_292),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_93),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_47),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_246),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_520),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_611),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_538),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_560),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_69),
.B(n_142),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_548),
.Y(n_831)
);

BUFx8_ASAP7_75t_SL g832 ( 
.A(n_154),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_509),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_582),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_578),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_99),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_461),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_389),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_332),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_541),
.Y(n_840)
);

CKINVDCx14_ASAP7_75t_R g841 ( 
.A(n_313),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_27),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_143),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_576),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_249),
.Y(n_845)
);

BUFx8_ASAP7_75t_SL g846 ( 
.A(n_276),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_195),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_471),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_533),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_495),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_19),
.Y(n_851)
);

BUFx8_ASAP7_75t_SL g852 ( 
.A(n_192),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_259),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_6),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_338),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_51),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_31),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_120),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_340),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_631),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_409),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_630),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_480),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_133),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_426),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_205),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_584),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_160),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_L g869 ( 
.A(n_514),
.B(n_486),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_140),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_472),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_247),
.Y(n_872)
);

BUFx8_ASAP7_75t_SL g873 ( 
.A(n_381),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_127),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_434),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_608),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_455),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_111),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_186),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_424),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_363),
.B(n_143),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_441),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_181),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_462),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_270),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_433),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_58),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_406),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_153),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_88),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_547),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_251),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_575),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_607),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_145),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_233),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_396),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_594),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_272),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_46),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_543),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_191),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_263),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_85),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_300),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_410),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_341),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_322),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_536),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_466),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_302),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_550),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_80),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_109),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_39),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_623),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_491),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_549),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_121),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_167),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_263),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_423),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_226),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_175),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_580),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_591),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_413),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_38),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_201),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_457),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_529),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_499),
.Y(n_932)
);

BUFx5_ASAP7_75t_L g933 ( 
.A(n_234),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_346),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_512),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_245),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_488),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_294),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_337),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_483),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_252),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_45),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_11),
.Y(n_943)
);

BUFx8_ASAP7_75t_SL g944 ( 
.A(n_61),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_432),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_181),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_261),
.Y(n_947)
);

BUFx2_ASAP7_75t_SL g948 ( 
.A(n_62),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_383),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_70),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_116),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_22),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_196),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_565),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_201),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_449),
.Y(n_956)
);

CKINVDCx14_ASAP7_75t_R g957 ( 
.A(n_227),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_77),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_402),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_341),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_139),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_41),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_149),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_77),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_57),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_221),
.B(n_5),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_245),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_256),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_479),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_238),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_172),
.Y(n_971)
);

CKINVDCx16_ASAP7_75t_R g972 ( 
.A(n_596),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_60),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_35),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_439),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_380),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_329),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_139),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_121),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_227),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_618),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_599),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_484),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_42),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_480),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_204),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_205),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_330),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_364),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_814),
.B(n_0),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_732),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_661),
.B(n_537),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_954),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_814),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_697),
.B(n_539),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_667),
.A2(n_544),
.B(n_540),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_732),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_821),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_851),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_732),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_732),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_661),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_851),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_742),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_841),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_756),
.Y(n_1006)
);

OA21x2_ASAP7_75t_L g1007 ( 
.A1(n_667),
.A2(n_552),
.B(n_551),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_756),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_SL g1009 ( 
.A1(n_642),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_875),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_900),
.B(n_4),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_957),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_732),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_967),
.A2(n_979),
.B1(n_897),
.B2(n_972),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_732),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_851),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_897),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_979),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_697),
.B(n_8),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_885),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_775),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_732),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_885),
.Y(n_1023)
);

BUFx8_ASAP7_75t_SL g1024 ( 
.A(n_813),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_954),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_775),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_690),
.B(n_946),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_742),
.Y(n_1028)
);

XNOR2x2_ASAP7_75t_L g1029 ( 
.A(n_656),
.B(n_8),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_823),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_857),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_803),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_803),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_954),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_803),
.Y(n_1035)
);

INVx6_ASAP7_75t_L g1036 ( 
.A(n_885),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_803),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_954),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_857),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_859),
.B(n_9),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_803),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_803),
.Y(n_1042)
);

AND2x6_ASAP7_75t_L g1043 ( 
.A(n_762),
.B(n_553),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_859),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_918),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_868),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_687),
.B(n_12),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_868),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_788),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_645),
.B(n_13),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_896),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_803),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_896),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_854),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_908),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_933),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_854),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_908),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_694),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_828),
.B(n_554),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_712),
.B(n_14),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_940),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_758),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_832),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_854),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_754),
.B(n_14),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_658),
.A2(n_16),
.B1(n_10),
.B2(n_15),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_940),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_658),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_662),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_678),
.A2(n_558),
.B(n_555),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_850),
.B(n_21),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_828),
.B(n_559),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_854),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_965),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_933),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_662),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_933),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_965),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_864),
.B(n_23),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_892),
.B(n_24),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_640),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_663),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_685),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_960),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_663),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_664),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_678),
.A2(n_562),
.B(n_561),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_685),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_960),
.Y(n_1091)
);

OAI22x1_ASAP7_75t_L g1092 ( 
.A1(n_765),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_744),
.A2(n_566),
.B(n_564),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_694),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_971),
.B(n_29),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_758),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_664),
.B(n_29),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_L g1098 ( 
.A(n_992),
.B(n_735),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_991),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_990),
.B(n_744),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_991),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_997),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_996),
.A2(n_646),
.B(n_639),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_992),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_997),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1003),
.B(n_1023),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_990),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1000),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1000),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1001),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_992),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1044),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1086),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1053),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1003),
.B(n_679),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1013),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1013),
.B(n_790),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1015),
.B(n_816),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1053),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1015),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_1088),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1023),
.B(n_707),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1077),
.A2(n_655),
.B1(n_659),
.B2(n_651),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1022),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1022),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1036),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1019),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_998),
.B(n_672),
.Y(n_1128)
);

INVxp33_ASAP7_75t_L g1129 ( 
.A(n_1088),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1032),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1012),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1033),
.B(n_891),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1040),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1025),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1033),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1035),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1006),
.Y(n_1137)
);

AO22x2_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_830),
.B1(n_948),
.B2(n_633),
.Y(n_1138)
);

INVx6_ASAP7_75t_L g1139 ( 
.A(n_1036),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_1014),
.B(n_989),
.C(n_988),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1008),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1039),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1005),
.B(n_665),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1018),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1039),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1041),
.A2(n_981),
.B(n_891),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1005),
.B(n_1058),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1042),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1068),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1045),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1010),
.B(n_668),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1010),
.B(n_668),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1068),
.B(n_669),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1042),
.B(n_981),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1059),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_994),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1052),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1027),
.B(n_676),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1052),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_992),
.A2(n_635),
.B1(n_638),
.B2(n_632),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1056),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1021),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_992),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1076),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_999),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1076),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1078),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1016),
.A2(n_770),
.B1(n_786),
.B2(n_763),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1002),
.B(n_672),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1020),
.B(n_648),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1026),
.Y(n_1174)
);

INVx8_ASAP7_75t_L g1175 ( 
.A(n_999),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1030),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1004),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_SL g1178 ( 
.A(n_1047),
.B(n_763),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1049),
.A2(n_676),
.B1(n_683),
.B2(n_673),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1078),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1087),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1028),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_1007),
.B(n_696),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1011),
.B(n_683),
.C(n_673),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1087),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1025),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1050),
.A2(n_1066),
.B(n_1061),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1031),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_995),
.B(n_735),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1046),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1048),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1051),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1024),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1025),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1063),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1055),
.B(n_688),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1059),
.B(n_691),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1043),
.Y(n_1198)
);

INVx8_ASAP7_75t_L g1199 ( 
.A(n_1094),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1062),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1075),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1097),
.B(n_691),
.C(n_689),
.Y(n_1202)
);

NOR2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_689),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_993),
.B(n_735),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1034),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1038),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1094),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1072),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1038),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1038),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1082),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1084),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1038),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1090),
.B(n_692),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1024),
.Y(n_1215)
);

INVxp33_ASAP7_75t_L g1216 ( 
.A(n_1080),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1054),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1092),
.B(n_1067),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1069),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1095),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1054),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_993),
.B(n_735),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1081),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1054),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1064),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_993),
.B(n_735),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1007),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1057),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1057),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_L g1231 ( 
.A(n_1043),
.B(n_735),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1017),
.B(n_910),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1065),
.Y(n_1233)
);

BUFx10_ASAP7_75t_L g1234 ( 
.A(n_1043),
.Y(n_1234)
);

BUFx10_ASAP7_75t_L g1235 ( 
.A(n_1043),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_SL g1236 ( 
.A(n_1043),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1060),
.Y(n_1237)
);

CKINVDCx11_ASAP7_75t_R g1238 ( 
.A(n_1070),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_1060),
.Y(n_1239)
);

INVx8_ASAP7_75t_L g1240 ( 
.A(n_1060),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1060),
.Y(n_1241)
);

BUFx4f_ASAP7_75t_L g1242 ( 
.A(n_1060),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1074),
.Y(n_1243)
);

AND3x2_ASAP7_75t_L g1244 ( 
.A(n_1029),
.B(n_968),
.C(n_719),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1083),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1085),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1091),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1073),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1073),
.B(n_695),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1073),
.A2(n_700),
.B1(n_703),
.B2(n_695),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1091),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1073),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1071),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1071),
.B(n_703),
.C(n_700),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1071),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1089),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1089),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1089),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1093),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1093),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1093),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1079),
.B(n_729),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1079),
.B(n_904),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_990),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1137),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1141),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_1129),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1221),
.B(n_1224),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1237),
.B(n_1248),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1208),
.B(n_800),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_SL g1272 ( 
.A(n_1248),
.B(n_770),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1216),
.B(n_909),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1166),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1187),
.B(n_909),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1216),
.B(n_912),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1177),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

AND2x6_ASAP7_75t_L g1279 ( 
.A(n_1166),
.B(n_831),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1175),
.B(n_706),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1187),
.B(n_912),
.Y(n_1281)
);

NOR3xp33_ASAP7_75t_L g1282 ( 
.A(n_1123),
.B(n_701),
.C(n_671),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1113),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1147),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_L g1285 ( 
.A(n_1240),
.B(n_926),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_SL g1286 ( 
.A(n_1129),
.B(n_786),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1148),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1161),
.A2(n_835),
.B1(n_905),
.B2(n_904),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1142),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1126),
.B(n_693),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1152),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_SL g1292 ( 
.A(n_1240),
.B(n_835),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1219),
.A2(n_906),
.B1(n_910),
.B2(n_905),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1163),
.B(n_911),
.C(n_906),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1150),
.B(n_1106),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1265),
.B(n_654),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1121),
.A2(n_914),
.B1(n_919),
.B2(n_911),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1107),
.B(n_916),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1142),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1198),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1127),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1175),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1131),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1128),
.B(n_921),
.Y(n_1304)
);

NAND2xp33_ASAP7_75t_L g1305 ( 
.A(n_1240),
.B(n_713),
.Y(n_1305)
);

NOR3xp33_ASAP7_75t_L g1306 ( 
.A(n_1123),
.B(n_743),
.C(n_708),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1172),
.B(n_725),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1154),
.B(n_914),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1127),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1156),
.B(n_777),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1211),
.Y(n_1311)
);

OA22x2_ASAP7_75t_L g1312 ( 
.A1(n_1244),
.A2(n_920),
.B1(n_921),
.B2(n_919),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1155),
.B(n_807),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1212),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1149),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1175),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1165),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1159),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1199),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1115),
.B(n_840),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1140),
.A2(n_923),
.B1(n_928),
.B2(n_920),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1174),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1198),
.B(n_1253),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1176),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1104),
.B(n_1111),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1115),
.B(n_844),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1144),
.B(n_936),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1242),
.B(n_860),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1188),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1190),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1122),
.B(n_867),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1249),
.A2(n_644),
.B1(n_647),
.B2(n_643),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1122),
.B(n_898),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1199),
.B(n_778),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1199),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1139),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1168),
.B(n_928),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1191),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1133),
.B(n_1112),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1139),
.B(n_982),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1192),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1114),
.B(n_931),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1119),
.B(n_723),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1100),
.B(n_761),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1201),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1232),
.A2(n_931),
.B1(n_932),
.B2(n_923),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1163),
.A2(n_653),
.B1(n_657),
.B2(n_650),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1173),
.B(n_932),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1099),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1158),
.Y(n_1351)
);

NOR3xp33_ASAP7_75t_L g1352 ( 
.A(n_1171),
.B(n_805),
.C(n_768),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1214),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1173),
.B(n_934),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1250),
.B(n_1241),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1263),
.B(n_934),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1179),
.A2(n_666),
.B(n_670),
.C(n_660),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1264),
.B(n_773),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1099),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1101),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1196),
.B(n_936),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1197),
.B(n_1207),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1255),
.B(n_949),
.C(n_941),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1202),
.B(n_949),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1219),
.A2(n_709),
.B1(n_731),
.B2(n_686),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1184),
.B(n_776),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_SL g1367 ( 
.A(n_1153),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1101),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1153),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1183),
.B(n_787),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1203),
.B(n_869),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1102),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1226),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1245),
.B(n_806),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1193),
.B(n_951),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1183),
.B(n_811),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1102),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1105),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1117),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1105),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1108),
.B(n_827),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1109),
.B(n_829),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1215),
.B(n_951),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1110),
.B(n_834),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1118),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1245),
.A2(n_953),
.B1(n_955),
.B2(n_952),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1189),
.B(n_862),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1116),
.B(n_876),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1118),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1120),
.B(n_893),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1189),
.B(n_674),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1178),
.B(n_894),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1236),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1178),
.B(n_901),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1234),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1124),
.B(n_925),
.Y(n_1397)
);

NOR2xp67_ASAP7_75t_L g1398 ( 
.A(n_1204),
.B(n_952),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1138),
.B(n_881),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1257),
.B(n_634),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1098),
.A2(n_677),
.B1(n_680),
.B2(n_675),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1124),
.B(n_953),
.Y(n_1402)
);

NOR3xp33_ASAP7_75t_L g1403 ( 
.A(n_1220),
.B(n_947),
.C(n_839),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1103),
.B(n_966),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1195),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1125),
.B(n_955),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1235),
.B(n_1239),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1125),
.B(n_956),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1130),
.B(n_956),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1231),
.B(n_637),
.C(n_636),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1132),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1257),
.B(n_641),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1157),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1130),
.B(n_726),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1254),
.A2(n_682),
.B(n_681),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1235),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1204),
.B(n_30),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1138),
.B(n_649),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1239),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1239),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1135),
.B(n_652),
.Y(n_1421)
);

O2A1O1Ixp5_ASAP7_75t_L g1422 ( 
.A1(n_1228),
.A2(n_733),
.B(n_740),
.C(n_728),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1136),
.B(n_705),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1138),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1257),
.B(n_714),
.Y(n_1425)
);

INVx8_ASAP7_75t_L g1426 ( 
.A(n_1257),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_L g1427 ( 
.A(n_1223),
.B(n_30),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1260),
.B(n_718),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1143),
.B(n_720),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1261),
.B(n_721),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1259),
.A2(n_686),
.B1(n_731),
.B2(n_709),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1223),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1145),
.B(n_728),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1227),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1145),
.B(n_733),
.Y(n_1435)
);

AO22x2_ASAP7_75t_L g1436 ( 
.A1(n_1220),
.A2(n_767),
.B1(n_799),
.B2(n_764),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1146),
.B(n_724),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1227),
.B(n_32),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1151),
.B(n_730),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1195),
.B(n_736),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1160),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1162),
.B(n_737),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1259),
.A2(n_698),
.B1(n_699),
.B2(n_684),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1164),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1256),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1167),
.B(n_740),
.Y(n_1447)
);

NOR3xp33_ASAP7_75t_L g1448 ( 
.A(n_1238),
.B(n_739),
.C(n_738),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_R g1449 ( 
.A(n_1238),
.B(n_977),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1262),
.A2(n_767),
.B1(n_799),
.B2(n_764),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1169),
.B(n_741),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1170),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1180),
.B(n_745),
.Y(n_1453)
);

AND2x2_ASAP7_75t_SL g1454 ( 
.A(n_1258),
.B(n_846),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1181),
.B(n_746),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1181),
.B(n_1185),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1262),
.B(n_748),
.C(n_747),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1185),
.B(n_750),
.Y(n_1458)
);

BUFx5_ASAP7_75t_L g1459 ( 
.A(n_1225),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1233),
.B(n_751),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1243),
.B(n_752),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1246),
.B(n_753),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1247),
.B(n_757),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1251),
.B(n_759),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_1252),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1217),
.B(n_766),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1134),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1218),
.A2(n_704),
.B(n_710),
.C(n_702),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1210),
.B(n_769),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1186),
.B(n_855),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1194),
.B(n_855),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1194),
.B(n_861),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1218),
.A2(n_715),
.B1(n_716),
.B2(n_711),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1222),
.A2(n_722),
.B1(n_727),
.B2(n_717),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1210),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1229),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1283),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1269),
.B(n_781),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1269),
.B(n_782),
.Y(n_1479)
);

AO22x1_ASAP7_75t_L g1480 ( 
.A1(n_1431),
.A2(n_815),
.B1(n_824),
.B2(n_802),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1295),
.B(n_783),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1303),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1415),
.A2(n_749),
.B(n_755),
.C(n_734),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1268),
.B(n_852),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1328),
.B(n_784),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1440),
.A2(n_771),
.B(n_760),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1415),
.A2(n_774),
.B(n_779),
.C(n_772),
.Y(n_1487)
);

AOI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1355),
.A2(n_1315),
.B(n_1370),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1266),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1404),
.A2(n_785),
.B(n_780),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1442),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1442),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1267),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1293),
.A2(n_791),
.B(n_792),
.C(n_789),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1271),
.B(n_798),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1422),
.A2(n_794),
.B(n_793),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1353),
.B(n_810),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1284),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1323),
.Y(n_1499)
);

O2A1O1Ixp5_ASAP7_75t_L g1500 ( 
.A1(n_1404),
.A2(n_888),
.B(n_903),
.C(n_879),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1451),
.B(n_817),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1272),
.A2(n_819),
.B(n_818),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1376),
.A2(n_1281),
.B(n_1275),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1316),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1458),
.B(n_1273),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1362),
.B(n_873),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1428),
.A2(n_796),
.B(n_797),
.C(n_795),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1276),
.B(n_822),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1323),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1323),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1325),
.A2(n_1206),
.B(n_1205),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1402),
.B(n_836),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1314),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1430),
.A2(n_804),
.B(n_808),
.C(n_801),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1352),
.B(n_843),
.C(n_842),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1373),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1274),
.B(n_845),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1357),
.A2(n_812),
.B(n_820),
.C(n_809),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1319),
.Y(n_1519)
);

AO32x1_ASAP7_75t_L g1520 ( 
.A1(n_1434),
.A2(n_903),
.A3(n_907),
.B1(n_888),
.B2(n_879),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1337),
.B(n_944),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1301),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1308),
.B(n_815),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1275),
.A2(n_1281),
.B(n_1270),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1402),
.B(n_848),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1323),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1444),
.A2(n_847),
.B1(n_866),
.B2(n_824),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_L g1528 ( 
.A(n_1302),
.B(n_32),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1304),
.B(n_847),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1381),
.A2(n_1209),
.B(n_1230),
.Y(n_1530)
);

AOI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1400),
.A2(n_1425),
.B(n_1412),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1406),
.B(n_856),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1274),
.B(n_863),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1335),
.B(n_33),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1274),
.B(n_865),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1327),
.B(n_866),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1288),
.B(n_874),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1300),
.B(n_871),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1393),
.A2(n_826),
.B(n_833),
.C(n_825),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1309),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1294),
.A2(n_878),
.B1(n_887),
.B2(n_874),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1369),
.B(n_837),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1300),
.B(n_872),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1406),
.B(n_1408),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_R g1545 ( 
.A(n_1286),
.B(n_878),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1383),
.A2(n_1407),
.B(n_1456),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1351),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1289),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1343),
.B(n_924),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1318),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1426),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1347),
.B(n_924),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1408),
.B(n_880),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1300),
.B(n_882),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1292),
.A2(n_886),
.B1(n_902),
.B2(n_884),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1426),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1324),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1282),
.A2(n_849),
.B(n_853),
.C(n_838),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1348),
.A2(n_1332),
.B1(n_1339),
.B2(n_1401),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1409),
.A2(n_1213),
.B(n_870),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1409),
.A2(n_877),
.B(n_858),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1317),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1356),
.B(n_942),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1339),
.A2(n_977),
.B1(n_942),
.B2(n_883),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1292),
.A2(n_970),
.B1(n_976),
.B2(n_962),
.Y(n_1565)
);

OAI21xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1311),
.A2(n_890),
.B(n_889),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1374),
.B(n_978),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1441),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1329),
.B(n_980),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1330),
.B(n_983),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1387),
.A2(n_984),
.B1(n_895),
.B2(n_899),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1367),
.Y(n_1572)
);

AO21x1_ASAP7_75t_L g1573 ( 
.A1(n_1388),
.A2(n_915),
.B(n_913),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1431),
.Y(n_1574)
);

BUFx4f_ASAP7_75t_L g1575 ( 
.A(n_1399),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1450),
.B(n_917),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1395),
.A2(n_922),
.B(n_929),
.C(n_927),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1405),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1365),
.A2(n_963),
.B1(n_964),
.B2(n_961),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1297),
.A2(n_930),
.B1(n_938),
.B2(n_935),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1338),
.B(n_1342),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1363),
.B(n_945),
.C(n_939),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1346),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1349),
.A2(n_958),
.B1(n_959),
.B2(n_950),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1365),
.B(n_969),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1336),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1358),
.B(n_973),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1358),
.B(n_974),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1354),
.A2(n_985),
.B1(n_987),
.B2(n_975),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1344),
.B(n_907),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1322),
.B(n_937),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1457),
.A2(n_986),
.B(n_943),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1306),
.B(n_34),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1466),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1379),
.A2(n_629),
.B(n_627),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1454),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1445),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1361),
.B(n_36),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1341),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1366),
.B(n_37),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1410),
.A2(n_570),
.B(n_569),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_L g1602 ( 
.A(n_1424),
.B(n_38),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1298),
.B(n_39),
.Y(n_1603)
);

CKINVDCx16_ASAP7_75t_R g1604 ( 
.A(n_1367),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1386),
.A2(n_579),
.B(n_574),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1390),
.A2(n_583),
.B(n_581),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1394),
.B(n_40),
.Y(n_1607)
);

NOR2x1p5_ASAP7_75t_SL g1608 ( 
.A(n_1459),
.B(n_585),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1298),
.B(n_43),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1416),
.A2(n_593),
.B(n_586),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1321),
.A2(n_43),
.B(n_44),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1296),
.B(n_1345),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1468),
.A2(n_48),
.B(n_44),
.C(n_47),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1398),
.B(n_1313),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1299),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1312),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1296),
.B(n_49),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1277),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1396),
.B(n_595),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1280),
.B(n_53),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1287),
.B(n_54),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1291),
.B(n_54),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1279),
.Y(n_1623)
);

AO21x1_ASAP7_75t_L g1624 ( 
.A1(n_1381),
.A2(n_55),
.B(n_56),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1414),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1364),
.B(n_55),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1414),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1452),
.A2(n_602),
.B(n_601),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1413),
.A2(n_604),
.B(n_603),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1433),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1399),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1310),
.B(n_61),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1320),
.B(n_63),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1307),
.B(n_63),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1326),
.B(n_64),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1433),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1280),
.B(n_64),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1350),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1359),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1331),
.B(n_65),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1333),
.B(n_65),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1299),
.B(n_1421),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1360),
.A2(n_1372),
.B(n_1368),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1382),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1382),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1377),
.A2(n_616),
.B(n_614),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1423),
.B(n_70),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1446),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1278),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1429),
.B(n_73),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1334),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1652)
);

O2A1O1Ixp5_ASAP7_75t_L g1653 ( 
.A1(n_1469),
.A2(n_622),
.B(n_626),
.C(n_621),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1446),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1443),
.B(n_1453),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1385),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1455),
.B(n_75),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1435),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1378),
.A2(n_80),
.B(n_81),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1396),
.B(n_83),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1385),
.B(n_85),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1411),
.A2(n_86),
.B(n_87),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1435),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1462),
.A2(n_89),
.B(n_90),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1463),
.A2(n_90),
.B(n_91),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1389),
.B(n_91),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1391),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1380),
.A2(n_92),
.B(n_94),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1399),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1391),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1397),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1312),
.A2(n_1418),
.B1(n_1371),
.B2(n_1285),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1436),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1436),
.B(n_104),
.Y(n_1674)
);

O2A1O1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1403),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1447),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1447),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1473),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1432),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_1679)
);

AO21x1_ASAP7_75t_L g1680 ( 
.A1(n_1470),
.A2(n_122),
.B(n_123),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1419),
.B(n_125),
.Y(n_1681)
);

NOR2x1p5_ASAP7_75t_SL g1682 ( 
.A(n_1459),
.B(n_126),
.Y(n_1682)
);

BUFx4f_ASAP7_75t_L g1683 ( 
.A(n_1334),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1420),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1470),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1305),
.A2(n_128),
.B(n_129),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1371),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1392),
.A2(n_131),
.B(n_132),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1417),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_1689)
);

BUFx4f_ASAP7_75t_L g1690 ( 
.A(n_1334),
.Y(n_1690)
);

INVxp33_ASAP7_75t_SL g1691 ( 
.A(n_1449),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1290),
.A2(n_1448),
.B1(n_1340),
.B2(n_1384),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1474),
.A2(n_140),
.B1(n_137),
.B2(n_138),
.Y(n_1693)
);

BUFx12f_ASAP7_75t_L g1694 ( 
.A(n_1279),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1375),
.B(n_141),
.C(n_144),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1427),
.A2(n_145),
.B1(n_141),
.B2(n_144),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1471),
.A2(n_146),
.B(n_147),
.Y(n_1697)
);

AOI221x1_ASAP7_75t_L g1698 ( 
.A1(n_1471),
.A2(n_150),
.B1(n_146),
.B2(n_148),
.C(n_151),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1438),
.A2(n_154),
.B1(n_151),
.B2(n_152),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1472),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1467),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1472),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1460),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1476),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1459),
.B(n_156),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1475),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1475),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1459),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1465),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1465),
.B(n_165),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1269),
.B(n_168),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1269),
.B(n_169),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1269),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1269),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1269),
.B(n_173),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1597),
.A2(n_177),
.B1(n_174),
.B2(n_176),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1559),
.B(n_176),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1551),
.Y(n_1719)
);

NAND3x1_ASAP7_75t_L g1720 ( 
.A(n_1674),
.B(n_1672),
.C(n_1616),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1594),
.B(n_1478),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1594),
.B(n_1489),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1597),
.B(n_178),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1654),
.B(n_179),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1537),
.B(n_179),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_R g1726 ( 
.A(n_1572),
.B(n_180),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_SL g1727 ( 
.A(n_1607),
.B(n_180),
.Y(n_1727)
);

AO221x1_ASAP7_75t_L g1728 ( 
.A1(n_1564),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.C(n_185),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1551),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1493),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1625),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1524),
.A2(n_186),
.B(n_187),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1530),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1710),
.B(n_189),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1598),
.B(n_189),
.C(n_190),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1646),
.A2(n_1628),
.B(n_1653),
.Y(n_1737)
);

AO21x1_ASAP7_75t_L g1738 ( 
.A1(n_1628),
.A2(n_190),
.B(n_191),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1544),
.A2(n_192),
.B(n_193),
.Y(n_1739)
);

INVx3_ASAP7_75t_SL g1740 ( 
.A(n_1604),
.Y(n_1740)
);

O2A1O1Ixp5_ASAP7_75t_L g1741 ( 
.A1(n_1531),
.A2(n_197),
.B(n_194),
.C(n_195),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1530),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1549),
.B(n_194),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1546),
.A2(n_197),
.B(n_198),
.Y(n_1744)
);

BUFx12f_ASAP7_75t_L g1745 ( 
.A(n_1607),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1545),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1498),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1654),
.B(n_199),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_SL g1749 ( 
.A1(n_1623),
.A2(n_199),
.B(n_200),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1652),
.A2(n_202),
.B(n_203),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1574),
.B(n_203),
.Y(n_1751)
);

O2A1O1Ixp5_ASAP7_75t_L g1752 ( 
.A1(n_1680),
.A2(n_1624),
.B(n_1706),
.C(n_1601),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1655),
.A2(n_204),
.B(n_206),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1550),
.B(n_207),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1557),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1558),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1646),
.A2(n_211),
.B(n_212),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1581),
.A2(n_1612),
.B(n_1643),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1643),
.A2(n_212),
.B(n_213),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1505),
.A2(n_213),
.B(n_214),
.Y(n_1760)
);

OAI21xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1627),
.A2(n_214),
.B(n_215),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1482),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1630),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1516),
.Y(n_1764)
);

NOR4xp25_ASAP7_75t_L g1765 ( 
.A(n_1631),
.B(n_1669),
.C(n_1675),
.D(n_1645),
.Y(n_1765)
);

NAND2x1_ASAP7_75t_L g1766 ( 
.A(n_1551),
.B(n_218),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1583),
.B(n_219),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1636),
.B(n_220),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1658),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1556),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1547),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1663),
.A2(n_222),
.B(n_223),
.Y(n_1772)
);

O2A1O1Ixp5_ASAP7_75t_L g1773 ( 
.A1(n_1601),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1500),
.A2(n_225),
.B(n_228),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1713),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1556),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1556),
.Y(n_1777)
);

OAI21x1_ASAP7_75t_L g1778 ( 
.A1(n_1595),
.A2(n_229),
.B(n_230),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1523),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1638),
.Y(n_1781)
);

AO31x2_ASAP7_75t_L g1782 ( 
.A1(n_1698),
.A2(n_235),
.A3(n_231),
.B(n_233),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1536),
.B(n_236),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1491),
.B(n_237),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1605),
.A2(n_238),
.B(n_239),
.Y(n_1785)
);

OAI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1606),
.A2(n_239),
.B(n_240),
.Y(n_1786)
);

OAI22x1_ASAP7_75t_L g1787 ( 
.A1(n_1673),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1576),
.B(n_241),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1568),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1716),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1584),
.B(n_246),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1702),
.A2(n_252),
.B1(n_248),
.B2(n_250),
.Y(n_1792)
);

AO31x2_ASAP7_75t_L g1793 ( 
.A1(n_1573),
.A2(n_254),
.A3(n_248),
.B(n_253),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1599),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1685),
.Y(n_1795)
);

OAI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1629),
.A2(n_253),
.B(n_254),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1529),
.A2(n_260),
.B1(n_255),
.B2(n_258),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1496),
.A2(n_258),
.B(n_260),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1491),
.Y(n_1799)
);

OAI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1496),
.A2(n_261),
.B(n_262),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1589),
.B(n_262),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1499),
.B(n_264),
.Y(n_1802)
);

OAI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1563),
.A2(n_264),
.B(n_265),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1684),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1642),
.A2(n_266),
.B(n_268),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1539),
.B(n_269),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1577),
.B(n_271),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1681),
.B(n_273),
.C(n_274),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1504),
.B(n_275),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1560),
.A2(n_275),
.B(n_276),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1495),
.A2(n_277),
.B(n_279),
.Y(n_1812)
);

AO31x2_ASAP7_75t_L g1813 ( 
.A1(n_1483),
.A2(n_283),
.A3(n_280),
.B(n_282),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1691),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1497),
.B(n_282),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1659),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1555),
.A2(n_286),
.B(n_288),
.Y(n_1817)
);

O2A1O1Ixp5_ASAP7_75t_SL g1818 ( 
.A1(n_1696),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1487),
.B(n_289),
.Y(n_1819)
);

INVx3_ASAP7_75t_SL g1820 ( 
.A(n_1504),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1542),
.Y(n_1821)
);

AO31x2_ASAP7_75t_L g1822 ( 
.A1(n_1613),
.A2(n_293),
.A3(n_290),
.B(n_291),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1513),
.Y(n_1823)
);

CKINVDCx12_ASAP7_75t_R g1824 ( 
.A(n_1585),
.Y(n_1824)
);

NOR3xp33_ASAP7_75t_L g1825 ( 
.A(n_1494),
.B(n_293),
.C(n_294),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1481),
.B(n_295),
.Y(n_1826)
);

AO21x1_ASAP7_75t_L g1827 ( 
.A1(n_1659),
.A2(n_297),
.B(n_298),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_SL g1828 ( 
.A1(n_1668),
.A2(n_297),
.B(n_298),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_SL g1829 ( 
.A1(n_1668),
.A2(n_299),
.B(n_301),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1587),
.B(n_299),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1683),
.B(n_1690),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1567),
.B(n_302),
.Y(n_1832)
);

BUFx2_ASAP7_75t_SL g1833 ( 
.A(n_1519),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1638),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1639),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1639),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1578),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1588),
.B(n_306),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1614),
.A2(n_307),
.B(n_308),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1561),
.B(n_308),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1580),
.B(n_309),
.Y(n_1841)
);

AO31x2_ASAP7_75t_L g1842 ( 
.A1(n_1676),
.A2(n_1677),
.A3(n_1656),
.B(n_1667),
.Y(n_1842)
);

OAI21xp33_ASAP7_75t_L g1843 ( 
.A1(n_1501),
.A2(n_310),
.B(n_311),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1512),
.A2(n_311),
.B(n_312),
.Y(n_1844)
);

AOI211x1_ASAP7_75t_L g1845 ( 
.A1(n_1486),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_SL g1846 ( 
.A1(n_1686),
.A2(n_314),
.B(n_315),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1542),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1700),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1562),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1525),
.A2(n_319),
.B(n_320),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1683),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1571),
.B(n_323),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1492),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1532),
.B(n_324),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1553),
.B(n_324),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1518),
.B(n_325),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1591),
.Y(n_1857)
);

AOI221x1_ASAP7_75t_L g1858 ( 
.A1(n_1611),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.C(n_329),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1592),
.A2(n_335),
.B(n_336),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1486),
.B(n_335),
.Y(n_1860)
);

AO31x2_ASAP7_75t_L g1861 ( 
.A1(n_1644),
.A2(n_339),
.A3(n_337),
.B(n_338),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1592),
.A2(n_340),
.B(n_342),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1661),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1633),
.A2(n_344),
.B(n_345),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1569),
.B(n_346),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1666),
.A2(n_347),
.B(n_348),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1621),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1570),
.B(n_349),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1519),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_SL g1870 ( 
.A(n_1690),
.B(n_350),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1541),
.B(n_350),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1635),
.A2(n_351),
.B(n_352),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1682),
.A2(n_351),
.B(n_352),
.C(n_353),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1506),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_L g1875 ( 
.A(n_1515),
.B(n_354),
.C(n_355),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1640),
.A2(n_356),
.B(n_357),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1647),
.A2(n_356),
.B(n_357),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1582),
.A2(n_358),
.B(n_359),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1704),
.B(n_360),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1650),
.A2(n_360),
.B(n_361),
.Y(n_1880)
);

OAI21x1_ASAP7_75t_SL g1881 ( 
.A1(n_1622),
.A2(n_362),
.B(n_366),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1704),
.B(n_1566),
.Y(n_1882)
);

AOI211x1_ASAP7_75t_L g1883 ( 
.A1(n_1678),
.A2(n_1712),
.B(n_1645),
.C(n_1714),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1522),
.Y(n_1884)
);

AO31x2_ASAP7_75t_L g1885 ( 
.A1(n_1670),
.A2(n_366),
.A3(n_367),
.B(n_368),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1484),
.B(n_367),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1590),
.B(n_368),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1586),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1603),
.B(n_369),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1609),
.B(n_369),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1540),
.B(n_370),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1641),
.A2(n_371),
.B(n_372),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1479),
.A2(n_374),
.B(n_375),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1617),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_SL g1895 ( 
.A1(n_1600),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.C(n_378),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1692),
.B(n_376),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1657),
.A2(n_377),
.B(n_378),
.Y(n_1897)
);

AO31x2_ASAP7_75t_L g1898 ( 
.A1(n_1671),
.A2(n_379),
.A3(n_380),
.B(n_381),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1508),
.B(n_382),
.Y(n_1899)
);

AO31x2_ASAP7_75t_L g1900 ( 
.A1(n_1705),
.A2(n_384),
.A3(n_385),
.B(n_386),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1593),
.B(n_384),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1626),
.A2(n_385),
.B(n_387),
.Y(n_1902)
);

CKINVDCx8_ASAP7_75t_R g1903 ( 
.A(n_1620),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1694),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1490),
.B(n_1703),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1618),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1664),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1490),
.B(n_390),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1565),
.B(n_391),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1509),
.B(n_391),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1509),
.B(n_392),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1665),
.A2(n_392),
.B(n_393),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1649),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1502),
.A2(n_394),
.B1(n_395),
.B2(n_398),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1521),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.C(n_401),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1678),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_SL g1917 ( 
.A(n_1660),
.B(n_403),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1510),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1637),
.B(n_405),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1632),
.A2(n_405),
.B(n_406),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1649),
.Y(n_1921)
);

AO21x1_ASAP7_75t_L g1922 ( 
.A1(n_1696),
.A2(n_407),
.B(n_408),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_SL g1923 ( 
.A1(n_1596),
.A2(n_408),
.B(n_409),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1510),
.A2(n_410),
.B(n_411),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1697),
.A2(n_411),
.B(n_412),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1693),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1708),
.Y(n_1927)
);

AOI211x1_ASAP7_75t_L g1928 ( 
.A1(n_1688),
.A2(n_415),
.B(n_416),
.C(n_417),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1526),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1602),
.B(n_418),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1634),
.A2(n_418),
.B(n_419),
.Y(n_1931)
);

OAI21x1_ASAP7_75t_L g1932 ( 
.A1(n_1548),
.A2(n_420),
.B(n_421),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1526),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1651),
.B(n_422),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1701),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1575),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1615),
.B(n_427),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1528),
.B(n_428),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1679),
.A2(n_429),
.B(n_430),
.C(n_431),
.Y(n_1939)
);

A2O1A1Ixp33_ASAP7_75t_L g1940 ( 
.A1(n_1662),
.A2(n_431),
.B(n_432),
.C(n_433),
.Y(n_1940)
);

OA22x2_ASAP7_75t_L g1941 ( 
.A1(n_1687),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1534),
.B(n_438),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1485),
.A2(n_438),
.B(n_439),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1517),
.A2(n_440),
.B(n_441),
.Y(n_1944)
);

AO31x2_ASAP7_75t_L g1945 ( 
.A1(n_1689),
.A2(n_442),
.A3(n_443),
.B(n_444),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1533),
.A2(n_1538),
.B(n_1554),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1648),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1535),
.A2(n_442),
.B(n_443),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1615),
.B(n_445),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1711),
.B(n_449),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1543),
.A2(n_450),
.B(n_451),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1660),
.A2(n_1695),
.B1(n_1709),
.B2(n_1715),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1699),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1608),
.A2(n_452),
.B(n_453),
.C(n_454),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1701),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1707),
.B(n_456),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_SL g1957 ( 
.A1(n_1619),
.A2(n_458),
.B(n_459),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1520),
.A2(n_458),
.B(n_459),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1520),
.A2(n_460),
.B(n_461),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1520),
.A2(n_460),
.B(n_463),
.C(n_464),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1551),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1559),
.B(n_465),
.Y(n_1962)
);

AOI211x1_ASAP7_75t_L g1963 ( 
.A1(n_1573),
.A2(n_470),
.B(n_471),
.C(n_473),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1489),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1503),
.A2(n_476),
.B(n_477),
.C(n_478),
.Y(n_1965)
);

OA22x2_ASAP7_75t_L g1966 ( 
.A1(n_1673),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1597),
.B(n_481),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1597),
.B(n_481),
.Y(n_1968)
);

O2A1O1Ixp5_ASAP7_75t_L g1969 ( 
.A1(n_1531),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1551),
.B(n_482),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1623),
.A2(n_485),
.B(n_486),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1559),
.B(n_487),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1489),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1559),
.B(n_490),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1559),
.B(n_492),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1551),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1559),
.B(n_492),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1597),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_1978)
);

OAI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1503),
.A2(n_493),
.B(n_494),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1489),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1537),
.B(n_497),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1530),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1489),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1559),
.B(n_498),
.Y(n_1984)
);

OR2x6_ASAP7_75t_L g1985 ( 
.A(n_1607),
.B(n_498),
.Y(n_1985)
);

NOR2x1_ASAP7_75t_L g1986 ( 
.A(n_1607),
.B(n_499),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1489),
.Y(n_1987)
);

AO31x2_ASAP7_75t_L g1988 ( 
.A1(n_1680),
.A2(n_501),
.A3(n_502),
.B(n_503),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1559),
.B(n_501),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1559),
.B(n_503),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1537),
.B(n_504),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1597),
.B(n_506),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1597),
.A2(n_507),
.B1(n_508),
.B2(n_510),
.Y(n_1993)
);

AO31x2_ASAP7_75t_L g1994 ( 
.A1(n_1680),
.A2(n_510),
.A3(n_511),
.B(n_513),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1530),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1597),
.B(n_511),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1489),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1505),
.B(n_515),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1559),
.B(n_516),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1537),
.B(n_516),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1489),
.Y(n_2001)
);

NAND2x1_ASAP7_75t_L g2002 ( 
.A(n_1551),
.B(n_517),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1559),
.B(n_519),
.Y(n_2003)
);

INVx3_ASAP7_75t_SL g2004 ( 
.A(n_1604),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1604),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1604),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1559),
.B(n_520),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1559),
.B(n_521),
.Y(n_2008)
);

OAI21x1_ASAP7_75t_SL g2009 ( 
.A1(n_1623),
.A2(n_522),
.B(n_523),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1559),
.B(n_523),
.Y(n_2010)
);

AOI211x1_ASAP7_75t_L g2011 ( 
.A1(n_1573),
.A2(n_524),
.B(n_525),
.C(n_526),
.Y(n_2011)
);

AO31x2_ASAP7_75t_L g2012 ( 
.A1(n_1680),
.A2(n_527),
.A3(n_528),
.B(n_529),
.Y(n_2012)
);

NAND2x1_ASAP7_75t_L g2013 ( 
.A(n_1551),
.B(n_527),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1551),
.Y(n_2014)
);

A2O1A1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1503),
.A2(n_528),
.B(n_530),
.C(n_531),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1551),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1503),
.A2(n_531),
.B(n_532),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1530),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1559),
.B(n_533),
.Y(n_2019)
);

BUFx12f_ASAP7_75t_L g2020 ( 
.A(n_1572),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1597),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1710),
.B(n_535),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1551),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1505),
.B(n_1269),
.Y(n_2024)
);

OAI22x1_ASAP7_75t_L g2025 ( 
.A1(n_1673),
.A2(n_1096),
.B1(n_1063),
.B2(n_1283),
.Y(n_2025)
);

NAND3x1_ASAP7_75t_L g2026 ( 
.A(n_1674),
.B(n_1672),
.C(n_1616),
.Y(n_2026)
);

OAI21x1_ASAP7_75t_L g2027 ( 
.A1(n_1610),
.A2(n_1488),
.B(n_1511),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1559),
.B(n_1269),
.Y(n_2028)
);

OAI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1610),
.A2(n_1488),
.B(n_1511),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1597),
.B(n_1503),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1489),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1559),
.B(n_1269),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1551),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1559),
.B(n_1269),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1477),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1559),
.B(n_1269),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1530),
.Y(n_2037)
);

AOI211x1_ASAP7_75t_L g2038 ( 
.A1(n_1573),
.A2(n_1659),
.B(n_1668),
.C(n_1559),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1559),
.B(n_1269),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1551),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1597),
.A2(n_1625),
.B1(n_1630),
.B2(n_1627),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1537),
.B(n_1283),
.Y(n_2042)
);

INVx5_ASAP7_75t_L g2043 ( 
.A(n_1551),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1551),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2024),
.B(n_1809),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1825),
.A2(n_1985),
.B1(n_1734),
.B2(n_1916),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_2030),
.A2(n_2032),
.B(n_2028),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1730),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2024),
.B(n_2042),
.Y(n_2049)
);

NAND2x1p5_ASAP7_75t_L g2050 ( 
.A(n_2043),
.B(n_2014),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1737),
.A2(n_2029),
.B(n_2027),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1825),
.A2(n_1985),
.B1(n_1927),
.B2(n_1728),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_2043),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1725),
.B(n_1981),
.Y(n_2054)
);

OAI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_2034),
.A2(n_2039),
.B(n_2036),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1824),
.A2(n_1847),
.B1(n_1821),
.B2(n_1762),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1991),
.B(n_2000),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1820),
.Y(n_2058)
);

OAI21x1_ASAP7_75t_L g2059 ( 
.A1(n_1733),
.A2(n_1982),
.B(n_1742),
.Y(n_2059)
);

BUFx4_ASAP7_75t_R g2060 ( 
.A(n_1727),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1733),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1742),
.Y(n_2062)
);

AO31x2_ASAP7_75t_L g2063 ( 
.A1(n_1738),
.A2(n_1995),
.A3(n_2018),
.B(n_1982),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1747),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_2021),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2021),
.B(n_1721),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_2043),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1755),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2037),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1795),
.B(n_1848),
.Y(n_2070)
);

BUFx2_ASAP7_75t_R g2071 ( 
.A(n_1740),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_1817),
.A2(n_1882),
.B(n_1922),
.C(n_1726),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1964),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1781),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1740),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1973),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1779),
.B(n_1722),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1980),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_2004),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1821),
.B(n_1879),
.Y(n_2080)
);

BUFx4_ASAP7_75t_SL g2081 ( 
.A(n_1851),
.Y(n_2081)
);

INVxp67_ASAP7_75t_SL g2082 ( 
.A(n_1781),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_1757),
.A2(n_1752),
.B(n_1959),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1983),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1745),
.A2(n_1998),
.B1(n_1926),
.B2(n_1941),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2041),
.A2(n_1834),
.B1(n_1836),
.B2(n_1998),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2035),
.B(n_1743),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1848),
.B(n_1987),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_1789),
.B(n_1764),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1997),
.Y(n_2090)
);

INVx2_ASAP7_75t_SL g2091 ( 
.A(n_2004),
.Y(n_2091)
);

AO31x2_ASAP7_75t_L g2092 ( 
.A1(n_1827),
.A2(n_1960),
.A3(n_1858),
.B(n_1954),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2001),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_2031),
.B(n_1775),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1745),
.A2(n_1941),
.B1(n_1751),
.B2(n_1832),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1783),
.B(n_1884),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1832),
.A2(n_1986),
.B1(n_1871),
.B2(n_1966),
.Y(n_2097)
);

INVx2_ASAP7_75t_SL g2098 ( 
.A(n_2020),
.Y(n_2098)
);

INVxp67_ASAP7_75t_L g2099 ( 
.A(n_1834),
.Y(n_2099)
);

INVx4_ASAP7_75t_SL g2100 ( 
.A(n_1729),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1794),
.Y(n_2101)
);

INVx3_ASAP7_75t_L g2102 ( 
.A(n_1729),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1823),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_2005),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1752),
.A2(n_1758),
.B(n_1815),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1836),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_2005),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1735),
.A2(n_2022),
.B1(n_1905),
.B2(n_1883),
.Y(n_2108)
);

CKINVDCx20_ASAP7_75t_R g2109 ( 
.A(n_2006),
.Y(n_2109)
);

BUFx12f_ASAP7_75t_L g2110 ( 
.A(n_2006),
.Y(n_2110)
);

NOR2x1_ASAP7_75t_SL g2111 ( 
.A(n_1833),
.B(n_1961),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1720),
.A2(n_2026),
.B1(n_2022),
.B2(n_1735),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1754),
.Y(n_2113)
);

AOI22x1_ASAP7_75t_L g2114 ( 
.A1(n_1744),
.A2(n_1828),
.B1(n_1829),
.B2(n_1774),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1767),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1966),
.A2(n_1856),
.B1(n_1815),
.B2(n_1894),
.Y(n_2116)
);

INVx6_ASAP7_75t_L g2117 ( 
.A(n_1961),
.Y(n_2117)
);

AO21x2_ASAP7_75t_L g2118 ( 
.A1(n_1954),
.A2(n_2017),
.B(n_1979),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1867),
.B(n_1857),
.Y(n_2119)
);

INVx5_ASAP7_75t_L g2120 ( 
.A(n_1961),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1784),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_SL g2122 ( 
.A1(n_1816),
.A2(n_1873),
.B(n_2015),
.C(n_1965),
.Y(n_2122)
);

AOI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_1765),
.A2(n_2025),
.B1(n_2038),
.B2(n_1837),
.C(n_1801),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_1806),
.A2(n_1807),
.B1(n_1819),
.B2(n_1791),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1788),
.B(n_1841),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1784),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2023),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_2023),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_2020),
.Y(n_2129)
);

NAND3xp33_ASAP7_75t_L g2130 ( 
.A(n_1818),
.B(n_1895),
.C(n_1928),
.Y(n_2130)
);

AO21x1_ASAP7_75t_L g2131 ( 
.A1(n_1723),
.A2(n_1968),
.B(n_1967),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1906),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1891),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1768),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2040),
.B(n_1719),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_1869),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1804),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1770),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1886),
.B(n_1771),
.Y(n_2139)
);

CKINVDCx11_ASAP7_75t_R g2140 ( 
.A(n_1851),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1866),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_1952),
.A2(n_1962),
.B(n_1718),
.Y(n_2142)
);

A2O1A1Ixp33_ASAP7_75t_L g2143 ( 
.A1(n_1761),
.A2(n_1816),
.B(n_2015),
.C(n_1965),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1899),
.A2(n_1890),
.B(n_1889),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_2044),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1972),
.A2(n_1975),
.B(n_1974),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_1746),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1901),
.B(n_1830),
.Y(n_2148)
);

A2O1A1Ixp33_ASAP7_75t_L g2149 ( 
.A1(n_1773),
.A2(n_1939),
.B(n_1798),
.C(n_1739),
.Y(n_2149)
);

NAND2x1p5_ASAP7_75t_L g2150 ( 
.A(n_1776),
.B(n_1777),
.Y(n_2150)
);

INVx5_ASAP7_75t_L g2151 ( 
.A(n_1935),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_1776),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_1746),
.B(n_1888),
.Y(n_2153)
);

OA21x2_ASAP7_75t_L g2154 ( 
.A1(n_1960),
.A2(n_1800),
.B(n_1785),
.Y(n_2154)
);

CKINVDCx11_ASAP7_75t_R g2155 ( 
.A(n_1903),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_1777),
.B(n_1976),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1810),
.Y(n_2157)
);

INVx4_ASAP7_75t_L g2158 ( 
.A(n_2016),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_L g2159 ( 
.A1(n_1780),
.A2(n_1797),
.B1(n_1874),
.B2(n_1970),
.Y(n_2159)
);

OAI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1870),
.A2(n_1917),
.B1(n_1860),
.B2(n_1936),
.Y(n_2160)
);

AOI21x1_ASAP7_75t_L g2161 ( 
.A1(n_1977),
.A2(n_1989),
.B(n_1984),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_2044),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1932),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_1937),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_1937),
.Y(n_2165)
);

AOI222xp33_ASAP7_75t_L g2166 ( 
.A1(n_1831),
.A2(n_1787),
.B1(n_1915),
.B2(n_1934),
.C1(n_1852),
.C2(n_1803),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_SL g2167 ( 
.A1(n_1957),
.A2(n_1862),
.B(n_1859),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1838),
.B(n_1990),
.Y(n_2168)
);

OAI21x1_ASAP7_75t_L g2169 ( 
.A1(n_1778),
.A2(n_1796),
.B(n_1786),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1877),
.Y(n_2170)
);

AO21x2_ASAP7_75t_L g2171 ( 
.A1(n_1732),
.A2(n_1873),
.B(n_1999),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_2033),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_SL g2173 ( 
.A1(n_1749),
.A2(n_2009),
.B1(n_1907),
.B2(n_1897),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1826),
.A2(n_2007),
.B(n_2003),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2008),
.A2(n_2019),
.B(n_2010),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1854),
.B(n_1855),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1720),
.B(n_2026),
.Y(n_2177)
);

O2A1O1Ixp33_ASAP7_75t_SL g2178 ( 
.A1(n_1939),
.A2(n_1763),
.B(n_1911),
.C(n_1910),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1919),
.B(n_1865),
.Y(n_2179)
);

AOI221x1_ASAP7_75t_L g2180 ( 
.A1(n_1958),
.A2(n_1843),
.B1(n_1759),
.B2(n_1763),
.C(n_1881),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_R g2181 ( 
.A(n_1814),
.B(n_2033),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1853),
.B(n_1949),
.Y(n_2182)
);

NAND3xp33_ASAP7_75t_L g2183 ( 
.A(n_1756),
.B(n_1963),
.C(n_2011),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_1814),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1731),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1868),
.B(n_1896),
.Y(n_2186)
);

O2A1O1Ixp33_ASAP7_75t_SL g2187 ( 
.A1(n_1802),
.A2(n_1910),
.B(n_1911),
.C(n_1724),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1947),
.B(n_1853),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1887),
.A2(n_1930),
.B(n_1748),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1769),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_1904),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1909),
.B(n_1842),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1842),
.B(n_1840),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_1953),
.A2(n_1923),
.B1(n_1880),
.B2(n_1850),
.C(n_1844),
.Y(n_2194)
);

NOR2xp67_ASAP7_75t_SL g2195 ( 
.A(n_1971),
.B(n_1904),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1946),
.B(n_1933),
.Y(n_2196)
);

CKINVDCx6p67_ASAP7_75t_R g2197 ( 
.A(n_1723),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_1908),
.B(n_1950),
.Y(n_2198)
);

INVxp67_ASAP7_75t_SL g2199 ( 
.A(n_1970),
.Y(n_2199)
);

INVx1_ASAP7_75t_SL g2200 ( 
.A(n_1918),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1913),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1921),
.B(n_1799),
.Y(n_2202)
);

AO21x2_ASAP7_75t_L g2203 ( 
.A1(n_1925),
.A2(n_1912),
.B(n_1846),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1792),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_SL g2205 ( 
.A1(n_1717),
.A2(n_1978),
.B1(n_1993),
.B2(n_1902),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_2013),
.A2(n_2002),
.B(n_1766),
.Y(n_2206)
);

BUFx2_ASAP7_75t_R g2207 ( 
.A(n_1968),
.Y(n_2207)
);

O2A1O1Ixp33_ASAP7_75t_SL g2208 ( 
.A1(n_1802),
.A2(n_1996),
.B(n_1992),
.C(n_1940),
.Y(n_2208)
);

NAND2x1p5_ASAP7_75t_L g2209 ( 
.A(n_1929),
.B(n_1992),
.Y(n_2209)
);

O2A1O1Ixp5_ASAP7_75t_L g2210 ( 
.A1(n_1996),
.A2(n_1741),
.B(n_1969),
.C(n_1811),
.Y(n_2210)
);

OR2x6_ASAP7_75t_L g2211 ( 
.A(n_1924),
.B(n_1845),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1940),
.A2(n_1956),
.B1(n_1736),
.B2(n_1753),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_1805),
.A2(n_1864),
.B(n_1892),
.Y(n_2213)
);

AOI22x1_ASAP7_75t_L g2214 ( 
.A1(n_1812),
.A2(n_1750),
.B1(n_1931),
.B2(n_1920),
.Y(n_2214)
);

NAND2x1p5_ASAP7_75t_L g2215 ( 
.A(n_1929),
.B(n_1938),
.Y(n_2215)
);

OAI21x1_ASAP7_75t_L g2216 ( 
.A1(n_1872),
.A2(n_1876),
.B(n_1760),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1842),
.B(n_1942),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_1772),
.A2(n_1878),
.B(n_1943),
.Y(n_2218)
);

OAI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_1893),
.A2(n_1951),
.B(n_1948),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1808),
.A2(n_1944),
.B(n_1875),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_1918),
.B(n_1839),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1790),
.B(n_1863),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1835),
.B(n_1849),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_1914),
.A2(n_1955),
.B(n_1782),
.Y(n_2224)
);

A2O1A1Ixp33_ASAP7_75t_L g2225 ( 
.A1(n_1861),
.A2(n_1898),
.B(n_1885),
.C(n_1945),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1782),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_SL g2227 ( 
.A1(n_1813),
.A2(n_1945),
.B(n_1861),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1988),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_1813),
.B(n_1945),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1822),
.B(n_1945),
.Y(n_2230)
);

A2O1A1Ixp33_ASAP7_75t_SL g2231 ( 
.A1(n_1988),
.A2(n_2012),
.B(n_1994),
.C(n_1822),
.Y(n_2231)
);

AOI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_1813),
.A2(n_1793),
.B1(n_1898),
.B2(n_1861),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1988),
.Y(n_2233)
);

A2O1A1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_1885),
.A2(n_1898),
.B(n_1822),
.C(n_1900),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1900),
.Y(n_2235)
);

OAI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_1822),
.A2(n_1793),
.B(n_1885),
.Y(n_2236)
);

OAI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_1898),
.A2(n_2024),
.B(n_2028),
.Y(n_2237)
);

NAND2x1p5_ASAP7_75t_L g2238 ( 
.A(n_2043),
.B(n_1551),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1740),
.Y(n_2239)
);

OAI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2028),
.Y(n_2240)
);

OAI222xp33_ASAP7_75t_L g2241 ( 
.A1(n_1985),
.A2(n_1966),
.B1(n_1734),
.B2(n_1673),
.C1(n_1941),
.C2(n_1986),
.Y(n_2241)
);

AO32x2_ASAP7_75t_L g2242 ( 
.A1(n_1717),
.A2(n_1993),
.A3(n_1978),
.B1(n_1769),
.B2(n_1792),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2024),
.B(n_1809),
.Y(n_2243)
);

NOR2x1_ASAP7_75t_R g2244 ( 
.A(n_1745),
.B(n_1063),
.Y(n_2244)
);

INVx3_ASAP7_75t_SL g2245 ( 
.A(n_1740),
.Y(n_2245)
);

O2A1O1Ixp33_ASAP7_75t_L g2246 ( 
.A1(n_1965),
.A2(n_2015),
.B(n_1939),
.C(n_1816),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2024),
.A2(n_2041),
.B1(n_2021),
.B2(n_1985),
.Y(n_2247)
);

A2O1A1Ixp33_ASAP7_75t_L g2248 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2034),
.C(n_2028),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_1809),
.A2(n_1825),
.B1(n_1673),
.B2(n_1985),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_1809),
.A2(n_1825),
.B1(n_1673),
.B2(n_1985),
.Y(n_2250)
);

OAI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2028),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_1985),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1809),
.B(n_1574),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1730),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2024),
.A2(n_2041),
.B1(n_2021),
.B2(n_1985),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_2043),
.Y(n_2256)
);

BUFx3_ASAP7_75t_L g2257 ( 
.A(n_2043),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2028),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1730),
.Y(n_2259)
);

A2O1A1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2034),
.C(n_2028),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1730),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_1740),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2024),
.B(n_1269),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_1762),
.B(n_1283),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2024),
.B(n_1269),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_1985),
.Y(n_2266)
);

NOR2x1_ASAP7_75t_R g2267 ( 
.A(n_1745),
.B(n_1063),
.Y(n_2267)
);

AOI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_1809),
.A2(n_1825),
.B1(n_1673),
.B2(n_1985),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1730),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_1809),
.A2(n_1825),
.B1(n_1673),
.B2(n_1985),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1733),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2024),
.A2(n_2041),
.B1(n_2021),
.B2(n_1985),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_1762),
.B(n_1283),
.Y(n_2273)
);

AOI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2024),
.A2(n_1123),
.B1(n_1306),
.B2(n_1282),
.C(n_1179),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2021),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_2043),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_1729),
.Y(n_2277)
);

OAI211xp5_ASAP7_75t_SL g2278 ( 
.A1(n_1882),
.A2(n_1673),
.B(n_1579),
.C(n_1494),
.Y(n_2278)
);

NOR2x1_ASAP7_75t_SL g2279 ( 
.A(n_1985),
.B(n_2043),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2024),
.A2(n_2032),
.B(n_2028),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2024),
.A2(n_2041),
.B1(n_2021),
.B2(n_1985),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1730),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_1729),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2048),
.Y(n_2284)
);

INVx2_ASAP7_75t_SL g2285 ( 
.A(n_2058),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2064),
.Y(n_2286)
);

OR2x6_ASAP7_75t_L g2287 ( 
.A(n_2165),
.B(n_2252),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_SL g2288 ( 
.A1(n_2266),
.A2(n_2255),
.B1(n_2272),
.B2(n_2247),
.Y(n_2288)
);

BUFx3_ASAP7_75t_L g2289 ( 
.A(n_2238),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_2053),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2068),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_2053),
.Y(n_2292)
);

O2A1O1Ixp5_ASAP7_75t_L g2293 ( 
.A1(n_2236),
.A2(n_2105),
.B(n_2210),
.C(n_2234),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_2061),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2073),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2076),
.Y(n_2296)
);

INVx1_ASAP7_75t_SL g2297 ( 
.A(n_2070),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2078),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2084),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_2067),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2248),
.B(n_2260),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2090),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2279),
.B(n_2067),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2093),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2254),
.Y(n_2305)
);

INVx6_ASAP7_75t_L g2306 ( 
.A(n_2120),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2259),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2049),
.B(n_2045),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2256),
.B(n_2257),
.Y(n_2309)
);

HB1xp67_ASAP7_75t_L g2310 ( 
.A(n_2061),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2261),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2269),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2160),
.B(n_2281),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2062),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_2256),
.Y(n_2315)
);

NOR2x1_ASAP7_75t_R g2316 ( 
.A(n_2140),
.B(n_2129),
.Y(n_2316)
);

INVxp67_ASAP7_75t_L g2317 ( 
.A(n_2065),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2243),
.B(n_2263),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2282),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2101),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_2069),
.Y(n_2321)
);

BUFx2_ASAP7_75t_L g2322 ( 
.A(n_2181),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2112),
.A2(n_2046),
.B1(n_2250),
.B2(n_2249),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2238),
.Y(n_2324)
);

HB1xp67_ASAP7_75t_L g2325 ( 
.A(n_2069),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2248),
.B(n_2260),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2103),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2132),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2119),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_2257),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2276),
.B(n_2088),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2240),
.B(n_2251),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2094),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2271),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2265),
.B(n_2253),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2065),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2275),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2275),
.Y(n_2338)
);

OAI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2149),
.A2(n_2210),
.B(n_2143),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_2276),
.Y(n_2340)
);

OAI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2149),
.A2(n_2143),
.B(n_2130),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2074),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2066),
.B(n_2264),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2253),
.B(n_2054),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2278),
.B(n_2273),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2057),
.B(n_2087),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2249),
.A2(n_2250),
.B1(n_2270),
.B2(n_2268),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2081),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2059),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2082),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2082),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2070),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2188),
.Y(n_2353)
);

INVx5_ASAP7_75t_L g2354 ( 
.A(n_2120),
.Y(n_2354)
);

BUFx12f_ASAP7_75t_L g2355 ( 
.A(n_2129),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_SL g2356 ( 
.A(n_2160),
.B(n_2241),
.Y(n_2356)
);

INVx2_ASAP7_75t_SL g2357 ( 
.A(n_2081),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_2050),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2099),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2063),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_2164),
.Y(n_2361)
);

INVx4_ASAP7_75t_L g2362 ( 
.A(n_2245),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2120),
.B(n_2100),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2120),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2140),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2099),
.Y(n_2366)
);

BUFx2_ASAP7_75t_L g2367 ( 
.A(n_2050),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2106),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2106),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2096),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2047),
.A2(n_2055),
.B(n_2258),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2157),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_2100),
.B(n_2121),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2089),
.Y(n_2374)
);

OAI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2142),
.A2(n_2246),
.B(n_2183),
.Y(n_2375)
);

INVx6_ASAP7_75t_L g2376 ( 
.A(n_2104),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2111),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2139),
.Y(n_2378)
);

BUFx2_ASAP7_75t_SL g2379 ( 
.A(n_2191),
.Y(n_2379)
);

AO21x2_ASAP7_75t_L g2380 ( 
.A1(n_2227),
.A2(n_2167),
.B(n_2231),
.Y(n_2380)
);

AO31x2_ASAP7_75t_L g2381 ( 
.A1(n_2234),
.A2(n_2225),
.A3(n_2230),
.B(n_2228),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2182),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2100),
.B(n_2126),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2063),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2201),
.Y(n_2385)
);

AO31x2_ASAP7_75t_L g2386 ( 
.A1(n_2225),
.A2(n_2230),
.A3(n_2233),
.B(n_2228),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2063),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2060),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2245),
.Y(n_2389)
);

NAND2x1p5_ASAP7_75t_L g2390 ( 
.A(n_2151),
.B(n_2195),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2060),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2141),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_2151),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2170),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2056),
.B(n_2136),
.Y(n_2395)
);

OR2x6_ASAP7_75t_L g2396 ( 
.A(n_2075),
.B(n_2091),
.Y(n_2396)
);

AND2x6_ASAP7_75t_L g2397 ( 
.A(n_2177),
.B(n_2163),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2046),
.A2(n_2270),
.B1(n_2268),
.B2(n_2097),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2197),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2113),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2079),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2115),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2133),
.Y(n_2403)
);

OR2x6_ASAP7_75t_L g2404 ( 
.A(n_2158),
.B(n_2110),
.Y(n_2404)
);

INVx4_ASAP7_75t_L g2405 ( 
.A(n_2079),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_2151),
.B(n_2128),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2134),
.Y(n_2407)
);

OR2x6_ASAP7_75t_L g2408 ( 
.A(n_2158),
.B(n_2110),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2077),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2196),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2274),
.B(n_2123),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2196),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2127),
.Y(n_2413)
);

AOI222xp33_ASAP7_75t_L g2414 ( 
.A1(n_2241),
.A2(n_2280),
.B1(n_2267),
.B2(n_2244),
.C1(n_2097),
.C2(n_2085),
.Y(n_2414)
);

AOI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2278),
.A2(n_2080),
.B1(n_2095),
.B2(n_2072),
.Y(n_2415)
);

OA21x2_ASAP7_75t_L g2416 ( 
.A1(n_2169),
.A2(n_2232),
.B(n_2180),
.Y(n_2416)
);

AO21x1_ASAP7_75t_L g2417 ( 
.A1(n_2246),
.A2(n_2086),
.B(n_2229),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2125),
.B(n_2184),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2148),
.B(n_2200),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2095),
.B(n_2085),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2235),
.Y(n_2421)
);

CKINVDCx6p67_ASAP7_75t_R g2422 ( 
.A(n_2191),
.Y(n_2422)
);

AO21x1_ASAP7_75t_L g2423 ( 
.A1(n_2229),
.A2(n_2108),
.B(n_2212),
.Y(n_2423)
);

AOI22xp33_ASAP7_75t_SL g2424 ( 
.A1(n_2114),
.A2(n_2199),
.B1(n_2223),
.B2(n_2118),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2196),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_SL g2426 ( 
.A1(n_2199),
.A2(n_2223),
.B1(n_2118),
.B2(n_2204),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2137),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2185),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2198),
.B(n_2186),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2190),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2207),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2052),
.A2(n_2116),
.B1(n_2205),
.B2(n_2124),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2080),
.B(n_2116),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2237),
.B(n_2124),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_2239),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2153),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2229),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2152),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2138),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2104),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2192),
.B(n_2174),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2138),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2145),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2162),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2131),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2051),
.Y(n_2446)
);

OR2x6_ASAP7_75t_L g2447 ( 
.A(n_2211),
.B(n_2098),
.Y(n_2447)
);

BUFx2_ASAP7_75t_L g2448 ( 
.A(n_2239),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2137),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2226),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_2343),
.B(n_2419),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2308),
.B(n_2217),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2294),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2346),
.B(n_2172),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2379),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2335),
.B(n_2329),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2354),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2344),
.B(n_2172),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2318),
.B(n_2166),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2370),
.B(n_2176),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2400),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2414),
.A2(n_2205),
.B1(n_2222),
.B2(n_2159),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2402),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2403),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2410),
.B(n_2221),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2407),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2284),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_2382),
.B(n_2193),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2286),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2354),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2291),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2354),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2354),
.Y(n_2473)
);

INVx8_ASAP7_75t_L g2474 ( 
.A(n_2404),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2295),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2296),
.Y(n_2476)
);

BUFx2_ASAP7_75t_SL g2477 ( 
.A(n_2362),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2378),
.B(n_2150),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2414),
.A2(n_2168),
.B1(n_2194),
.B2(n_2179),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2412),
.B(n_2221),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2298),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2309),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2299),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2425),
.B(n_2437),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2436),
.B(n_2156),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2374),
.B(n_2202),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2418),
.B(n_2135),
.Y(n_2487)
);

AND2x4_ASAP7_75t_L g2488 ( 
.A(n_2392),
.B(n_2221),
.Y(n_2488)
);

BUFx2_ASAP7_75t_L g2489 ( 
.A(n_2303),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2302),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2411),
.B(n_2146),
.Y(n_2491)
);

OR2x2_ASAP7_75t_L g2492 ( 
.A(n_2317),
.B(n_2262),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2331),
.B(n_2147),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2304),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2305),
.Y(n_2495)
);

INVxp67_ASAP7_75t_SL g2496 ( 
.A(n_2294),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2307),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2311),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2312),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2319),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2320),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2327),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_2415),
.B(n_2071),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2310),
.B(n_2154),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2310),
.B(n_2154),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2314),
.B(n_2154),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2314),
.B(n_2203),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2321),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2328),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2359),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2366),
.Y(n_2511)
);

OR2x2_ASAP7_75t_L g2512 ( 
.A(n_2336),
.B(n_2262),
.Y(n_2512)
);

INVxp67_ASAP7_75t_L g2513 ( 
.A(n_2321),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2368),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2363),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2325),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2325),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2429),
.B(n_2242),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2369),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2334),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2334),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2340),
.B(n_2242),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2420),
.B(n_2242),
.Y(n_2523)
);

HB1xp67_ASAP7_75t_L g2524 ( 
.A(n_2413),
.Y(n_2524)
);

NOR2x1_ASAP7_75t_L g2525 ( 
.A(n_2362),
.B(n_2211),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2337),
.B(n_2107),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2350),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2351),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2338),
.B(n_2107),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2309),
.B(n_2433),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2345),
.B(n_2242),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2342),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2353),
.B(n_2175),
.Y(n_2533)
);

BUFx3_ASAP7_75t_L g2534 ( 
.A(n_2358),
.Y(n_2534)
);

INVx2_ASAP7_75t_SL g2535 ( 
.A(n_2363),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2345),
.B(n_2155),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2428),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2394),
.B(n_2211),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2347),
.B(n_2173),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2430),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2285),
.B(n_2173),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2413),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2372),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2398),
.B(n_2283),
.Y(n_2544)
);

INVxp67_ASAP7_75t_R g2545 ( 
.A(n_2422),
.Y(n_2545)
);

OR2x2_ASAP7_75t_L g2546 ( 
.A(n_2398),
.B(n_2277),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2409),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2367),
.B(n_2219),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2446),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2385),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2434),
.B(n_2171),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2322),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2434),
.B(n_2171),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2438),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2332),
.B(n_2144),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2332),
.B(n_2122),
.Y(n_2556)
);

AO31x2_ASAP7_75t_L g2557 ( 
.A1(n_2417),
.A2(n_2423),
.A3(n_2371),
.B(n_2301),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2431),
.B(n_2102),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2355),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_2349),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2358),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2349),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2288),
.A2(n_2209),
.B(n_2215),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2323),
.B(n_2215),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2432),
.B(n_2122),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2333),
.B(n_2155),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2306),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2421),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2323),
.B(n_2092),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2395),
.B(n_2092),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2432),
.B(n_2178),
.Y(n_2571)
);

BUFx2_ASAP7_75t_SL g2572 ( 
.A(n_2348),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2290),
.B(n_2161),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_R g2574 ( 
.A(n_2365),
.B(n_2109),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2290),
.B(n_2216),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2375),
.B(n_2178),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2300),
.B(n_2117),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2297),
.B(n_2092),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2300),
.B(n_2117),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2292),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2375),
.B(n_2208),
.Y(n_2581)
);

INVxp67_ASAP7_75t_L g2582 ( 
.A(n_2356),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2339),
.B(n_2083),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2339),
.B(n_2083),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2301),
.B(n_2208),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2315),
.B(n_2117),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_L g2587 ( 
.A(n_2503),
.B(n_2399),
.C(n_2389),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2549),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2518),
.B(n_2288),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2547),
.B(n_2326),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2461),
.Y(n_2591)
);

OR2x2_ASAP7_75t_L g2592 ( 
.A(n_2452),
.B(n_2297),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2451),
.B(n_2456),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2468),
.B(n_2441),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2463),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2523),
.B(n_2551),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2462),
.A2(n_2356),
.B1(n_2313),
.B2(n_2388),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2530),
.B(n_2487),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2538),
.B(n_2380),
.Y(n_2599)
);

AOI222xp33_ASAP7_75t_L g2600 ( 
.A1(n_2462),
.A2(n_2479),
.B1(n_2539),
.B2(n_2459),
.C1(n_2491),
.C2(n_2503),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2454),
.B(n_2361),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2551),
.B(n_2381),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2464),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2466),
.Y(n_2604)
);

NAND3xp33_ASAP7_75t_L g2605 ( 
.A(n_2479),
.B(n_2341),
.C(n_2445),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2531),
.B(n_2326),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2553),
.B(n_2381),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2532),
.B(n_2533),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2460),
.B(n_2447),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2553),
.B(n_2381),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2583),
.B(n_2381),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2453),
.B(n_2441),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2467),
.Y(n_2613)
);

NAND2x1p5_ASAP7_75t_L g2614 ( 
.A(n_2470),
.B(n_2472),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2469),
.Y(n_2615)
);

BUFx2_ASAP7_75t_L g2616 ( 
.A(n_2474),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2471),
.B(n_2313),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2583),
.B(n_2386),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2584),
.B(n_2386),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2584),
.B(n_2386),
.Y(n_2620)
);

BUFx2_ASAP7_75t_L g2621 ( 
.A(n_2474),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2453),
.B(n_2361),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2475),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2522),
.B(n_2386),
.Y(n_2624)
);

AND2x4_ASAP7_75t_L g2625 ( 
.A(n_2538),
.B(n_2380),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2538),
.B(n_2397),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2474),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2476),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2477),
.A2(n_2391),
.B1(n_2447),
.B2(n_2390),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2508),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2481),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2504),
.B(n_2384),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2483),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2504),
.B(n_2384),
.Y(n_2634)
);

AND2x4_ASAP7_75t_L g2635 ( 
.A(n_2488),
.B(n_2397),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2490),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2488),
.B(n_2397),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2458),
.B(n_2486),
.Y(n_2638)
);

HB1xp67_ASAP7_75t_L g2639 ( 
.A(n_2496),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2494),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2495),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2497),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2498),
.Y(n_2643)
);

INVx2_ASAP7_75t_SL g2644 ( 
.A(n_2482),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2499),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2500),
.B(n_2371),
.Y(n_2646)
);

AND2x4_ASAP7_75t_SL g2647 ( 
.A(n_2515),
.B(n_2404),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2501),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2502),
.B(n_2341),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2505),
.B(n_2450),
.Y(n_2650)
);

BUFx2_ASAP7_75t_L g2651 ( 
.A(n_2489),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2509),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2525),
.B(n_2426),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2543),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2541),
.B(n_2447),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2493),
.B(n_2352),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2465),
.B(n_2397),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2510),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2511),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2514),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2519),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2537),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_2496),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2540),
.Y(n_2664)
);

INVx1_ASAP7_75t_SL g2665 ( 
.A(n_2574),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2527),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2528),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2568),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2554),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2506),
.B(n_2360),
.Y(n_2670)
);

AND2x2_ASAP7_75t_SL g2671 ( 
.A(n_2568),
.B(n_2516),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2550),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2507),
.B(n_2516),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2524),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2507),
.B(n_2387),
.Y(n_2675)
);

OR2x2_ASAP7_75t_L g2676 ( 
.A(n_2513),
.B(n_2287),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2524),
.Y(n_2677)
);

NOR2xp67_ASAP7_75t_L g2678 ( 
.A(n_2457),
.B(n_2357),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2517),
.B(n_2426),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2589),
.B(n_2571),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2611),
.B(n_2618),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2611),
.B(n_2480),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2639),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2646),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2618),
.B(n_2480),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2596),
.B(n_2570),
.Y(n_2686)
);

NAND2x1_ASAP7_75t_L g2687 ( 
.A(n_2635),
.B(n_2520),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2619),
.B(n_2480),
.Y(n_2688)
);

AND2x4_ASAP7_75t_L g2689 ( 
.A(n_2599),
.B(n_2575),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2599),
.B(n_2484),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2588),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2596),
.B(n_2569),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2619),
.B(n_2578),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2606),
.B(n_2565),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2599),
.B(n_2484),
.Y(n_2695)
);

NOR2x1_ASAP7_75t_L g2696 ( 
.A(n_2678),
.B(n_2572),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2620),
.B(n_2520),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2620),
.B(n_2521),
.Y(n_2698)
);

NAND2xp33_ASAP7_75t_SL g2699 ( 
.A(n_2616),
.B(n_2574),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2602),
.B(n_2521),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2602),
.B(n_2484),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2672),
.Y(n_2702)
);

AND2x2_ASAP7_75t_SL g2703 ( 
.A(n_2635),
.B(n_2637),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2617),
.B(n_2594),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2607),
.B(n_2548),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2607),
.B(n_2416),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2612),
.B(n_2513),
.Y(n_2707)
);

NOR2x1_ASAP7_75t_L g2708 ( 
.A(n_2665),
.B(n_2470),
.Y(n_2708)
);

HB1xp67_ASAP7_75t_L g2709 ( 
.A(n_2639),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2591),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2610),
.B(n_2416),
.Y(n_2711)
);

INVxp67_ASAP7_75t_L g2712 ( 
.A(n_2651),
.Y(n_2712)
);

BUFx2_ASAP7_75t_L g2713 ( 
.A(n_2668),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2595),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2603),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2604),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2610),
.B(n_2624),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2624),
.B(n_2560),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2613),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2625),
.B(n_2573),
.Y(n_2720)
);

NOR2x1_ASAP7_75t_L g2721 ( 
.A(n_2621),
.B(n_2472),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2625),
.B(n_2560),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2615),
.Y(n_2723)
);

OR2x2_ASAP7_75t_L g2724 ( 
.A(n_2673),
.B(n_2542),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2623),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2628),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2670),
.B(n_2675),
.Y(n_2727)
);

NAND2x1p5_ASAP7_75t_L g2728 ( 
.A(n_2671),
.B(n_2473),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2670),
.B(n_2562),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2631),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2673),
.B(n_2542),
.Y(n_2731)
);

INVx3_ASAP7_75t_L g2732 ( 
.A(n_2728),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2702),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2717),
.B(n_2681),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2702),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2690),
.B(n_2657),
.Y(n_2736)
);

NOR2xp67_ASAP7_75t_L g2737 ( 
.A(n_2712),
.B(n_2663),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2710),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2710),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2714),
.Y(n_2740)
);

OR2x2_ASAP7_75t_L g2741 ( 
.A(n_2692),
.B(n_2593),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2727),
.B(n_2632),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2692),
.B(n_2663),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2727),
.B(n_2632),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2696),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2713),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2713),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2681),
.B(n_2634),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2714),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2717),
.B(n_2598),
.Y(n_2750)
);

OR2x2_ASAP7_75t_L g2751 ( 
.A(n_2724),
.B(n_2630),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2724),
.B(n_2630),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2715),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2715),
.Y(n_2754)
);

INVx3_ASAP7_75t_L g2755 ( 
.A(n_2728),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2716),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2716),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2719),
.Y(n_2758)
);

INVxp33_ASAP7_75t_L g2759 ( 
.A(n_2708),
.Y(n_2759)
);

INVxp33_ASAP7_75t_L g2760 ( 
.A(n_2728),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2680),
.B(n_2674),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_SL g2762 ( 
.A(n_2721),
.B(n_2627),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2719),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2706),
.B(n_2634),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2723),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2694),
.B(n_2605),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2731),
.B(n_2592),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2731),
.B(n_2622),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2684),
.B(n_2718),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2706),
.B(n_2679),
.Y(n_2770)
);

OR2x2_ASAP7_75t_L g2771 ( 
.A(n_2686),
.B(n_2677),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2684),
.B(n_2600),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2704),
.B(n_2650),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2718),
.B(n_2650),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2699),
.B(n_2671),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2685),
.B(n_2688),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2690),
.B(n_2657),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2691),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2683),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2691),
.Y(n_2780)
);

AOI32xp33_ASAP7_75t_L g2781 ( 
.A1(n_2701),
.A2(n_2587),
.A3(n_2455),
.B1(n_2647),
.B2(n_2552),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2711),
.B(n_2679),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2685),
.B(n_2601),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2743),
.Y(n_2784)
);

OAI21xp33_ASAP7_75t_L g2785 ( 
.A1(n_2772),
.A2(n_2597),
.B(n_2705),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2732),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2751),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2752),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2766),
.A2(n_2597),
.B1(n_2609),
.B2(n_2536),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2733),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2735),
.Y(n_2791)
);

OAI32xp33_ASAP7_75t_L g2792 ( 
.A1(n_2759),
.A2(n_2614),
.A3(n_2709),
.B1(n_2707),
.B2(n_2473),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2745),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2746),
.Y(n_2794)
);

AOI32xp33_ASAP7_75t_L g2795 ( 
.A1(n_2759),
.A2(n_2647),
.A3(n_2701),
.B1(n_2688),
.B2(n_2682),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2770),
.B(n_2711),
.Y(n_2796)
);

NAND2x1p5_ASAP7_75t_L g2797 ( 
.A(n_2732),
.B(n_2687),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2746),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2766),
.B(n_2693),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2738),
.Y(n_2800)
);

AOI21xp33_ASAP7_75t_SL g2801 ( 
.A1(n_2775),
.A2(n_2703),
.B(n_2629),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2747),
.Y(n_2802)
);

AOI32xp33_ASAP7_75t_L g2803 ( 
.A1(n_2762),
.A2(n_2775),
.A3(n_2760),
.B1(n_2750),
.B2(n_2748),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2764),
.B(n_2690),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2770),
.B(n_2693),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2739),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2782),
.B(n_2729),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2782),
.B(n_2729),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2747),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2737),
.A2(n_2536),
.B1(n_2655),
.B2(n_2609),
.Y(n_2810)
);

AOI22xp33_ASAP7_75t_L g2811 ( 
.A1(n_2741),
.A2(n_2655),
.B1(n_2582),
.B2(n_2656),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2761),
.B(n_2723),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2742),
.B(n_2700),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2748),
.B(n_2682),
.Y(n_2814)
);

OAI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2779),
.A2(n_2653),
.B(n_2563),
.Y(n_2815)
);

INVxp67_ASAP7_75t_L g2816 ( 
.A(n_2768),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2764),
.B(n_2697),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2740),
.Y(n_2818)
);

OAI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2760),
.A2(n_2653),
.B(n_2582),
.Y(n_2819)
);

O2A1O1Ixp33_ASAP7_75t_L g2820 ( 
.A1(n_2769),
.A2(n_2440),
.B(n_2555),
.C(n_2529),
.Y(n_2820)
);

AOI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2736),
.A2(n_2703),
.B1(n_2720),
.B2(n_2689),
.Y(n_2821)
);

INVxp67_ASAP7_75t_L g2822 ( 
.A(n_2767),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2776),
.B(n_2695),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2734),
.B(n_2725),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2774),
.B(n_2707),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2778),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2749),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2778),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2742),
.B(n_2697),
.Y(n_2829)
);

OAI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2732),
.A2(n_2614),
.B(n_2457),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2753),
.Y(n_2831)
);

NAND3xp33_ASAP7_75t_L g2832 ( 
.A(n_2803),
.B(n_2781),
.C(n_2365),
.Y(n_2832)
);

AOI21xp33_ASAP7_75t_L g2833 ( 
.A1(n_2793),
.A2(n_2396),
.B(n_2492),
.Y(n_2833)
);

O2A1O1Ixp33_ASAP7_75t_SL g2834 ( 
.A1(n_2801),
.A2(n_2687),
.B(n_2755),
.C(n_2535),
.Y(n_2834)
);

OAI21xp5_ASAP7_75t_SL g2835 ( 
.A1(n_2815),
.A2(n_2795),
.B(n_2797),
.Y(n_2835)
);

OAI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2821),
.A2(n_2755),
.B1(n_2644),
.B2(n_2773),
.Y(n_2836)
);

OAI32xp33_ASAP7_75t_L g2837 ( 
.A1(n_2797),
.A2(n_2755),
.A3(n_2744),
.B1(n_2771),
.B2(n_2783),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2790),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2785),
.B(n_2744),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_SL g2840 ( 
.A(n_2786),
.B(n_2820),
.Y(n_2840)
);

CKINVDCx20_ASAP7_75t_R g2841 ( 
.A(n_2810),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2786),
.Y(n_2842)
);

AOI211xp5_ASAP7_75t_SL g2843 ( 
.A1(n_2786),
.A2(n_2576),
.B(n_2581),
.C(n_2564),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2792),
.A2(n_2830),
.B(n_2819),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2799),
.B(n_2754),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2812),
.B(n_2756),
.Y(n_2846)
);

OAI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2811),
.A2(n_2777),
.B1(n_2736),
.B2(n_2695),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2812),
.B(n_2757),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2791),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2800),
.Y(n_2850)
);

NAND2x1p5_ASAP7_75t_L g2851 ( 
.A(n_2794),
.B(n_2534),
.Y(n_2851)
);

OR2x2_ASAP7_75t_L g2852 ( 
.A(n_2825),
.B(n_2698),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2806),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2789),
.A2(n_2777),
.B1(n_2736),
.B2(n_2720),
.Y(n_2854)
);

AOI221xp5_ASAP7_75t_L g2855 ( 
.A1(n_2824),
.A2(n_2822),
.B1(n_2816),
.B2(n_2789),
.C(n_2784),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2824),
.B(n_2758),
.Y(n_2856)
);

O2A1O1Ixp33_ASAP7_75t_L g2857 ( 
.A1(n_2794),
.A2(n_2526),
.B(n_2396),
.C(n_2512),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2807),
.B(n_2698),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2805),
.B(n_2763),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2818),
.Y(n_2860)
);

AOI211xp5_ASAP7_75t_L g2861 ( 
.A1(n_2832),
.A2(n_2545),
.B(n_2316),
.C(n_2559),
.Y(n_2861)
);

OAI21xp5_ASAP7_75t_L g2862 ( 
.A1(n_2832),
.A2(n_2802),
.B(n_2798),
.Y(n_2862)
);

AOI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2841),
.A2(n_2835),
.B1(n_2855),
.B2(n_2847),
.Y(n_2863)
);

OAI21xp33_ASAP7_75t_L g2864 ( 
.A1(n_2854),
.A2(n_2811),
.B(n_2788),
.Y(n_2864)
);

NOR2x1_ASAP7_75t_L g2865 ( 
.A(n_2840),
.B(n_2404),
.Y(n_2865)
);

OAI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2839),
.A2(n_2814),
.B1(n_2808),
.B2(n_2805),
.Y(n_2866)
);

AOI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2834),
.A2(n_2802),
.B(n_2798),
.Y(n_2867)
);

OAI21xp33_ASAP7_75t_L g2868 ( 
.A1(n_2837),
.A2(n_2787),
.B(n_2809),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2846),
.B(n_2796),
.Y(n_2869)
);

AOI222xp33_ASAP7_75t_L g2870 ( 
.A1(n_2836),
.A2(n_2809),
.B1(n_2796),
.B2(n_2827),
.C1(n_2831),
.C2(n_2669),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2859),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2851),
.B(n_2804),
.Y(n_2872)
);

AOI211xp5_ASAP7_75t_SL g2873 ( 
.A1(n_2844),
.A2(n_2566),
.B(n_2109),
.C(n_2558),
.Y(n_2873)
);

NOR4xp25_ASAP7_75t_L g2874 ( 
.A(n_2833),
.B(n_2814),
.C(n_2633),
.D(n_2640),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2848),
.B(n_2829),
.Y(n_2875)
);

OAI221xp5_ASAP7_75t_L g2876 ( 
.A1(n_2843),
.A2(n_2765),
.B1(n_2813),
.B2(n_2828),
.C(n_2826),
.Y(n_2876)
);

NOR2x1_ASAP7_75t_L g2877 ( 
.A(n_2842),
.B(n_2408),
.Y(n_2877)
);

OAI221xp5_ASAP7_75t_L g2878 ( 
.A1(n_2857),
.A2(n_2828),
.B1(n_2826),
.B2(n_2376),
.C(n_2424),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2845),
.A2(n_2777),
.B1(n_2720),
.B2(n_2817),
.Y(n_2879)
);

AOI221xp5_ASAP7_75t_L g2880 ( 
.A1(n_2856),
.A2(n_2849),
.B1(n_2853),
.B2(n_2850),
.C(n_2838),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2860),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2852),
.B(n_2829),
.Y(n_2882)
);

OAI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2842),
.A2(n_2817),
.B(n_2424),
.Y(n_2883)
);

OAI21xp33_ASAP7_75t_SL g2884 ( 
.A1(n_2858),
.A2(n_2823),
.B(n_2644),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_SL g2885 ( 
.A1(n_2835),
.A2(n_2390),
.B(n_2401),
.Y(n_2885)
);

AOI21xp33_ASAP7_75t_SL g2886 ( 
.A1(n_2832),
.A2(n_2559),
.B(n_2408),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2859),
.Y(n_2887)
);

NAND3xp33_ASAP7_75t_SL g2888 ( 
.A(n_2835),
.B(n_2435),
.C(n_2448),
.Y(n_2888)
);

AOI221xp5_ASAP7_75t_L g2889 ( 
.A1(n_2837),
.A2(n_2730),
.B1(n_2726),
.B2(n_2725),
.C(n_2659),
.Y(n_2889)
);

OAI21xp5_ASAP7_75t_SL g2890 ( 
.A1(n_2835),
.A2(n_2626),
.B(n_2695),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2881),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2871),
.B(n_2726),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2887),
.B(n_2730),
.Y(n_2893)
);

OR2x2_ASAP7_75t_L g2894 ( 
.A(n_2866),
.B(n_2780),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2875),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2888),
.A2(n_2408),
.B(n_2396),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2863),
.B(n_2638),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2880),
.B(n_2658),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2874),
.B(n_2660),
.Y(n_2899)
);

HB1xp67_ASAP7_75t_L g2900 ( 
.A(n_2862),
.Y(n_2900)
);

NOR3x1_ASAP7_75t_L g2901 ( 
.A(n_2885),
.B(n_2535),
.C(n_2515),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2882),
.B(n_2661),
.Y(n_2902)
);

NAND3xp33_ASAP7_75t_L g2903 ( 
.A(n_2873),
.B(n_2435),
.C(n_2405),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2864),
.B(n_2636),
.Y(n_2904)
);

OAI211xp5_ASAP7_75t_L g2905 ( 
.A1(n_2886),
.A2(n_2405),
.B(n_2561),
.C(n_2534),
.Y(n_2905)
);

INVx2_ASAP7_75t_SL g2906 ( 
.A(n_2877),
.Y(n_2906)
);

NOR3xp33_ASAP7_75t_L g2907 ( 
.A(n_2862),
.B(n_2330),
.C(n_2315),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2869),
.B(n_2780),
.Y(n_2908)
);

NAND3xp33_ASAP7_75t_L g2909 ( 
.A(n_2873),
.B(n_2214),
.C(n_2641),
.Y(n_2909)
);

NAND3xp33_ASAP7_75t_L g2910 ( 
.A(n_2865),
.B(n_2643),
.C(n_2642),
.Y(n_2910)
);

NAND3xp33_ASAP7_75t_L g2911 ( 
.A(n_2890),
.B(n_2648),
.C(n_2645),
.Y(n_2911)
);

HB1xp67_ASAP7_75t_L g2912 ( 
.A(n_2884),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2895),
.B(n_2872),
.Y(n_2913)
);

NOR3xp33_ASAP7_75t_L g2914 ( 
.A(n_2912),
.B(n_2861),
.C(n_2878),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2892),
.Y(n_2915)
);

NOR2x1_ASAP7_75t_L g2916 ( 
.A(n_2903),
.B(n_2876),
.Y(n_2916)
);

NOR2x1p5_ASAP7_75t_L g2917 ( 
.A(n_2903),
.B(n_2870),
.Y(n_2917)
);

AOI211x1_ASAP7_75t_SL g2918 ( 
.A1(n_2897),
.A2(n_2883),
.B(n_2867),
.C(n_2868),
.Y(n_2918)
);

NAND4xp75_ASAP7_75t_L g2919 ( 
.A(n_2901),
.B(n_2896),
.C(n_2906),
.D(n_2889),
.Y(n_2919)
);

NOR3xp33_ASAP7_75t_L g2920 ( 
.A(n_2905),
.B(n_2879),
.C(n_2330),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2891),
.B(n_2652),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_SL g2922 ( 
.A1(n_2910),
.A2(n_2376),
.B1(n_2561),
.B2(n_2306),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2893),
.Y(n_2923)
);

NOR3xp33_ASAP7_75t_SL g2924 ( 
.A(n_2909),
.B(n_2376),
.C(n_2608),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_L g2925 ( 
.A(n_2900),
.B(n_2449),
.C(n_2427),
.Y(n_2925)
);

NOR2x1_ASAP7_75t_L g2926 ( 
.A(n_2899),
.B(n_2911),
.Y(n_2926)
);

NAND3xp33_ASAP7_75t_L g2927 ( 
.A(n_2904),
.B(n_2189),
.C(n_2439),
.Y(n_2927)
);

NOR3xp33_ASAP7_75t_L g2928 ( 
.A(n_2898),
.B(n_2449),
.C(n_2427),
.Y(n_2928)
);

NOR3xp33_ASAP7_75t_SL g2929 ( 
.A(n_2902),
.B(n_2649),
.C(n_2590),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2894),
.B(n_2364),
.Y(n_2930)
);

XOR2xp5_ASAP7_75t_L g2931 ( 
.A(n_2918),
.B(n_2908),
.Y(n_2931)
);

NOR3xp33_ASAP7_75t_L g2932 ( 
.A(n_2919),
.B(n_2907),
.C(n_2377),
.Y(n_2932)
);

NOR2x1_ASAP7_75t_L g2933 ( 
.A(n_2916),
.B(n_2393),
.Y(n_2933)
);

NAND4xp75_ASAP7_75t_L g2934 ( 
.A(n_2926),
.B(n_2567),
.C(n_2579),
.D(n_2577),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2913),
.B(n_2654),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2915),
.B(n_2662),
.Y(n_2936)
);

NAND4xp75_ASAP7_75t_L g2937 ( 
.A(n_2924),
.B(n_2567),
.C(n_2586),
.D(n_2220),
.Y(n_2937)
);

NAND3xp33_ASAP7_75t_L g2938 ( 
.A(n_2914),
.B(n_2443),
.C(n_2442),
.Y(n_2938)
);

AND2x4_ASAP7_75t_L g2939 ( 
.A(n_2928),
.B(n_2664),
.Y(n_2939)
);

XOR2x1_ASAP7_75t_L g2940 ( 
.A(n_2917),
.B(n_2373),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2922),
.A2(n_2585),
.B(n_2556),
.Y(n_2941)
);

OAI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2925),
.A2(n_2293),
.B(n_2224),
.Y(n_2942)
);

OR2x2_ASAP7_75t_L g2943 ( 
.A(n_2923),
.B(n_2557),
.Y(n_2943)
);

NOR2x1_ASAP7_75t_L g2944 ( 
.A(n_2921),
.B(n_2393),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2933),
.B(n_2929),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2931),
.B(n_2921),
.Y(n_2946)
);

NOR2xp67_ASAP7_75t_L g2947 ( 
.A(n_2938),
.B(n_2930),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2932),
.B(n_2920),
.Y(n_2948)
);

NOR2x1_ASAP7_75t_L g2949 ( 
.A(n_2934),
.B(n_2927),
.Y(n_2949)
);

NOR2x1_ASAP7_75t_L g2950 ( 
.A(n_2937),
.B(n_2289),
.Y(n_2950)
);

NOR3xp33_ASAP7_75t_L g2951 ( 
.A(n_2944),
.B(n_2942),
.C(n_2941),
.Y(n_2951)
);

OR2x2_ASAP7_75t_L g2952 ( 
.A(n_2935),
.B(n_2557),
.Y(n_2952)
);

OAI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2943),
.A2(n_2206),
.B(n_2213),
.Y(n_2953)
);

NOR2xp67_ASAP7_75t_SL g2954 ( 
.A(n_2940),
.B(n_2306),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2939),
.Y(n_2955)
);

AOI222xp33_ASAP7_75t_L g2956 ( 
.A1(n_2946),
.A2(n_2936),
.B1(n_2666),
.B2(n_2667),
.C1(n_2485),
.C2(n_2478),
.Y(n_2956)
);

XNOR2x2_ASAP7_75t_L g2957 ( 
.A(n_2950),
.B(n_2218),
.Y(n_2957)
);

XNOR2xp5_ASAP7_75t_L g2958 ( 
.A(n_2948),
.B(n_2373),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2955),
.B(n_2945),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2947),
.B(n_2722),
.Y(n_2960)
);

OAI221xp5_ASAP7_75t_SL g2961 ( 
.A1(n_2951),
.A2(n_2287),
.B1(n_2544),
.B2(n_2546),
.C(n_2676),
.Y(n_2961)
);

OAI22xp5_ASAP7_75t_SL g2962 ( 
.A1(n_2950),
.A2(n_2406),
.B1(n_2364),
.B2(n_2324),
.Y(n_2962)
);

XNOR2xp5_ASAP7_75t_L g2963 ( 
.A(n_2949),
.B(n_2383),
.Y(n_2963)
);

AND2x4_ASAP7_75t_L g2964 ( 
.A(n_2952),
.B(n_2689),
.Y(n_2964)
);

OAI22x1_ASAP7_75t_L g2965 ( 
.A1(n_2959),
.A2(n_2954),
.B1(n_2953),
.B2(n_2383),
.Y(n_2965)
);

AOI22x1_ASAP7_75t_L g2966 ( 
.A1(n_2963),
.A2(n_2406),
.B1(n_2364),
.B2(n_2580),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2960),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2956),
.Y(n_2968)
);

BUFx2_ASAP7_75t_L g2969 ( 
.A(n_2957),
.Y(n_2969)
);

OAI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2967),
.A2(n_2958),
.B(n_2961),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2970),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2971),
.B(n_2968),
.Y(n_2972)
);

AO21x2_ASAP7_75t_L g2973 ( 
.A1(n_2972),
.A2(n_2969),
.B(n_2964),
.Y(n_2973)
);

AOI221xp5_ASAP7_75t_L g2974 ( 
.A1(n_2973),
.A2(n_2965),
.B1(n_2962),
.B2(n_2966),
.C(n_2444),
.Y(n_2974)
);

AOI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2974),
.A2(n_2965),
.B(n_2187),
.Y(n_2975)
);


endmodule