module fake_jpeg_6416_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_27),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.C(n_20),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_26),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_4),
.C(n_7),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_40),
.B(n_22),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_26),
.B(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_15),
.B1(n_20),
.B2(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_56),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_20),
.B1(n_10),
.B2(n_9),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_36),
.B1(n_37),
.B2(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_52),
.B1(n_59),
.B2(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_67),
.B1(n_64),
.B2(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_20),
.B1(n_33),
.B2(n_11),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_77),
.B1(n_47),
.B2(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_9),
.B1(n_33),
.B2(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_84),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_42),
.C(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_41),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_52),
.B(n_75),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_78),
.B(n_63),
.C(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_87),
.C(n_91),
.Y(n_104)
);

XOR2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_63),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_90),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_90),
.B1(n_89),
.B2(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_105),
.B1(n_93),
.B2(n_106),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_96),
.C(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_117),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_112),
.B(n_118),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_122),
.C(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_109),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_96),
.B(n_97),
.C(n_95),
.D(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_100),
.Y(n_125)
);


endmodule