module fake_jpeg_13127_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_17),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_35),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_12),
.B1(n_21),
.B2(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_20),
.B1(n_25),
.B2(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_30),
.B1(n_18),
.B2(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_48),
.B1(n_52),
.B2(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_24),
.B1(n_23),
.B2(n_14),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_24),
.C(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_37),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_16),
.B2(n_23),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_59),
.B1(n_41),
.B2(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_20),
.B1(n_41),
.B2(n_40),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_4),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_65),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.C(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_42),
.C(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_42),
.B1(n_20),
.B2(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_63),
.B1(n_64),
.B2(n_60),
.C(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_70),
.C(n_68),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_55),
.B1(n_59),
.B2(n_8),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.C(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);


endmodule