module fake_jpeg_22729_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_34),
.B1(n_22),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_51),
.B1(n_57),
.B2(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_20),
.B(n_32),
.C(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_17),
.B1(n_31),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_17),
.B1(n_35),
.B2(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_19),
.B1(n_25),
.B2(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_68),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_30),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_76),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_80),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_74),
.Y(n_103)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_17),
.B1(n_31),
.B2(n_27),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_43),
.B1(n_35),
.B2(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_17),
.B1(n_43),
.B2(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_42),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_101),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_117),
.Y(n_127)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_68),
.A3(n_64),
.B1(n_50),
.B2(n_27),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_113),
.C(n_120),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_43),
.B1(n_51),
.B2(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_82),
.B1(n_71),
.B2(n_79),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_73),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_65),
.B1(n_58),
.B2(n_38),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_116),
.B1(n_79),
.B2(n_70),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_58),
.B1(n_38),
.B2(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_0),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_122),
.B(n_33),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_42),
.C(n_40),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_16),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_92),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_56),
.B(n_42),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_107),
.B(n_85),
.C(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_133),
.A2(n_29),
.B(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_140),
.B1(n_147),
.B2(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_126),
.B(n_138),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_94),
.B1(n_88),
.B2(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_78),
.B1(n_60),
.B2(n_23),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_60),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_99),
.B1(n_115),
.B2(n_97),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_146),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_102),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_159),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_120),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_162),
.C(n_166),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_104),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_144),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_117),
.B1(n_119),
.B2(n_98),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_118),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_137),
.C(n_125),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_118),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_178),
.C(n_151),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_106),
.B1(n_100),
.B2(n_96),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_95),
.B1(n_61),
.B2(n_67),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_180),
.B(n_42),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_42),
.C(n_40),
.Y(n_178)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.C(n_21),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_42),
.B(n_40),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_13),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_11),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_134),
.C(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_207),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_191),
.B(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_188),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_130),
.C(n_143),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_209),
.C(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_197),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_143),
.B1(n_67),
.B2(n_61),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_201),
.B1(n_164),
.B2(n_95),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

OAI322xp33_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_176),
.A3(n_167),
.B1(n_169),
.B2(n_153),
.C1(n_179),
.C2(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_124),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_42),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_40),
.C(n_95),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_171),
.B1(n_181),
.B2(n_175),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_161),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_194),
.B(n_0),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_221),
.C(n_229),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_187),
.B(n_195),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_194),
.B(n_2),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_159),
.C(n_166),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_162),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_180),
.B1(n_29),
.B2(n_24),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_24),
.B1(n_23),
.B2(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_40),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_40),
.C(n_21),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_18),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_2),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_0),
.C(n_1),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_202),
.C(n_204),
.Y(n_243)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_247),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_208),
.B(n_188),
.C(n_210),
.D(n_196),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_186),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_225),
.B(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_256),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_236),
.B1(n_238),
.B2(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_242),
.C(n_223),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_271),
.C(n_218),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_262),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_240),
.B1(n_235),
.B2(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_265),
.B1(n_4),
.B2(n_5),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_249),
.B1(n_239),
.B2(n_244),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_227),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_216),
.C(n_229),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_231),
.B(n_250),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_255),
.C(n_245),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_222),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_230),
.C(n_226),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_271),
.B(n_272),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_252),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_7),
.B(n_8),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_224),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_270),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_283),
.C(n_9),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_269),
.B(n_272),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_298),
.B(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_257),
.B1(n_266),
.B2(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_9),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_8),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_278),
.B(n_281),
.Y(n_299)
);

AOI311xp33_ASAP7_75t_SL g311 ( 
.A1(n_299),
.A2(n_306),
.A3(n_10),
.B(n_12),
.C(n_13),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_15),
.C(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_8),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_298),
.A3(n_307),
.B1(n_288),
.B2(n_292),
.C1(n_306),
.C2(n_304),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_293),
.C(n_11),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B(n_10),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_293),
.B1(n_12),
.B2(n_13),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_12),
.B1(n_15),
.B2(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_15),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.Y(n_322)
);


endmodule