module fake_aes_560_n_676 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_676);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_676;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_69), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_22), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_23), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_14), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_11), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_76), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_57), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_70), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_34), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_68), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_17), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_71), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_48), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_49), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_52), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_55), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_43), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_16), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_67), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_12), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_15), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_2), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_1), .Y(n_120) );
INVxp33_ASAP7_75t_SL g121 ( .A(n_18), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_39), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_10), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_66), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_123), .B(n_0), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_109), .B(n_0), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_87), .B(n_1), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_113), .B(n_2), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_113), .B(n_81), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_81), .B(n_4), .Y(n_138) );
CKINVDCx11_ASAP7_75t_R g139 ( .A(n_82), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_106), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_88), .A2(n_32), .B(n_74), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_83), .B(n_84), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
NOR2xp33_ASAP7_75t_SL g155 ( .A(n_79), .B(n_30), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_98), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_99), .B(n_5), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_122), .Y(n_159) );
BUFx8_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_118), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_84), .Y(n_164) );
AND3x2_ASAP7_75t_L g165 ( .A(n_94), .B(n_5), .C(n_6), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_101), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_103), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_159), .B(n_100), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_136), .B(n_107), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_137), .B(n_92), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
CKINVDCx8_ASAP7_75t_R g180 ( .A(n_140), .Y(n_180) );
CKINVDCx8_ASAP7_75t_R g181 ( .A(n_140), .Y(n_181) );
AND2x6_ASAP7_75t_L g182 ( .A(n_136), .B(n_110), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_137), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_148), .B(n_89), .Y(n_187) );
OR2x6_ASAP7_75t_L g188 ( .A(n_130), .B(n_111), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_164), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_160), .B(n_112), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_132), .A2(n_121), .B1(n_120), .B2(n_102), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_164), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_125), .B(n_105), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_132), .B(n_97), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_149), .B(n_119), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_137), .B(n_119), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
INVx8_ASAP7_75t_L g201 ( .A(n_132), .Y(n_201) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_125), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_160), .B(n_104), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_141), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_141), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
NAND3x1_ASAP7_75t_L g208 ( .A(n_130), .B(n_92), .C(n_93), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_149), .A2(n_93), .B1(n_114), .B2(n_111), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_141), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_150), .B(n_114), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_138), .A2(n_96), .B1(n_115), .B2(n_85), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_150), .B(n_96), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_141), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_128), .B(n_108), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
AND2x6_ASAP7_75t_L g220 ( .A(n_143), .B(n_117), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_152), .B(n_6), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_161), .B(n_33), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_152), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_128), .B(n_7), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_224), .B(n_162), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_189), .A2(n_142), .B(n_161), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_221), .A2(n_161), .B1(n_134), .B2(n_129), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_224), .B(n_139), .Y(n_235) );
CKINVDCx11_ASAP7_75t_R g236 ( .A(n_180), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_202), .B(n_143), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_184), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_153), .B1(n_129), .B2(n_134), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_184), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_195), .B(n_153), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_208), .A2(n_162), .B1(n_156), .B2(n_163), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_186), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_188), .A2(n_138), .B1(n_163), .B2(n_156), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_221), .A2(n_143), .B1(n_166), .B2(n_126), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_183), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_221), .Y(n_248) );
AND3x2_ASAP7_75t_SL g249 ( .A(n_180), .B(n_165), .C(n_126), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_218), .B(n_166), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_201), .B(n_143), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_187), .B(n_211), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_201), .B(n_166), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_201), .B(n_146), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_201), .B(n_146), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_200), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_205), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_192), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_227), .Y(n_263) );
CKINVDCx6p67_ASAP7_75t_R g264 ( .A(n_215), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_174), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_176), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_193), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_181), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_176), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_202), .B(n_147), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_211), .B(n_146), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_181), .Y(n_272) );
AND3x2_ASAP7_75t_SL g273 ( .A(n_208), .B(n_165), .C(n_126), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_211), .B(n_127), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_175), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_214), .B(n_127), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_127), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_175), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_182), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_199), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_214), .B(n_131), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_172), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_174), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_174), .Y(n_287) );
OAI21xp33_ASAP7_75t_L g288 ( .A1(n_196), .A2(n_194), .B(n_188), .Y(n_288) );
AND2x6_ASAP7_75t_L g289 ( .A(n_175), .B(n_131), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_188), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_182), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_284), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_289), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_259), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
AND2x2_ASAP7_75t_SL g298 ( .A(n_246), .B(n_234), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_248), .A2(n_220), .B1(n_182), .B2(n_188), .Y(n_299) );
INVx5_ASAP7_75t_L g300 ( .A(n_233), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_252), .B(n_220), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_252), .A2(n_178), .B(n_202), .C(n_196), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_212), .B1(n_209), .B2(n_191), .C(n_217), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_228), .B(n_220), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_236), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_290), .B(n_220), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_245), .B(n_220), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_235), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_263), .B(n_172), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_233), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_242), .B(n_220), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_265), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
INVx5_ASAP7_75t_L g318 ( .A(n_233), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_288), .A2(n_182), .B1(n_172), .B2(n_178), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_261), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_232), .B(n_178), .Y(n_321) );
OAI21xp33_ASAP7_75t_SL g322 ( .A1(n_243), .A2(n_203), .B(n_142), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_264), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_265), .Y(n_324) );
OR2x2_ASAP7_75t_SL g325 ( .A(n_236), .B(n_131), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_266), .A2(n_182), .B1(n_190), .B2(n_171), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_264), .B(n_144), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_240), .B(n_135), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_271), .A2(n_151), .B1(n_144), .B2(n_157), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_254), .B(n_158), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_261), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_269), .B(n_151), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_274), .A2(n_167), .B1(n_145), .B2(n_144), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_281), .B(n_151), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_256), .B(n_145), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_267), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_239), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_322), .A2(n_250), .B(n_230), .C(n_257), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_298), .A2(n_282), .B1(n_285), .B2(n_244), .Y(n_344) );
CKINVDCx6p67_ASAP7_75t_R g345 ( .A(n_323), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_292), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_308), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_303), .A2(n_250), .B1(n_275), .B2(n_283), .C(n_278), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_298), .A2(n_244), .B1(n_229), .B2(n_272), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_298), .A2(n_244), .B1(n_229), .B2(n_272), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_292), .B(n_268), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_332), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_268), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_322), .A2(n_251), .B(n_277), .C(n_260), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_328), .A2(n_259), .B1(n_291), .B2(n_249), .Y(n_357) );
BUFx12f_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_312), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_313), .B(n_309), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_309), .A2(n_229), .B1(n_289), .B2(n_287), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_309), .B(n_232), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_299), .A2(n_291), .B1(n_259), .B2(n_280), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_309), .B(n_259), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_299), .A2(n_280), .B1(n_232), .B2(n_249), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_329), .A2(n_255), .B1(n_241), .B2(n_238), .C(n_231), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_300), .B(n_232), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_293), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_358), .A2(n_310), .B1(n_330), .B2(n_320), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_343), .A2(n_310), .B(n_302), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_360), .A2(n_301), .B1(n_307), .B2(n_315), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_358), .A2(n_330), .B1(n_301), .B2(n_339), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_355), .A2(n_341), .B(n_339), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_346), .B(n_300), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_362), .B1(n_360), .B2(n_356), .C(n_344), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_315), .B1(n_331), .B2(n_338), .C(n_333), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_341), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_372), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_346), .B(n_341), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_372), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_326), .B(n_319), .C(n_337), .Y(n_389) );
AOI221xp5_ASAP7_75t_SL g390 ( .A1(n_349), .A2(n_325), .B1(n_237), .B2(n_338), .C(n_270), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_351), .A2(n_304), .B1(n_306), .B2(n_336), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_361), .B(n_145), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_361), .B(n_340), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_370), .A2(n_294), .B1(n_305), .B2(n_311), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_304), .B1(n_336), .B2(n_293), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_350), .A2(n_237), .B1(n_157), .B2(n_296), .C(n_327), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_361), .A2(n_305), .B1(n_294), .B2(n_311), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_369), .A2(n_324), .B1(n_335), .B2(n_316), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_353), .A2(n_324), .B1(n_335), .B2(n_316), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_157), .B1(n_297), .B2(n_342), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_353), .A2(n_306), .B1(n_334), .B2(n_155), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_354), .A2(n_297), .B(n_342), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_383), .B(n_273), .C(n_363), .D(n_155), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_345), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_393), .B(n_345), .Y(n_406) );
INVxp67_ASAP7_75t_R g407 ( .A(n_392), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_387), .B(n_354), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_388), .A2(n_373), .B1(n_374), .B2(n_367), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_375), .B(n_373), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_147), .B1(n_154), .B2(n_167), .C(n_347), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_382), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_397), .B(n_367), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_374), .B(n_359), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_390), .B(n_167), .C(n_147), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_384), .A2(n_368), .B1(n_154), .B2(n_147), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_397), .B(n_368), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_375), .A2(n_368), .B1(n_327), .B2(n_296), .C(n_335), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_379), .B(n_368), .Y(n_422) );
OAI21x1_ASAP7_75t_L g423 ( .A1(n_402), .A2(n_371), .B(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_394), .B(n_365), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_394), .B(n_295), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_400), .B(n_295), .Y(n_427) );
OAI211xp5_ASAP7_75t_SL g428 ( .A1(n_379), .A2(n_223), .B(n_270), .C(n_273), .Y(n_428) );
AOI33xp33_ASAP7_75t_L g429 ( .A1(n_391), .A2(n_170), .A3(n_179), .B1(n_185), .B2(n_207), .B3(n_210), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_400), .B(n_297), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_154), .B1(n_167), .B2(n_347), .C(n_253), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_389), .A2(n_321), .B(n_142), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_378), .A2(n_335), .B1(n_327), .B2(n_324), .C(n_296), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_395), .A2(n_334), .B1(n_359), .B2(n_296), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_365), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_359), .B1(n_380), .B2(n_300), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_405), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_422), .B(n_380), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_412), .B1(n_422), .B2(n_421), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_415), .B(n_154), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_418), .A2(n_409), .B1(n_436), .B2(n_407), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_428), .A2(n_365), .B1(n_154), .B2(n_167), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_413), .B(n_154), .C(n_167), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_434), .B(n_359), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_408), .B(n_154), .Y(n_449) );
AOI21xp33_ASAP7_75t_SL g450 ( .A1(n_406), .A2(n_7), .B(n_8), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_414), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_435), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_417), .B(n_167), .C(n_318), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_426), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_428), .A2(n_327), .B1(n_324), .B2(n_316), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_411), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_406), .A2(n_316), .B1(n_318), .B2(n_300), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_424), .B(n_9), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_411), .B(n_10), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_429), .B(n_418), .C(n_432), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_419), .B(n_300), .Y(n_462) );
OAI211xp5_ASAP7_75t_L g463 ( .A1(n_404), .A2(n_321), .B(n_300), .C(n_318), .Y(n_463) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_425), .A2(n_170), .A3(n_179), .B1(n_185), .B2(n_207), .B3(n_210), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_430), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_437), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_409), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_431), .A2(n_318), .B1(n_314), .B2(n_258), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_427), .Y(n_471) );
INVx5_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_433), .B(n_11), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_429), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_403), .A2(n_239), .B1(n_253), .B2(n_226), .C(n_216), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_405), .B(n_318), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_405), .B(n_12), .Y(n_477) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_417), .A2(n_213), .B(n_216), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_405), .B(n_13), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_408), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_405), .B(n_14), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_405), .B(n_318), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_405), .B(n_18), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_405), .B(n_19), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_454), .B(n_19), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_454), .B(n_20), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_441), .A2(n_371), .B1(n_21), .B2(n_314), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_454), .B(n_21), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_481), .Y(n_493) );
OAI222xp33_ASAP7_75t_L g494 ( .A1(n_444), .A2(n_371), .B1(n_280), .B2(n_232), .C1(n_286), .C2(n_226), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_465), .B(n_24), .Y(n_495) );
NOR3xp33_ASAP7_75t_SL g496 ( .A(n_444), .B(n_213), .C(n_25), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_479), .B(n_314), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_448), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_448), .Y(n_499) );
AND2x4_ASAP7_75t_SL g500 ( .A(n_451), .B(n_314), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_457), .Y(n_501) );
AND2x4_ASAP7_75t_SL g502 ( .A(n_482), .B(n_314), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_471), .B(n_204), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_465), .B(n_26), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_442), .B(n_204), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_460), .A2(n_222), .A3(n_219), .B(n_206), .Y(n_507) );
NAND2x1_ASAP7_75t_SL g508 ( .A(n_467), .B(n_222), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_442), .B(n_219), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_450), .B(n_486), .C(n_485), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_452), .B(n_206), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_440), .B(n_471), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_440), .B(n_28), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_452), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_440), .B(n_29), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_466), .B(n_198), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_457), .B(n_258), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_466), .B(n_198), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
OAI211xp5_ASAP7_75t_SL g521 ( .A1(n_475), .A2(n_169), .B(n_168), .C(n_286), .Y(n_521) );
INVxp67_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_450), .B(n_225), .C(n_173), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_479), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_440), .B(n_35), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_466), .B(n_37), .Y(n_526) );
OAI211xp5_ASAP7_75t_SL g527 ( .A1(n_475), .A2(n_169), .B(n_168), .C(n_286), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_443), .B(n_225), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_447), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_474), .A2(n_258), .B1(n_233), .B2(n_225), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_477), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_467), .B(n_38), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_443), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_477), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_462), .B(n_225), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_480), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_462), .B(n_225), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_480), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_459), .B(n_173), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_483), .Y(n_540) );
OAI31xp33_ASAP7_75t_SL g541 ( .A1(n_438), .A2(n_40), .A3(n_41), .B(n_42), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_476), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
AOI322xp5_ASAP7_75t_L g545 ( .A1(n_510), .A2(n_486), .A3(n_485), .B1(n_483), .B2(n_459), .C1(n_474), .C2(n_468), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_498), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_522), .B(n_473), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_512), .B(n_468), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_512), .B(n_455), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_491), .A2(n_474), .B1(n_438), .B2(n_473), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_488), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_501), .B(n_461), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_542), .B(n_476), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_498), .B(n_455), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_523), .A2(n_453), .B(n_461), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_502), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_531), .B(n_449), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_488), .B(n_455), .Y(n_559) );
CKINVDCx6p67_ASAP7_75t_R g560 ( .A(n_520), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_499), .B(n_484), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_489), .B(n_484), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_493), .B(n_472), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_445), .B(n_449), .Y(n_565) );
NAND2x1_ASAP7_75t_L g566 ( .A(n_520), .B(n_453), .Y(n_566) );
NOR3xp33_ASAP7_75t_SL g567 ( .A(n_494), .B(n_463), .C(n_446), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_493), .B(n_472), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_502), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_524), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_524), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_534), .B(n_472), .Y(n_572) );
AOI21xp33_ASAP7_75t_L g573 ( .A1(n_541), .A2(n_472), .B(n_458), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_520), .A2(n_472), .B1(n_446), .B2(n_478), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_536), .B(n_458), .C(n_456), .D(n_464), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_515), .B(n_472), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_529), .B(n_472), .Y(n_578) );
NAND3xp33_ASAP7_75t_SL g579 ( .A(n_507), .B(n_470), .C(n_47), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_529), .B(n_447), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_487), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_538), .B(n_447), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_533), .B(n_447), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_540), .B(n_478), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_492), .B(n_478), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_492), .B(n_478), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_533), .B(n_173), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_490), .B(n_46), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_495), .B(n_173), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_490), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_553), .B(n_539), .C(n_537), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_546), .B(n_537), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_543), .Y(n_593) );
AOI21xp33_ASAP7_75t_SL g594 ( .A1(n_573), .A2(n_497), .B(n_525), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_549), .B(n_535), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_560), .A2(n_500), .B1(n_497), .B2(n_532), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_544), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_545), .A2(n_500), .B(n_508), .C(n_532), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_574), .B(n_497), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_576), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_550), .B(n_549), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_553), .B(n_504), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_581), .B(n_495), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_554), .B(n_535), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_548), .B(n_508), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_552), .Y(n_606) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_551), .A2(n_525), .B(n_514), .C(n_516), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_563), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_590), .B(n_526), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_577), .B(n_526), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_560), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_570), .B(n_528), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_561), .B(n_571), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_582), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_548), .B(n_503), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_558), .B(n_572), .Y(n_617) );
NAND2x1_ASAP7_75t_SL g618 ( .A(n_578), .B(n_516), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_547), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_584), .B(n_503), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_559), .B(n_514), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_559), .B(n_528), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_556), .A2(n_518), .B(n_527), .Y(n_623) );
OAI321xp33_ASAP7_75t_L g624 ( .A1(n_579), .A2(n_521), .A3(n_519), .B1(n_517), .B2(n_509), .C(n_505), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_555), .Y(n_625) );
AOI31xp33_ASAP7_75t_L g626 ( .A1(n_569), .A2(n_530), .A3(n_511), .B(n_58), .Y(n_626) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_569), .B(n_54), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_555), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_567), .A2(n_56), .B(n_60), .C(n_61), .Y(n_629) );
NAND4xp75_ASAP7_75t_L g630 ( .A(n_578), .B(n_63), .C(n_64), .D(n_65), .Y(n_630) );
AOI211x1_ASAP7_75t_SL g631 ( .A1(n_575), .A2(n_173), .B(n_75), .C(n_73), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_580), .B(n_258), .Y(n_632) );
AO22x2_ASAP7_75t_L g633 ( .A1(n_564), .A2(n_280), .B1(n_568), .B2(n_580), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_587), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_557), .A2(n_280), .B1(n_566), .B2(n_565), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_585), .B(n_586), .C(n_568), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_583), .B(n_564), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_588), .A2(n_560), .B1(n_551), .B2(n_441), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_587), .B(n_589), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_639), .A2(n_607), .B1(n_605), .B2(n_611), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_613), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_636), .B(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
INVx2_ASAP7_75t_SL g645 ( .A(n_592), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_594), .B(n_598), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_598), .A2(n_635), .B1(n_599), .B2(n_628), .C(n_625), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_628), .A2(n_615), .B1(n_614), .B2(n_616), .C(n_637), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_599), .A2(n_605), .B(n_624), .C(n_596), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_633), .A2(n_595), .B1(n_604), .B2(n_591), .Y(n_650) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_593), .A2(n_597), .B1(n_600), .B2(n_612), .Y(n_651) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_629), .A2(n_626), .B(n_620), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_612), .Y(n_653) );
AOI31xp33_ASAP7_75t_L g654 ( .A1(n_627), .A2(n_623), .A3(n_602), .B(n_601), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_650), .A2(n_633), .B1(n_623), .B2(n_601), .C(n_608), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_641), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_644), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_654), .A2(n_629), .B(n_632), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_618), .B(n_638), .C(n_610), .Y(n_659) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_646), .B(n_633), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_653), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_647), .A2(n_640), .B1(n_622), .B2(n_606), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_655), .A2(n_651), .B1(n_648), .B2(n_652), .C(n_643), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_656), .A2(n_651), .B1(n_642), .B2(n_645), .Y(n_664) );
XNOR2x1_ASAP7_75t_L g665 ( .A(n_660), .B(n_630), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g666 ( .A1(n_662), .A2(n_631), .B1(n_621), .B2(n_603), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_661), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_667), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_666), .A2(n_658), .B1(n_657), .B2(n_634), .Y(n_669) );
XOR2xp5_ASAP7_75t_L g670 ( .A(n_665), .B(n_609), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_668), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_670), .B(n_663), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_671), .B(n_669), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_673), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_674), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_672), .B1(n_664), .B2(n_659), .C(n_619), .Y(n_676) );
endmodule