module real_jpeg_15650_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_535),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_0),
.B(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_1),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_1),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_1),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_1),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_1),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_1),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_3),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_3),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_3),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_4),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_4),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_5),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_5),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g323 ( 
.A(n_5),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_5),
.B(n_420),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_5),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_6),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_6),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_6),
.B(n_52),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_7),
.B(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_7),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_7),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_7),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_7),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_9),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_10),
.Y(n_536)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_12),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_12),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_12),
.B(n_145),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_12),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_12),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_12),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_12),
.B(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_15),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_16),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_16),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_16),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_16),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_16),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_16),
.B(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_16),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_520),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_253),
.B(n_514),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_205),
.C(n_248),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_166),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_24),
.B(n_166),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_99),
.C(n_132),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_26),
.B(n_99),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_70),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_71),
.C(n_91),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_45),
.C(n_61),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_28),
.B(n_45),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_29),
.B(n_178),
.C(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_39),
.B(n_43),
.C(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_42),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_60),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_55),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_47),
.A2(n_49),
.B1(n_68),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_47),
.B(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_47),
.A2(n_136),
.B1(n_314),
.B2(n_315),
.Y(n_375)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_48),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_48),
.Y(n_457)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_48),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_62),
.C(n_69),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_49),
.B(n_419),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_50),
.B(n_143),
.Y(n_142)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g178 ( 
.A(n_51),
.B(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_52),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_52),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_135),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_58),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_60),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_60),
.A2(n_346),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_61),
.B(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_62),
.A2(n_165),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_62),
.B(n_165),
.Y(n_530)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_69),
.B1(n_102),
.B2(n_106),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_65),
.B(n_158),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_67),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_68),
.B(n_419),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_69),
.B(n_107),
.C(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_91),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_84),
.C(n_86),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_72),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.C(n_80),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_73),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_73),
.B(n_192),
.C(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_80),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_76),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_98),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_86),
.B(n_94),
.C(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_86),
.A2(n_87),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_87),
.B(n_209),
.C(n_215),
.Y(n_234)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_92),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_94),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2x2_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_115),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_100),
.B(n_116),
.C(n_118),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_102),
.A2(n_106),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_102),
.B(n_172),
.C(n_178),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_102),
.B(n_322),
.C(n_323),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_102),
.A2(n_106),
.B1(n_322),
.B2(n_374),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_103),
.Y(n_488)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_112),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_113),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_113),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_117),
.B(n_177),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_119),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_119),
.A2(n_185),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_119),
.B(n_142),
.C(n_165),
.Y(n_526)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_126),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_138),
.C(n_142),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_131),
.C(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_127),
.A2(n_130),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_129),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_132),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_148),
.C(n_152),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_133),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_146),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_134),
.B(n_137),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_225),
.Y(n_332)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_142),
.A2(n_177),
.B1(n_178),
.B2(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_146),
.Y(n_335)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_150),
.Y(n_298)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_161),
.C(n_165),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_154),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_159),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_155),
.B(n_158),
.Y(n_262)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_159),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_161),
.A2(n_165),
.B1(n_240),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_161),
.Y(n_294)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_164),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_165),
.A2(n_225),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_167),
.B(n_170),
.C(n_186),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_186),
.B2(n_187),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2x2_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_182),
.C(n_184),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_174),
.Y(n_353)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_218),
.C(n_239),
.Y(n_245)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_204),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_201),
.B2(n_202),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_202),
.C(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_191),
.A2(n_192),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_198),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_205),
.A2(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_231),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_206),
.B(n_231),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_227),
.C(n_228),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_227),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_217),
.C(n_226),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_232),
.B(n_234),
.C(n_235),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_236),
.B(n_245),
.C(n_246),
.Y(n_524)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_249),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_250),
.B(n_252),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_397),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_336),
.B(n_389),
.C(n_390),
.D(n_396),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_256),
.B(n_391),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_303),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_257),
.B(n_303),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_295),
.Y(n_257)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_258),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_279),
.C(n_290),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.C(n_270),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_261),
.B(n_356),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_263),
.A2(n_264),
.B1(n_270),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_264),
.A2(n_265),
.B(n_267),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_270),
.Y(n_357)
);

MAJx3_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_271),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_273),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_276),
.Y(n_311)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_279),
.A2(n_291),
.B1(n_292),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_281),
.B(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_286),
.Y(n_329)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_299),
.B(n_301),
.C(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_333),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_333),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_328),
.C(n_330),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_321),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_312),
.A2(n_313),
.B1(n_321),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_319),
.Y(n_494)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_322),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_323),
.B(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_327),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_330),
.Y(n_340)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_360),
.B(n_388),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_358),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_358),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.C(n_354),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_355),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.C(n_345),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_344),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.C(n_350),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_347),
.A2(n_350),
.B1(n_351),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_347),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_363),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.C(n_371),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_364),
.A2(n_365),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_367),
.A2(n_368),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.C(n_376),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_372),
.B(n_375),
.C(n_376),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_376),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_380),
.C(n_386),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_377),
.A2(n_378),
.B1(n_386),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_380),
.B(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_386),
.Y(n_449)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_394),
.Y(n_396)
);

NAND4xp25_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_399),
.C(n_400),
.D(n_401),
.Y(n_397)
);

OAI21x1_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_505),
.B(n_513),
.Y(n_401)
);

AOI21x1_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_450),
.B(n_504),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_426),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_426),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_424),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_410),
.C(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.C(n_418),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_411),
.A2(n_412),
.B1(n_413),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_428),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.C(n_447),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_465),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_447),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_443),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_439),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_466),
.B(n_503),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_464),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_452),
.B(n_464),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_462),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_500),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_455),
.A2(n_462),
.B1(n_463),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_455),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_458),
.Y(n_476)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_497),
.B(n_502),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_485),
.B(n_496),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_475),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_469),
.B(n_475),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_473),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_479),
.C(n_482),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_483),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_490),
.B(n_495),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_489),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_499),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_511),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_511),
.Y(n_513)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_534),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_533),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_533),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_527),
.B1(n_531),
.B2(n_532),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_526),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule