module real_jpeg_30199_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_18),
.B(n_20),
.C(n_21),
.D(n_28),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_25),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_1),
.A2(n_25),
.B(n_36),
.C(n_77),
.D(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_1),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_55),
.B(n_70),
.Y(n_101)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_4),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_5),
.A2(n_41),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_69)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_7),
.B(n_25),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_38),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_41),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_9),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_73),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_60),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_60),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_47),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_32),
.Y(n_16)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI32xp33_ASAP7_75t_L g57 ( 
.A1(n_19),
.A2(n_20),
.A3(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_24),
.B(n_26),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_24),
.A2(n_38),
.A3(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_40),
.B2(n_45),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_53),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_44),
.B(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_54),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_88),
.B(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.C(n_68),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_84),
.B(n_108),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_81),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_94),
.B(n_107),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_93),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_100),
.B(n_106),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);


endmodule