module fake_aes_9310_n_20 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_0), .A2(n_9), .B1(n_10), .B2(n_7), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_3), .B(n_4), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_1), .B(n_5), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_15), .B(n_13), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_16), .B1(n_11), .B2(n_15), .C(n_6), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_19) );
AOI222xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_2), .B1(n_6), .B2(n_7), .C1(n_8), .C2(n_18), .Y(n_20) );
endmodule