module fake_jpeg_19067_n_235 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx8_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_14),
.B1(n_22),
.B2(n_21),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_16),
.B(n_25),
.Y(n_51)
);

XOR2x1_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_65),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_44),
.B(n_40),
.C(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_59),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_35),
.B1(n_29),
.B2(n_45),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_27),
.B(n_26),
.C(n_17),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_32),
.B1(n_37),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_70),
.B1(n_79),
.B2(n_63),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_28),
.B1(n_16),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_81),
.B1(n_80),
.B2(n_35),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_25),
.C(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_76),
.B1(n_68),
.B2(n_71),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_57),
.C(n_59),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_38),
.C(n_29),
.Y(n_116)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_56),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_82),
.B1(n_63),
.B2(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_53),
.B(n_55),
.C(n_56),
.D(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_109),
.B1(n_115),
.B2(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_82),
.B1(n_83),
.B2(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_85),
.B1(n_94),
.B2(n_65),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_53),
.B1(n_49),
.B2(n_78),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_48),
.B(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_49),
.B1(n_16),
.B2(n_13),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_49),
.B1(n_43),
.B2(n_42),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_31),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_31),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_115),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_100),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_131),
.B(n_48),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_123),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_135),
.C(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_129),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_75),
.B1(n_43),
.B2(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_21),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_117),
.C(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_31),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_75),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_38),
.C(n_45),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_18),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_58),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_54),
.B1(n_42),
.B2(n_58),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_33),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_54),
.B1(n_87),
.B2(n_19),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_127),
.B1(n_19),
.B2(n_13),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_135),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_48),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_15),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_87),
.C(n_34),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_123),
.C(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_173),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_157),
.C(n_155),
.Y(n_167)
);

BUFx12f_ASAP7_75t_SL g184 ( 
.A(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_158),
.B(n_149),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_24),
.C(n_33),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_24),
.C(n_20),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_159),
.B1(n_144),
.B2(n_18),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_141),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_147),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_189),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_143),
.B1(n_153),
.B2(n_154),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_15),
.B1(n_8),
.B2(n_12),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_163),
.C(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_194),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_188),
.B(n_146),
.CI(n_172),
.CON(n_193),
.SN(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_174),
.C(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_167),
.C(n_15),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_198),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_20),
.C(n_7),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_20),
.C(n_7),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_176),
.C(n_185),
.Y(n_209)
);

OAI321xp33_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_197),
.A3(n_193),
.B1(n_8),
.B2(n_9),
.C(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_189),
.B(n_176),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_210),
.B(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_186),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_196),
.C(n_201),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_218),
.C(n_10),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_219),
.B(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_9),
.B1(n_10),
.B2(n_2),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_9),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_0),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_0),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_214),
.B(n_1),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_229),
.C(n_222),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_1),
.C(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_228),
.B(n_1),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_3),
.C(n_103),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_234),
.B(n_3),
.Y(n_235)
);


endmodule