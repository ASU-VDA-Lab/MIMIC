module fake_jpeg_16883_n_55 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_18),
.B(n_17),
.C(n_16),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_26),
.B(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_25),
.B1(n_23),
.B2(n_4),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_28),
.B1(n_5),
.B2(n_6),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

AND2x4_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_23),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_24),
.C(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_34),
.B2(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_49),
.B1(n_41),
.B2(n_8),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_51),
.B(n_48),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_45),
.Y(n_54)
);

OAI321xp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_8),
.A3(n_9),
.B1(n_45),
.B2(n_46),
.C(n_53),
.Y(n_55)
);


endmodule