module fake_jpeg_4257_n_148 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_32),
.Y(n_53)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_24),
.B1(n_17),
.B2(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_19),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_2),
.Y(n_39)
);

NOR2x1_ASAP7_75t_R g48 ( 
.A(n_39),
.B(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_20),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_27),
.B(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_18),
.B1(n_14),
.B2(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_42),
.C(n_11),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_50),
.C(n_51),
.Y(n_93)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_82),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_87),
.B1(n_67),
.B2(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_95),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_54),
.B(n_44),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_77),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_47),
.Y(n_100)
);

XOR2x2_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_43),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_73),
.A3(n_77),
.B1(n_59),
.B2(n_58),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_66),
.B(n_53),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_79),
.B1(n_75),
.B2(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_82),
.B1(n_60),
.B2(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_93),
.B(n_89),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_92),
.B(n_100),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_126),
.B(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_97),
.C(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_125),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_114),
.B1(n_113),
.B2(n_107),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_96),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_91),
.B(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_104),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_130),
.B(n_109),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_110),
.B1(n_108),
.B2(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_111),
.B1(n_78),
.B2(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_138),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_104),
.B(n_111),
.Y(n_136)
);

AOI31xp67_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_129),
.A3(n_134),
.B(n_7),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_7),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_128),
.C(n_132),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_145),
.B1(n_8),
.B2(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_8),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);


endmodule