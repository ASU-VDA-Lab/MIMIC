module real_aes_15563_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g823 ( .A(n_0), .B(n_824), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_1), .A2(n_4), .B1(n_271), .B2(n_272), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_2), .A2(n_42), .B1(n_128), .B2(n_198), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_3), .A2(n_23), .B1(n_198), .B2(n_207), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_5), .A2(n_15), .B1(n_504), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_6), .A2(n_59), .B1(n_156), .B2(n_157), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_7), .A2(n_16), .B1(n_128), .B2(n_130), .Y(n_127) );
INVx1_ASAP7_75t_L g824 ( .A(n_8), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_9), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_10), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_11), .A2(n_17), .B1(n_505), .B2(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g110 ( .A(n_12), .B(n_37), .Y(n_110) );
BUFx2_ASAP7_75t_L g818 ( .A(n_12), .Y(n_818) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_13), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_14), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_18), .A2(n_97), .B1(n_272), .B2(n_504), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_19), .A2(n_38), .B1(n_164), .B2(n_521), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_20), .B(n_163), .Y(n_518) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_21), .A2(n_57), .B(n_141), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_22), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_24), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_25), .B(n_133), .Y(n_227) );
INVx4_ASAP7_75t_R g180 ( .A(n_26), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_27), .A2(n_46), .B1(n_135), .B2(n_269), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_28), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_29), .A2(n_52), .B1(n_135), .B2(n_504), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_30), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_31), .B(n_521), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_32), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_33), .B(n_198), .Y(n_233) );
INVx1_ASAP7_75t_L g276 ( .A(n_34), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_SL g204 ( .A1(n_35), .A2(n_128), .B(n_132), .C(n_205), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_36), .A2(n_54), .B1(n_128), .B2(n_135), .Y(n_216) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_37), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_39), .A2(n_85), .B1(n_128), .B2(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_40), .A2(n_113), .B1(n_114), .B2(n_786), .Y(n_112) );
INVx1_ASAP7_75t_L g786 ( .A(n_40), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_41), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_43), .A2(n_45), .B1(n_128), .B2(n_130), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_44), .A2(n_58), .B1(n_504), .B2(n_556), .Y(n_572) );
INVx1_ASAP7_75t_L g230 ( .A(n_47), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_48), .B(n_128), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_49), .Y(n_249) );
INVx2_ASAP7_75t_L g791 ( .A(n_50), .Y(n_791) );
INVx1_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
BUFx3_ASAP7_75t_L g794 ( .A(n_51), .Y(n_794) );
INVx1_ASAP7_75t_L g801 ( .A(n_53), .Y(n_801) );
AOI31xp33_ASAP7_75t_L g804 ( .A1(n_53), .A2(n_101), .A3(n_103), .B(n_805), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_55), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_56), .A2(n_86), .B1(n_128), .B2(n_135), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_60), .A2(n_74), .B1(n_269), .B2(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_61), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_62), .A2(n_77), .B1(n_128), .B2(n_130), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_63), .A2(n_96), .B1(n_504), .B2(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
AND2x4_ASAP7_75t_L g143 ( .A(n_65), .B(n_144), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_66), .A2(n_88), .B1(n_135), .B2(n_269), .Y(n_268) );
AO22x1_ASAP7_75t_L g161 ( .A1(n_67), .A2(n_75), .B1(n_162), .B2(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g144 ( .A(n_68), .Y(n_144) );
AND2x2_ASAP7_75t_L g208 ( .A(n_69), .B(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_70), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_71), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_72), .B(n_156), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_73), .A2(n_100), .B1(n_814), .B2(n_825), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_76), .B(n_198), .Y(n_250) );
INVx2_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_79), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_80), .B(n_209), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_81), .A2(n_95), .B1(n_135), .B2(n_156), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_82), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_83), .B(n_139), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_84), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_87), .B(n_209), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_89), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_90), .B(n_209), .Y(n_246) );
INVx1_ASAP7_75t_L g108 ( .A(n_91), .Y(n_108) );
NAND2xp33_ASAP7_75t_L g522 ( .A(n_92), .B(n_163), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_93), .A2(n_137), .B(n_156), .C(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g185 ( .A(n_94), .B(n_186), .Y(n_185) );
NAND2xp33_ASAP7_75t_L g254 ( .A(n_98), .B(n_181), .Y(n_254) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_111), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_103), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND3x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .C(n_109), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR3x1_ASAP7_75t_L g821 ( .A(n_107), .B(n_794), .C(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g482 ( .A(n_108), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_109), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_L g813 ( .A(n_110), .B(n_794), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_787), .B(n_795), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AO22x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_479), .B1(n_480), .B2(n_483), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
NOR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_393), .Y(n_116) );
NAND4xp75_ASAP7_75t_L g117 ( .A(n_118), .B(n_298), .C(n_340), .D(n_364), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI211xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_187), .B(n_235), .C(n_277), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g384 ( .A(n_122), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g478 ( .A(n_122), .B(n_415), .Y(n_478) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_148), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g293 ( .A(n_124), .B(n_245), .Y(n_293) );
AND2x2_ASAP7_75t_L g334 ( .A(n_124), .B(n_295), .Y(n_334) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g241 ( .A(n_125), .B(n_170), .Y(n_241) );
OR2x2_ASAP7_75t_L g259 ( .A(n_125), .B(n_170), .Y(n_259) );
INVx2_ASAP7_75t_L g285 ( .A(n_125), .Y(n_285) );
AND2x2_ASAP7_75t_L g315 ( .A(n_125), .B(n_245), .Y(n_315) );
AND2x2_ASAP7_75t_L g344 ( .A(n_125), .B(n_169), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_125), .B(n_296), .Y(n_380) );
AO31x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_138), .A3(n_142), .B(n_145), .Y(n_125) );
OAI22x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B1(n_134), .B2(n_136), .Y(n_126) );
INVx4_ASAP7_75t_L g130 ( .A(n_128), .Y(n_130) );
INVx1_ASAP7_75t_L g505 ( .A(n_128), .Y(n_505) );
INVx1_ASAP7_75t_L g556 ( .A(n_128), .Y(n_556) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
INVx1_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_129), .Y(n_200) );
INVx2_ASAP7_75t_L g207 ( .A(n_129), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_130), .A2(n_249), .B(n_250), .C(n_251), .Y(n_248) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_130), .A2(n_132), .B(n_517), .C(n_518), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_131), .A2(n_152), .B1(n_215), .B2(n_216), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_131), .A2(n_136), .B1(n_268), .B2(n_270), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_131), .A2(n_136), .B1(n_493), .B2(n_495), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_131), .A2(n_503), .B1(n_506), .B2(n_507), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_131), .A2(n_520), .B(n_522), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_131), .A2(n_528), .B1(n_529), .B2(n_530), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_131), .A2(n_507), .B1(n_539), .B2(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_131), .A2(n_529), .B1(n_548), .B2(n_549), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_131), .A2(n_529), .B1(n_555), .B2(n_557), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_131), .A2(n_529), .B1(n_571), .B2(n_572), .Y(n_570) );
INVx6_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_132), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_132), .A2(n_254), .B(n_255), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_132), .A2(n_151), .B(n_161), .C(n_167), .Y(n_297) );
BUFx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_133), .Y(n_137) );
INVx2_ASAP7_75t_L g154 ( .A(n_133), .Y(n_154) );
INVx1_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_135), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g271 ( .A(n_135), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_136), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_SL g507 ( .A(n_137), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_138), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_138), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
OAI21xp33_ASAP7_75t_L g167 ( .A1(n_139), .A2(n_159), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
INVx2_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
AO31x2_ASAP7_75t_L g526 ( .A1(n_142), .A2(n_217), .A3(n_527), .B(n_531), .Y(n_526) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_142), .A2(n_193), .A3(n_538), .B(n_542), .Y(n_537) );
AO31x2_ASAP7_75t_L g546 ( .A1(n_142), .A2(n_491), .A3(n_547), .B(n_551), .Y(n_546) );
BUFx10_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
BUFx10_ASAP7_75t_L g218 ( .A(n_143), .Y(n_218) );
INVx1_ASAP7_75t_L g274 ( .A(n_143), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx2_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
BUFx2_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_147), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_147), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g357 ( .A(n_148), .B(n_286), .Y(n_357) );
INVx2_ASAP7_75t_L g452 ( .A(n_148), .Y(n_452) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_169), .Y(n_148) );
INVx2_ASAP7_75t_L g240 ( .A(n_149), .Y(n_240) );
AND2x4_ASAP7_75t_L g283 ( .A(n_149), .B(n_170), .Y(n_283) );
AOI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_160), .B(n_166), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_159), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_152), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g529 ( .A(n_153), .Y(n_529) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g252 ( .A(n_154), .Y(n_252) );
INVx1_ASAP7_75t_L g540 ( .A(n_157), .Y(n_540) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_158), .B(n_177), .Y(n_176) );
INVxp67_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g504 ( .A(n_163), .Y(n_504) );
OAI21xp33_ASAP7_75t_SL g226 ( .A1(n_164), .A2(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_195), .B(n_204), .Y(n_194) );
AND2x2_ASAP7_75t_L g442 ( .A(n_169), .B(n_240), .Y(n_442) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g306 ( .A(n_170), .Y(n_306) );
AND2x2_ASAP7_75t_L g363 ( .A(n_170), .B(n_245), .Y(n_363) );
AND2x2_ASAP7_75t_L g378 ( .A(n_170), .B(n_286), .Y(n_378) );
AND2x2_ASAP7_75t_L g400 ( .A(n_170), .B(n_240), .Y(n_400) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_185), .Y(n_170) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_171), .A2(n_273), .A3(n_554), .B(n_558), .Y(n_553) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_171), .A2(n_508), .A3(n_570), .B(n_573), .Y(n_569) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_173), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_SL g542 ( .A(n_173), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_184), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_179) );
INVx2_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
INVx1_ASAP7_75t_L g521 ( .A(n_181), .Y(n_521) );
INVx1_ASAP7_75t_L g550 ( .A(n_182), .Y(n_550) );
INVx1_ASAP7_75t_L g508 ( .A(n_184), .Y(n_508) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_187), .A2(n_448), .B(n_450), .C(n_457), .Y(n_447) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_221), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g434 ( .A(n_190), .B(n_370), .Y(n_434) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_211), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_191), .B(n_223), .Y(n_333) );
INVxp67_ASAP7_75t_L g347 ( .A(n_191), .Y(n_347) );
AND2x2_ASAP7_75t_L g367 ( .A(n_191), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_191), .B(n_280), .Y(n_374) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g263 ( .A(n_192), .Y(n_263) );
AOI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_208), .Y(n_192) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_193), .A2(n_267), .A3(n_273), .B(n_275), .Y(n_266) );
AO31x2_ASAP7_75t_L g501 ( .A1(n_193), .A2(n_502), .A3(n_508), .B(n_509), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B(n_202), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g272 ( .A(n_200), .Y(n_272) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_203), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
INVx2_ASAP7_75t_SL g494 ( .A(n_207), .Y(n_494) );
INVx2_ASAP7_75t_L g217 ( .A(n_209), .Y(n_217) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_209), .B(n_257), .Y(n_256) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g234 ( .A(n_210), .B(n_218), .Y(n_234) );
BUFx3_ASAP7_75t_L g491 ( .A(n_210), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_210), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g514 ( .A(n_210), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_210), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_210), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g308 ( .A(n_211), .B(n_290), .Y(n_308) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g356 ( .A(n_212), .B(n_263), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_212), .B(n_266), .Y(n_362) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g262 ( .A(n_213), .B(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g331 ( .A(n_213), .B(n_266), .Y(n_331) );
BUFx2_ASAP7_75t_L g338 ( .A(n_213), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_213), .B(n_266), .Y(n_418) );
AO31x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .A3(n_218), .B(n_219), .Y(n_213) );
INVx1_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g348 ( .A(n_222), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g477 ( .A(n_222), .B(n_262), .Y(n_477) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g280 ( .A(n_223), .Y(n_280) );
AND2x2_ASAP7_75t_L g291 ( .A(n_223), .B(n_266), .Y(n_291) );
AND2x2_ASAP7_75t_L g337 ( .A(n_223), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g370 ( .A(n_223), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_223), .B(n_281), .Y(n_387) );
AND2x2_ASAP7_75t_L g426 ( .A(n_223), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_231), .B(n_234), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_242), .B(n_260), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_237), .A2(n_405), .B1(n_406), .B2(n_408), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_241), .Y(n_237) );
AND2x2_ASAP7_75t_L g402 ( .A(n_238), .B(n_293), .Y(n_402) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g466 ( .A(n_240), .B(n_286), .Y(n_466) );
AND2x2_ASAP7_75t_L g430 ( .A(n_241), .B(n_325), .Y(n_430) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_258), .Y(n_242) );
OR2x2_ASAP7_75t_L g327 ( .A(n_243), .B(n_304), .Y(n_327) );
OR2x2_ASAP7_75t_L g439 ( .A(n_243), .B(n_259), .Y(n_439) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g302 ( .A(n_244), .Y(n_302) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g286 ( .A(n_245), .Y(n_286) );
BUFx3_ASAP7_75t_L g368 ( .A(n_245), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_253), .B(n_256), .Y(n_247) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g436 ( .A(n_259), .B(n_295), .Y(n_436) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g278 ( .A(n_262), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g319 ( .A(n_262), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g456 ( .A(n_262), .Y(n_456) );
INVx1_ASAP7_75t_L g475 ( .A(n_262), .Y(n_475) );
INVx2_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_263), .B(n_266), .Y(n_339) );
INVx1_ASAP7_75t_L g403 ( .A(n_264), .Y(n_403) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g464 ( .A(n_265), .Y(n_464) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g281 ( .A(n_266), .Y(n_281) );
INVx1_ASAP7_75t_L g371 ( .A(n_266), .Y(n_371) );
AO31x2_ASAP7_75t_L g490 ( .A1(n_273), .A2(n_491), .A3(n_492), .B(n_496), .Y(n_490) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_SL g523 ( .A(n_274), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B1(n_287), .B2(n_292), .Y(n_277) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g322 ( .A(n_280), .B(n_307), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_280), .B(n_290), .Y(n_382) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx3_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_283), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g407 ( .A(n_283), .B(n_391), .Y(n_407) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_284), .A2(n_322), .B1(n_323), .B2(n_328), .C1(n_334), .C2(n_335), .Y(n_321) );
OAI21xp33_ASAP7_75t_SL g351 ( .A1(n_284), .A2(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g375 ( .A(n_284), .B(n_294), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_284), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OR2x2_ASAP7_75t_L g304 ( .A(n_285), .B(n_296), .Y(n_304) );
INVx1_ASAP7_75t_L g392 ( .A(n_285), .Y(n_392) );
BUFx2_ASAP7_75t_L g326 ( .A(n_286), .Y(n_326) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_289), .B(n_330), .Y(n_359) );
OR2x2_ASAP7_75t_L g471 ( .A(n_289), .B(n_331), .Y(n_471) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g354 ( .A(n_291), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g469 ( .A(n_291), .Y(n_469) );
OAI31xp33_ASAP7_75t_L g450 ( .A1(n_292), .A2(n_451), .A3(n_453), .B(n_454), .Y(n_450) );
AND2x4_ASAP7_75t_SL g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_293), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_321), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_307), .B(n_309), .Y(n_299) );
NOR2x1_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x6_ASAP7_75t_L g420 ( .A(n_302), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g443 ( .A(n_306), .B(n_380), .Y(n_443) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_308), .A2(n_397), .B1(n_399), .B2(n_401), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_308), .A2(n_369), .B(n_431), .C(n_458), .Y(n_457) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B(n_318), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_313), .B(n_411), .C(n_412), .D(n_414), .Y(n_410) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_315), .B(n_317), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_315), .B(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g389 ( .A(n_320), .B(n_349), .Y(n_389) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_327), .A2(n_471), .B1(n_472), .B2(n_474), .Y(n_470) );
AOI221x1_ASAP7_75t_L g409 ( .A1(n_328), .A2(n_410), .B1(n_416), .B2(n_419), .C(n_422), .Y(n_409) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g361 ( .A(n_333), .B(n_362), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_334), .B(n_415), .Y(n_424) );
O2A1O1Ixp5_ASAP7_75t_L g437 ( .A1(n_335), .A2(n_419), .B(n_438), .C(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx2_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_350), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_342), .A2(n_360), .B1(n_430), .B2(n_431), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g366 ( .A(n_344), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_344), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g465 ( .A(n_344), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_347), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g468 ( .A(n_347), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_357), .B2(n_358), .C1(n_360), .C2(n_363), .Y(n_350) );
INVx1_ASAP7_75t_L g435 ( .A(n_354), .Y(n_435) );
INVx1_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g432 ( .A(n_356), .Y(n_432) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g373 ( .A(n_362), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_383), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B1(n_372), .B2(n_375), .C1(n_376), .C2(n_381), .Y(n_365) );
INVx3_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
BUFx2_ASAP7_75t_L g473 ( .A(n_368), .Y(n_473) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g445 ( .A(n_370), .Y(n_445) );
OR2x2_ASAP7_75t_L g455 ( .A(n_370), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_SL g413 ( .A(n_378), .Y(n_413) );
AND2x2_ASAP7_75t_L g458 ( .A(n_379), .B(n_415), .Y(n_458) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_418), .Y(n_417) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g474 ( .A(n_387), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g405 ( .A(n_389), .Y(n_405) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g412 ( .A(n_392), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g462 ( .A(n_392), .Y(n_462) );
NAND4xp75_ASAP7_75t_L g393 ( .A(n_394), .B(n_428), .C(n_446), .D(n_459), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_409), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_403), .B(n_404), .Y(n_395) );
INVxp33_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_398), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
AND2x2_ASAP7_75t_L g461 ( .A(n_400), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g431 ( .A(n_403), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g449 ( .A(n_414), .Y(n_449) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_SL g440 ( .A1(n_417), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_440) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_437), .Y(n_428) );
AOI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_476), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B1(n_465), .B2(n_467), .C(n_470), .Y(n_460) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx12f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g812 ( .A(n_482), .B(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_483), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_483), .Y(n_805) );
NAND4xp75_ASAP7_75t_L g483 ( .A(n_484), .B(n_626), .C(n_702), .D(n_754), .Y(n_483) );
AND3x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_599), .C(n_612), .Y(n_484) );
AOI221x1_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_533), .B1(n_560), .B2(n_564), .C(n_576), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_486), .A2(n_600), .B(n_602), .C(n_603), .Y(n_599) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g563 ( .A(n_490), .Y(n_563) );
BUFx2_ASAP7_75t_L g581 ( .A(n_490), .Y(n_581) );
OR2x2_ASAP7_75t_L g623 ( .A(n_490), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_490), .B(n_501), .Y(n_630) );
AND2x4_ASAP7_75t_L g665 ( .A(n_490), .B(n_500), .Y(n_665) );
OR2x2_ASAP7_75t_L g708 ( .A(n_490), .B(n_526), .Y(n_708) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_500), .B(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_500), .Y(n_595) );
INVx2_ASAP7_75t_L g622 ( .A(n_500), .Y(n_622) );
INVx3_ASAP7_75t_L g635 ( .A(n_500), .Y(n_635) );
AND2x2_ASAP7_75t_L g753 ( .A(n_500), .B(n_582), .Y(n_753) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g562 ( .A(n_501), .B(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g618 ( .A(n_501), .Y(n_618) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
INVx1_ASAP7_75t_L g765 ( .A(n_512), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .Y(n_512) );
AND2x2_ASAP7_75t_L g561 ( .A(n_513), .B(n_526), .Y(n_561) );
INVx1_ASAP7_75t_L g624 ( .A(n_513), .Y(n_624) );
OAI21x1_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_524), .Y(n_513) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_514), .A2(n_515), .B(n_524), .Y(n_583) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_519), .B(n_523), .Y(n_515) );
INVx2_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
AND2x2_ASAP7_75t_L g631 ( .A(n_525), .B(n_582), .Y(n_631) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g593 ( .A(n_526), .Y(n_593) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_526), .Y(n_653) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_535), .A2(n_625), .B1(n_629), .B2(n_632), .Y(n_628) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_544), .Y(n_535) );
INVx1_ASAP7_75t_L g646 ( .A(n_536), .Y(n_646) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g566 ( .A(n_537), .B(n_546), .Y(n_566) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_553), .Y(n_597) );
INVx4_ASAP7_75t_SL g608 ( .A(n_537), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_537), .B(n_642), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_537), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g679 ( .A(n_545), .B(n_657), .Y(n_679) );
OR2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_694), .Y(n_712) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_553), .Y(n_545) );
INVx2_ASAP7_75t_L g586 ( .A(n_546), .Y(n_586) );
INVx1_ASAP7_75t_L g591 ( .A(n_546), .Y(n_591) );
AND2x2_ASAP7_75t_L g598 ( .A(n_546), .B(n_568), .Y(n_598) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_546), .Y(n_614) );
INVx1_ASAP7_75t_L g642 ( .A(n_546), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_546), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g575 ( .A(n_553), .Y(n_575) );
AND2x4_ASAP7_75t_L g585 ( .A(n_553), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g611 ( .A(n_553), .Y(n_611) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_553), .Y(n_688) );
INVx1_ASAP7_75t_L g781 ( .A(n_553), .Y(n_781) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_561), .B(n_634), .Y(n_701) );
AND2x2_ASAP7_75t_L g714 ( .A(n_561), .B(n_630), .Y(n_714) );
AND2x2_ASAP7_75t_L g784 ( .A(n_561), .B(n_635), .Y(n_784) );
AND2x4_ASAP7_75t_L g619 ( .A(n_563), .B(n_582), .Y(n_619) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g686 ( .A(n_566), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g700 ( .A(n_566), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_566), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g602 ( .A(n_567), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_567), .B(n_640), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_567), .A2(n_697), .B(n_700), .C(n_701), .Y(n_696) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_575), .Y(n_567) );
AND2x2_ASAP7_75t_L g667 ( .A(n_568), .B(n_608), .Y(n_667) );
INVx3_ASAP7_75t_L g694 ( .A(n_568), .Y(n_694) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g589 ( .A(n_569), .Y(n_589) );
AND2x4_ASAP7_75t_L g615 ( .A(n_569), .B(n_575), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_575), .B(n_608), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_584), .B1(n_592), .B2(n_596), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g733 ( .A(n_578), .Y(n_733) );
AND2x4_ASAP7_75t_L g644 ( .A(n_579), .B(n_624), .Y(n_644) );
INVx1_ASAP7_75t_L g664 ( .A(n_579), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_581), .A2(n_637), .B1(n_647), .B2(n_649), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_581), .B(n_638), .Y(n_695) );
NAND2x1_ASAP7_75t_L g752 ( .A(n_581), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g767 ( .A(n_581), .Y(n_767) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g706 ( .A(n_583), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g625 ( .A(n_585), .B(n_607), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_585), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g666 ( .A(n_585), .B(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_585), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_585), .B(n_648), .Y(n_747) );
AND2x4_ASAP7_75t_L g770 ( .A(n_585), .B(n_698), .Y(n_770) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx3_ASAP7_75t_L g648 ( .A(n_588), .Y(n_648) );
AND2x2_ASAP7_75t_L g660 ( .A(n_588), .B(n_653), .Y(n_660) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g610 ( .A(n_589), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
INVx1_ASAP7_75t_L g601 ( .A(n_590), .Y(n_601) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g758 ( .A(n_591), .B(n_608), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g684 ( .A(n_593), .B(n_665), .Y(n_684) );
INVx2_ASAP7_75t_L g725 ( .A(n_593), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_593), .B(n_619), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_594), .B(n_644), .Y(n_774) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_597), .B(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g669 ( .A(n_597), .B(n_614), .Y(n_669) );
INVx1_ASAP7_75t_L g761 ( .A(n_597), .Y(n_761) );
AND2x2_ASAP7_75t_L g760 ( .A(n_598), .B(n_687), .Y(n_760) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_602), .A2(n_732), .B1(n_734), .B2(n_736), .Y(n_731) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g640 ( .A(n_608), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g676 ( .A(n_608), .Y(n_676) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_608), .Y(n_682) );
INVx2_ASAP7_75t_L g699 ( .A(n_608), .Y(n_699) );
OR2x2_ASAP7_75t_L g720 ( .A(n_608), .B(n_683), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_608), .B(n_678), .Y(n_730) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g697 ( .A(n_610), .B(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_610), .Y(n_751) );
INVx1_ASAP7_75t_L g678 ( .A(n_611), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B(n_620), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_615), .B(n_646), .Y(n_645) );
INVx3_ASAP7_75t_L g683 ( .A(n_615), .Y(n_683) );
AND2x2_ASAP7_75t_L g757 ( .A(n_615), .B(n_758), .Y(n_757) );
AOI211x1_ASAP7_75t_SL g685 ( .A1(n_616), .A2(n_686), .B(n_689), .C(n_696), .Y(n_685) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g742 ( .A(n_618), .B(n_619), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_619), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_619), .Y(n_735) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g650 ( .A(n_622), .Y(n_650) );
NOR2x1p5_ASAP7_75t_L g707 ( .A(n_622), .B(n_708), .Y(n_707) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_623), .B(n_652), .Y(n_651) );
NOR2xp67_ASAP7_75t_SL g724 ( .A(n_623), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g785 ( .A(n_625), .B(n_693), .Y(n_785) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_670), .Y(n_626) );
NAND3xp33_ASAP7_75t_SL g627 ( .A(n_628), .B(n_636), .C(n_654), .Y(n_627) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_630), .Y(n_661) );
AND2x2_ASAP7_75t_L g668 ( .A(n_630), .B(n_664), .Y(n_668) );
AND2x4_ASAP7_75t_SL g782 ( .A(n_630), .B(n_644), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_631), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_633), .A2(n_675), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g764 ( .A(n_635), .B(n_765), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_643), .B2(n_645), .Y(n_637) );
NAND2x1_ASAP7_75t_L g713 ( .A(n_640), .B(n_693), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_640), .B(n_687), .Y(n_723) );
INVx1_ASAP7_75t_L g750 ( .A(n_640), .Y(n_750) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_643), .A2(n_769), .B(n_772), .Y(n_768) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_644), .A2(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g729 ( .A(n_648), .Y(n_729) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g673 ( .A(n_651), .Y(n_673) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_661), .B1(n_662), .B2(n_666), .C1(n_668), .C2(n_669), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_656), .A2(n_690), .B(n_695), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_657), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g771 ( .A(n_657), .Y(n_771) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_658), .Y(n_777) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g741 ( .A(n_663), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g734 ( .A(n_664), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_685), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_680), .B2(n_684), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g691 ( .A(n_677), .Y(n_691) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx4_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g719 ( .A(n_694), .B(n_711), .Y(n_719) );
OR2x2_ASAP7_75t_L g779 ( .A(n_694), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND5xp2_ASAP7_75t_L g755 ( .A(n_700), .B(n_747), .C(n_756), .D(n_759), .E(n_761), .Y(n_755) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_738), .Y(n_702) );
NAND2xp67_ASAP7_75t_SL g703 ( .A(n_704), .B(n_721), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_709), .B1(n_714), .B2(n_715), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_712), .C(n_713), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g744 ( .A(n_713), .Y(n_744) );
NAND3xp33_ASAP7_75t_SL g715 ( .A(n_716), .B(n_719), .C(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g737 ( .A(n_718), .Y(n_737) );
O2A1O1Ixp33_ASAP7_75t_SL g749 ( .A1(n_719), .A2(n_750), .B(n_751), .C(n_752), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_726), .B2(n_727), .C(n_731), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_728), .B(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g745 ( .A(n_732), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
AOI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_746), .C(n_749), .Y(n_743) );
AOI211x1_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_762), .B(n_768), .C(n_783), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2x1p5_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .B1(n_778), .B2(n_782), .Y(n_772) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
BUFx12f_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x6_ASAP7_75t_SL g789 ( .A(n_790), .B(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx3_ASAP7_75t_L g798 ( .A(n_791), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_791), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_799), .B(n_806), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
BUFx8_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B(n_804), .Y(n_799) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx10_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx12f_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_816), .Y(n_825) );
AND2x6_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVxp33_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
endmodule