module fake_jpeg_25546_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_64),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_22),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_31),
.B1(n_18),
.B2(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_23),
.Y(n_85)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_69),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_79),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_40),
.B1(n_42),
.B2(n_27),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_67),
.B1(n_55),
.B2(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_27),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_23),
.B(n_21),
.C(n_34),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_59),
.B1(n_18),
.B2(n_34),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_85),
.Y(n_114)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_94),
.Y(n_120)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_49),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_96),
.B(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_60),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_72),
.B(n_91),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_115),
.B1(n_83),
.B2(n_101),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_118),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_91),
.B1(n_89),
.B2(n_74),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_47),
.B1(n_63),
.B2(n_53),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_65),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_123),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_72),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_128),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_110),
.C(n_119),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_18),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_96),
.B(n_21),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_77),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_77),
.B1(n_79),
.B2(n_76),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_90),
.B1(n_109),
.B2(n_124),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_76),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_93),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_150),
.B1(n_112),
.B2(n_100),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_144),
.Y(n_162)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_87),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_123),
.B1(n_102),
.B2(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_152),
.B1(n_90),
.B2(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_92),
.B1(n_73),
.B2(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_31),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_99),
.B1(n_106),
.B2(n_108),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_25),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_33),
.C(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_155),
.A2(n_170),
.B(n_127),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_92),
.C(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_179),
.C(n_158),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_16),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_157),
.A2(n_159),
.B(n_145),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_122),
.B(n_34),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_179),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_181),
.B1(n_182),
.B2(n_142),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_167),
.B1(n_174),
.B2(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_112),
.B1(n_57),
.B2(n_86),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_169),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_150),
.B1(n_128),
.B2(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_57),
.B1(n_21),
.B2(n_32),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_31),
.B1(n_32),
.B2(n_65),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_60),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_65),
.B1(n_25),
.B2(n_17),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_25),
.B1(n_27),
.B2(n_24),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_144),
.B1(n_163),
.B2(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_143),
.Y(n_203)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_206),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_192),
.B(n_15),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_196),
.B1(n_155),
.B2(n_185),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_132),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_131),
.B1(n_150),
.B2(n_136),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_214),
.B1(n_181),
.B2(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_141),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_211),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_171),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_15),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_164),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_183),
.B1(n_185),
.B2(n_156),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_226),
.B1(n_238),
.B2(n_214),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_213),
.B1(n_198),
.B2(n_193),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_157),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_173),
.C(n_171),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_216),
.C(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_173),
.B1(n_9),
.B2(n_10),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_12),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_261),
.B1(n_262),
.B2(n_218),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_250),
.B1(n_224),
.B2(n_218),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_194),
.B1(n_206),
.B2(n_191),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_228),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_217),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_258),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_190),
.C(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.C(n_263),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_212),
.C(n_202),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_220),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_10),
.C(n_1),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_239),
.C(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_256),
.C(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_241),
.C(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_277),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_250),
.B1(n_243),
.B2(n_255),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_253),
.B1(n_265),
.B2(n_274),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_237),
.B(n_233),
.C(n_227),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_251),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_277),
.B1(n_275),
.B2(n_2),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_260),
.C(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_292),
.C(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_236),
.B1(n_219),
.B2(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_0),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_6),
.C(n_1),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_0),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_0),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_270),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_300),
.C(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_285),
.A2(n_0),
.B(n_1),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_292),
.B(n_4),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_2),
.C(n_3),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_3),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_4),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_282),
.C(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_301),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_305),
.B(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_300),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_311),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_323),
.B(n_317),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_293),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_307),
.B(n_321),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_310),
.B(n_315),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_318),
.C(n_323),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_298),
.B(n_5),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_5),
.Y(n_329)
);


endmodule