module fake_netlist_5_332_n_7877 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_256, n_305, n_533, n_52, n_278, n_110, n_7877);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_7877;

wire n_924;
wire n_6643;
wire n_6122;
wire n_2253;
wire n_977;
wire n_2756;
wire n_2417;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_7164;
wire n_5287;
wire n_6546;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_7710;
wire n_5035;
wire n_2391;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_7461;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_6649;
wire n_7154;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_6810;
wire n_7660;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_7686;
wire n_4211;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_6742;
wire n_3019;
wire n_2096;
wire n_6694;
wire n_877;
wire n_3776;
wire n_7616;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_6913;
wire n_7867;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_4131;
wire n_7772;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_7641;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_1242;
wire n_7468;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_7861;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_5648;
wire n_7667;
wire n_1314;
wire n_1512;
wire n_6931;
wire n_1490;
wire n_6618;
wire n_6408;
wire n_3214;
wire n_7523;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_1449;
wire n_6698;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_6214;
wire n_7493;
wire n_3868;
wire n_1948;
wire n_3183;
wire n_3437;
wire n_7804;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_6939;
wire n_882;
wire n_2384;
wire n_7528;
wire n_3156;
wire n_3376;
wire n_7562;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_6707;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_7402;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_901;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_7801;
wire n_1151;
wire n_1405;
wire n_7463;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_6725;
wire n_7613;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_2968;
wire n_7316;
wire n_1585;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_1000;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6062;
wire n_6191;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_5909;
wire n_1385;
wire n_7575;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_1527;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_7701;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_6793;
wire n_7873;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_7568;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_4983;
wire n_2379;
wire n_5695;
wire n_7814;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_3649;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_2514;
wire n_5862;
wire n_6304;
wire n_5189;
wire n_6956;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_1027;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_7002;
wire n_1412;
wire n_3981;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_6027;
wire n_6598;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_1711;
wire n_870;
wire n_6638;
wire n_1891;
wire n_7308;
wire n_5254;
wire n_3526;
wire n_6900;
wire n_2546;
wire n_965;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_7457;
wire n_4613;
wire n_7718;
wire n_4649;
wire n_7617;
wire n_1888;
wire n_6269;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_7768;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_6013;
wire n_7357;
wire n_2449;
wire n_5083;
wire n_6927;
wire n_1194;
wire n_6503;
wire n_5888;
wire n_2297;
wire n_4186;
wire n_7310;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_7593;
wire n_6256;
wire n_7716;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_5870;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_7076;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_6982;
wire n_1680;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_3317;
wire n_7539;
wire n_1121;
wire n_7229;
wire n_4391;
wire n_949;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_1195;
wire n_7797;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_757;
wire n_7869;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_2805;
wire n_7781;
wire n_1145;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_1153;
wire n_3856;
wire n_741;
wire n_7624;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_1163;
wire n_6805;
wire n_6185;
wire n_1207;
wire n_5010;
wire n_7762;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_940;
wire n_6351;
wire n_7552;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_6901;
wire n_2947;
wire n_978;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_6411;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_7746;
wire n_5435;
wire n_1431;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_7139;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_7857;
wire n_962;
wire n_723;
wire n_2536;
wire n_6387;
wire n_1336;
wire n_7223;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_6019;
wire n_6222;
wire n_7165;
wire n_3505;
wire n_6223;
wire n_4610;
wire n_6435;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_974;
wire n_727;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_5657;
wire n_957;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_6844;
wire n_3001;
wire n_7795;
wire n_7404;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_6295;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_3185;
wire n_1300;
wire n_6087;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_7822;
wire n_2017;
wire n_2604;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_6790;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_3984;
wire n_6807;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_7708;
wire n_1823;
wire n_7696;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_7115;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_6218;
wire n_7281;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_1552;
wire n_6189;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_815;
wire n_4594;
wire n_6153;
wire n_3424;
wire n_5970;
wire n_1381;
wire n_6418;
wire n_1037;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_3215;
wire n_2419;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_1437;
wire n_6591;
wire n_6266;
wire n_7161;
wire n_7580;
wire n_7153;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_7350;
wire n_5690;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_6967;
wire n_5885;
wire n_2254;
wire n_6433;
wire n_1382;
wire n_925;
wire n_3546;
wire n_7535;
wire n_6893;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_7632;
wire n_3244;
wire n_6501;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_6798;
wire n_5702;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_7844;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_6986;
wire n_802;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_6745;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_7594;
wire n_7766;
wire n_3715;
wire n_7803;
wire n_7340;
wire n_6699;
wire n_7747;
wire n_6073;
wire n_972;
wire n_5767;
wire n_6324;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_6138;
wire n_7603;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_6477;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_6159;
wire n_6283;
wire n_7396;
wire n_5322;
wire n_856;
wire n_7116;
wire n_1793;
wire n_4352;
wire n_7519;
wire n_4441;
wire n_6943;
wire n_918;
wire n_4761;
wire n_6827;
wire n_6173;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_6312;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_4043;
wire n_2291;
wire n_1636;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_7770;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1096;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_7664;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_6300;
wire n_7815;
wire n_2043;
wire n_2751;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_7023;
wire n_1807;
wire n_2618;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_6783;
wire n_4748;
wire n_7465;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_7847;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_7149;
wire n_2795;
wire n_6459;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_7700;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_6869;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_7117;
wire n_789;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_6555;
wire n_3877;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_6490;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_5460;
wire n_2097;
wire n_7628;
wire n_4304;
wire n_6761;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_6294;
wire n_6767;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_4805;
wire n_4885;
wire n_7838;
wire n_7786;
wire n_5983;
wire n_1661;
wire n_5804;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_861;
wire n_6582;
wire n_1658;
wire n_7752;
wire n_1904;
wire n_6996;
wire n_1345;
wire n_1899;
wire n_6974;
wire n_7731;
wire n_6765;
wire n_7577;
wire n_1003;
wire n_6921;
wire n_2067;
wire n_2219;
wire n_7845;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_7709;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_1657;
wire n_5886;
wire n_768;
wire n_7080;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_7744;
wire n_1491;
wire n_754;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_6960;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_6836;
wire n_2605;
wire n_1310;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_6972;
wire n_2924;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_5785;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_766;
wire n_6010;
wire n_7247;
wire n_1117;
wire n_6833;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_7481;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_7687;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_6265;
wire n_1650;
wire n_1137;
wire n_6821;
wire n_3934;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_7742;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_7758;
wire n_7547;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_5630;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_7513;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_7540;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_7622;
wire n_7005;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_7353;
wire n_6219;
wire n_1889;
wire n_6965;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_6720;
wire n_1569;
wire n_2188;
wire n_6032;
wire n_7174;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_756;
wire n_1429;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_7816;
wire n_3170;
wire n_7591;
wire n_5775;
wire n_2748;
wire n_3311;
wire n_7830;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_1861;
wire n_760;
wire n_5731;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_5831;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_2939;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_886;
wire n_5653;
wire n_6258;
wire n_7070;
wire n_1221;
wire n_5394;
wire n_6755;
wire n_2774;
wire n_7276;
wire n_7351;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_6084;
wire n_4827;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_7666;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_7211;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_7368;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_2526;
wire n_6389;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_6910;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_816;
wire n_5678;
wire n_5935;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6331;
wire n_1555;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_6278;
wire n_6787;
wire n_6872;
wire n_4899;
wire n_796;
wire n_6208;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_1012;
wire n_5411;
wire n_7754;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_6990;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_5185;
wire n_1193;
wire n_6359;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_7763;
wire n_1487;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_6301;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_6744;
wire n_4981;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_7381;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_7291;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_3267;
wire n_4995;
wire n_7870;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_6104;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6475;
wire n_3884;
wire n_6465;
wire n_3726;
wire n_6496;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_7305;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_1074;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_7545;
wire n_7846;
wire n_1448;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_6194;
wire n_7695;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_7537;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_7489;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_1186;
wire n_5883;
wire n_6985;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_7451;
wire n_6238;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_6366;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_7236;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_3256;
wire n_7560;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_1501;
wire n_7572;
wire n_3086;
wire n_1007;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_6529;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_7140;
wire n_7233;
wire n_819;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_5457;
wire n_7352;
wire n_951;
wire n_7134;
wire n_5532;
wire n_1494;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_6525;
wire n_7650;
wire n_3434;
wire n_1806;
wire n_933;
wire n_6631;
wire n_6892;
wire n_1563;
wire n_7663;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_7729;
wire n_3987;
wire n_7339;
wire n_902;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_6658;
wire n_6264;
wire n_6925;
wire n_5919;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_7767;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_7672;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_7482;
wire n_6864;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_6494;
wire n_5503;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_6199;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_3022;
wire n_7839;
wire n_4264;
wire n_7504;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_7360;
wire n_7681;
wire n_7301;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_7794;
wire n_7366;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_6947;
wire n_1723;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_7309;
wire n_4626;
wire n_1097;
wire n_1036;
wire n_6863;
wire n_6637;
wire n_798;
wire n_6100;
wire n_7860;
wire n_6735;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_6358;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_7876;
wire n_6050;
wire n_2470;
wire n_7244;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_7610;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_5903;
wire n_6371;
wire n_813;
wire n_1284;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_7751;
wire n_6510;
wire n_1748;
wire n_4569;
wire n_6468;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_7788;
wire n_1064;
wire n_5842;
wire n_858;
wire n_6352;
wire n_2985;
wire n_5722;
wire n_7534;
wire n_5636;
wire n_7719;
wire n_5065;
wire n_2753;
wire n_7287;
wire n_1582;
wire n_7032;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_7851;
wire n_1211;
wire n_6332;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_5877;
wire n_907;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_6751;
wire n_7068;
wire n_892;
wire n_4556;
wire n_6322;
wire n_5454;
wire n_7704;
wire n_2620;
wire n_7773;
wire n_6667;
wire n_7526;
wire n_1581;
wire n_6530;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_6405;
wire n_6613;
wire n_4353;
wire n_2042;
wire n_6248;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_7821;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_6894;
wire n_1856;
wire n_7267;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_7387;
wire n_7431;
wire n_7654;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_847;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_822;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_6140;
wire n_1779;
wire n_7441;
wire n_4738;
wire n_6211;
wire n_1369;
wire n_3909;
wire n_6307;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_809;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_5697;
wire n_7188;
wire n_1810;
wire n_7573;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_6515;
wire n_6011;
wire n_7722;
wire n_6645;
wire n_3150;
wire n_747;
wire n_6984;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_7193;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_2181;
wire n_1829;
wire n_6183;
wire n_7522;
wire n_5882;
wire n_4030;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_1710;
wire n_7502;
wire n_1128;
wire n_2928;
wire n_7335;
wire n_7103;
wire n_1734;
wire n_4820;
wire n_6246;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_6383;
wire n_4938;
wire n_7020;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_7825;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_7533;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_3667;
wire n_1987;
wire n_878;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_6611;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_6116;
wire n_919;
wire n_7186;
wire n_4356;
wire n_6819;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_6473;
wire n_1586;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_6310;
wire n_7840;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_7658;
wire n_7828;
wire n_4935;
wire n_6365;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_7401;
wire n_6828;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_6355;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_7835;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_7356;
wire n_1721;
wire n_2338;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_6754;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_7585;
wire n_4570;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_2418;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_7544;
wire n_3458;
wire n_5712;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_7255;
wire n_4093;
wire n_1486;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_6237;
wire n_834;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_893;
wire n_6341;
wire n_1965;
wire n_1902;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_6697;
wire n_874;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_3189;
wire n_2066;
wire n_6449;
wire n_993;
wire n_7832;
wire n_3154;
wire n_1551;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_7584;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_6983;
wire n_970;
wire n_7843;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_7222;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_3486;
wire n_6808;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_6571;
wire n_921;
wire n_5100;
wire n_7470;
wire n_1795;
wire n_5849;
wire n_6251;
wire n_7400;
wire n_2578;
wire n_3483;
wire n_6635;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_7623;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_5034;
wire n_6733;
wire n_1708;
wire n_7071;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_7859;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_1776;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_5754;
wire n_6016;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_7212;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_6726;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_967;
wire n_6689;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_7777;
wire n_2998;
wire n_6277;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_6095;
wire n_7671;
wire n_6247;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_6616;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_7871;
wire n_6946;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_1228;
wire n_6317;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_7649;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_945;
wire n_6693;
wire n_3743;
wire n_6734;
wire n_7135;
wire n_7014;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_984;
wire n_6382;
wire n_7328;
wire n_1983;
wire n_7635;
wire n_6404;
wire n_5975;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_6379;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_1977;
wire n_1147;
wire n_2153;
wire n_6235;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_6417;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_7728;
wire n_3442;
wire n_1201;
wire n_7690;
wire n_1114;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_7270;
wire n_1176;
wire n_5940;
wire n_1149;
wire n_7390;
wire n_1020;
wire n_7805;
wire n_7807;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_6914;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_6272;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_6236;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_849;
wire n_6871;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_7506;
wire n_2340;
wire n_3552;
wire n_875;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_5578;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_969;
wire n_1401;
wire n_4113;
wire n_1998;
wire n_1019;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_6992;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7304;
wire n_5792;
wire n_1187;
wire n_6657;
wire n_7756;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_1174;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_7612;
wire n_6113;
wire n_7789;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_6242;
wire n_7088;
wire n_6519;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_6842;
wire n_7588;
wire n_3390;
wire n_1573;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_6801;
wire n_774;
wire n_2493;
wire n_4930;
wire n_7680;
wire n_5276;
wire n_6308;
wire n_1059;
wire n_7398;
wire n_1133;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_2885;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_4282;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_6415;
wire n_2994;
wire n_6857;
wire n_3135;
wire n_2401;
wire n_5476;
wire n_7842;
wire n_2003;
wire n_5856;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_6361;
wire n_3438;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_872;
wire n_5684;
wire n_5861;
wire n_1297;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_7862;
wire n_2806;
wire n_1184;
wire n_5312;
wire n_2184;
wire n_985;
wire n_5850;
wire n_3404;
wire n_3217;
wire n_3425;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7820;
wire n_7167;
wire n_7833;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_7643;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_6712;
wire n_1602;
wire n_1178;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_6953;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_780;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_5674;
wire n_3600;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_1388;
wire n_2836;
wire n_5682;
wire n_6392;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_5612;
wire n_6125;
wire n_6599;
wire n_6685;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_6560;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_5301;
wire n_7800;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_7615;
wire n_5898;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1024;
wire n_7298;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_7581;
wire n_4049;
wire n_6641;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_1238;
wire n_7190;
wire n_7112;
wire n_7678;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_6195;
wire n_862;
wire n_3584;
wire n_6356;
wire n_3756;
wire n_2889;
wire n_7001;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_7829;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_6559;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_6653;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_786;
wire n_1142;
wire n_2579;
wire n_6923;
wire n_6825;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_6399;
wire n_1873;
wire n_3201;
wire n_6275;
wire n_1087;
wire n_5666;
wire n_6575;
wire n_3472;
wire n_7732;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_1247;
wire n_7459;
wire n_7096;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_7551;
wire n_4045;
wire n_6678;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_7750;
wire n_5015;
wire n_2702;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_6752;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_2209;
wire n_7652;
wire n_7808;
wire n_6500;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_7051;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_6628;
wire n_844;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_1601;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_5688;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_6293;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2505;
wire n_2427;
wire n_7676;
wire n_4061;
wire n_3250;
wire n_2070;
wire n_7553;
wire n_6905;
wire n_7425;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_1379;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_6577;
wire n_6899;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_6370;
wire n_3266;
wire n_7210;
wire n_4646;
wire n_5769;
wire n_6065;
wire n_1130;
wire n_7039;
wire n_6987;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_6190;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_6309;
wire n_6623;
wire n_7723;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_7811;
wire n_5341;
wire n_4320;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_7348;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_3688;
wire n_6865;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_6535;
wire n_904;
wire n_3338;
wire n_7213;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_5966;
wire n_1542;
wire n_7456;
wire n_5041;
wire n_7420;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_6482;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_7715;
wire n_1780;
wire n_3732;
wire n_6605;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_5908;
wire n_6018;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_7736;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_7177;
wire n_5939;
wire n_3766;
wire n_1353;
wire n_800;
wire n_7780;
wire n_2880;
wire n_7379;
wire n_3350;
wire n_4165;
wire n_2389;
wire n_1666;
wire n_4866;
wire n_7444;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_7813;
wire n_864;
wire n_7030;
wire n_5420;
wire n_1264;
wire n_6311;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_1607;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_5679;
wire n_947;
wire n_3710;
wire n_5938;
wire n_6702;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_1230;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_6452;
wire n_929;
wire n_3379;
wire n_4374;
wire n_6791;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_7280;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_6915;
wire n_7110;
wire n_1104;
wire n_1294;
wire n_7511;
wire n_1257;
wire n_6856;
wire n_1182;
wire n_7791;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_7232;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_6364;
wire n_6451;
wire n_6552;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_4816;
wire n_7827;
wire n_1483;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_6978;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_1374;
wire n_4793;
wire n_7363;
wire n_6612;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_955;
wire n_5511;
wire n_7863;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_7295;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_897;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_1428;
wire n_6866;
wire n_7831;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_7466;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_1513;
wire n_2970;
wire n_7651;
wire n_2235;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_6935;
wire n_1590;
wire n_7530;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6907;
wire n_6158;
wire n_7661;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_6338;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_7823;
wire n_7467;
wire n_736;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_7541;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_7241;
wire n_7717;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_7464;
wire n_2590;
wire n_6302;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_6706;
wire n_944;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_7434;
wire n_7636;
wire n_7054;
wire n_6999;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_6228;
wire n_857;
wire n_5650;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_4702;
wire n_6888;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_971;
wire n_6800;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_6922;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_7503;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7273;
wire n_6647;
wire n_7296;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_7543;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_7507;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_7555;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_914;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_759;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_7033;
wire n_6121;
wire n_1571;
wire n_3119;
wire n_7531;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_6646;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_7131;
wire n_7769;
wire n_6903;
wire n_1647;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_6941;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_6106;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_7688;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_7806;
wire n_6566;
wire n_1443;
wire n_946;
wire n_1539;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_7204;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_6047;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_7354;
wire n_7448;
wire n_6244;
wire n_2290;
wire n_6861;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_7852;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_5163;
wire n_2039;
wire n_7748;
wire n_5768;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_6588;
wire n_3396;
wire n_1445;
wire n_7050;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_7136;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_6108;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_6165;
wire n_1828;
wire n_6621;
wire n_2320;
wire n_1045;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_7810;
wire n_4640;
wire n_2583;
wire n_6323;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_7817;
wire n_2523;
wire n_6933;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_1578;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_3719;
wire n_7855;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_7764;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_6216;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_7263;
wire n_743;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_6911;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_6327;
wire n_2595;
wire n_761;
wire n_6607;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_7240;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_7725;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_1015;
wire n_7278;
wire n_1651;
wire n_7630;
wire n_2775;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_6695;
wire n_3557;
wire n_2230;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_1455;
wire n_6600;
wire n_767;
wire n_2490;
wire n_1407;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_5969;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_6458;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_6746;
wire n_2508;
wire n_4031;
wire n_7586;
wire n_7720;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_2461;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_6851;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_1082;
wire n_3961;
wire n_716;
wire n_1630;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_7841;
wire n_6619;
wire n_1023;
wire n_5603;
wire n_6804;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_1056;
wire n_3588;
wire n_7792;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_7809;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3298;
wire n_3033;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_2333;
wire n_2916;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_7569;
wire n_7003;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_7419;
wire n_5827;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_7784;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_7500;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_7864;
wire n_5228;
wire n_1504;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_7790;
wire n_3572;
wire n_992;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_842;
wire n_7642;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_7045;
wire n_1643;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3078;
wire n_6979;
wire n_6203;
wire n_7405;
wire n_7739;
wire n_894;
wire n_3253;
wire n_7207;
wire n_4027;
wire n_831;
wire n_2280;
wire n_7454;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_6870;
wire n_7639;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_7251;
wire n_2303;
wire n_7776;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_830;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_1655;
wire n_749;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_7782;
wire n_7220;
wire n_717;
wire n_4316;
wire n_3697;
wire n_939;
wire n_7438;
wire n_1232;
wire n_734;
wire n_2638;
wire n_7515;
wire n_7574;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_7065;
wire n_1338;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_1522;
wire n_7868;
wire n_6973;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_5200;
wire n_1653;
wire n_5659;
wire n_1506;
wire n_5618;
wire n_6325;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_7008;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_6111;
wire n_1834;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_6260;
wire n_7501;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_6665;
wire n_7566;
wire n_7055;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_726;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_7872;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_7819;
wire n_6570;
wire n_1410;
wire n_707;
wire n_6498;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_6692;
wire n_937;
wire n_6074;
wire n_2779;
wire n_7561;
wire n_1584;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_6045;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_2811;
wire n_3348;
wire n_7415;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_895;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_6772;
wire n_1991;
wire n_2224;
wire n_1543;
wire n_6823;
wire n_6877;
wire n_732;
wire n_6806;
wire n_7426;
wire n_5906;
wire n_4743;
wire n_3805;
wire n_1067;
wire n_3825;
wire n_6831;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_7217;
wire n_2692;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_799;
wire n_6785;
wire n_1213;
wire n_6374;
wire n_6930;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_7735;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_6838;
wire n_869;
wire n_5736;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_1352;
wire n_2197;
wire n_7558;
wire n_2199;
wire n_5069;
wire n_7442;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_2480;
wire n_6034;
wire n_7499;
wire n_2363;
wire n_4072;
wire n_916;
wire n_5579;
wire n_1115;
wire n_7085;
wire n_4781;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_4424;
wire n_823;
wire n_725;
wire n_7611;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_719;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_1683;
wire n_1530;
wire n_997;
wire n_7627;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_5793;
wire n_5591;
wire n_7856;
wire n_1320;
wire n_4050;
wire n_7496;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_5623;
wire n_1063;
wire n_5681;
wire n_4853;
wire n_981;
wire n_7399;
wire n_867;
wire n_2422;
wire n_6213;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_7605;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_905;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_782;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_6858;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_1330;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_7837;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_6430;
wire n_6193;
wire n_934;
wire n_5314;
wire n_6462;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_787;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_7812;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_5777;
wire n_2764;
wire n_1498;
wire n_7046;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_7579;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_928;
wire n_1943;
wire n_7460;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_7698;
wire n_6154;
wire n_7344;
wire n_1396;
wire n_1348;
wire n_6020;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_7079;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_7774;
wire n_5797;
wire n_6696;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_6210;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_6964;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_6681;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_6661;
wire n_3303;
wire n_1654;
wire n_6640;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_3591;
wire n_2196;
wire n_7721;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_6832;
wire n_7836;
wire n_1595;
wire n_2161;
wire n_6160;
wire n_7564;
wire n_2404;
wire n_2083;
wire n_6718;
wire n_2503;
wire n_6542;
wire n_1540;
wire n_1936;
wire n_6031;
wire n_5568;
wire n_2027;
wire n_5502;
wire n_2642;
wire n_720;
wire n_2500;
wire n_7653;
wire n_1918;
wire n_5656;
wire n_863;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_3480;
wire n_2695;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_2414;
wire n_6438;
wire n_1402;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_6758;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_6874;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_6030;
wire n_6077;
wire n_4119;
wire n_3799;
wire n_7743;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_4474;
wire n_1089;
wire n_6386;
wire n_5217;
wire n_1004;
wire n_5957;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7737;
wire n_7433;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_7347;
wire n_4580;
wire n_6792;
wire n_7633;
wire n_1263;
wire n_6177;
wire n_5912;
wire n_1126;
wire n_7798;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_5396;
wire n_7693;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_6557;
wire n_7300;
wire n_956;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_7532;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_1545;
wire n_2374;
wire n_5859;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_1152;
wire n_7118;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6285;
wire n_6778;
wire n_6025;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_7669;
wire n_5268;
wire n_6318;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_6315;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_6343;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_920;
wire n_2515;
wire n_7865;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_6912;
wire n_5914;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_7133;
wire n_1850;
wire n_6883;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_7518;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_1547;
wire n_777;
wire n_6407;
wire n_1755;
wire n_6749;
wire n_6839;
wire n_7711;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_7705;
wire n_2915;
wire n_1239;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_1521;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_7854;
wire n_2337;
wire n_7707;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_6736;
wire n_5344;
wire n_923;
wire n_6526;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_6350;
wire n_7013;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_7656;
wire n_3885;
wire n_6845;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_6508;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_7570;
wire n_7771;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_5626;
wire n_6603;
wire n_6114;
wire n_1463;
wire n_6576;
wire n_3651;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_7714;
wire n_4815;
wire n_7202;
wire n_4246;
wire n_3580;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_7621;
wire n_5291;
wire n_5876;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_1565;
wire n_4088;
wire n_6876;
wire n_7778;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_7028;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_7320;
wire n_6255;
wire n_7313;
wire n_7343;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_7875;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_7337;
wire n_6989;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_7753;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_887;
wire n_6270;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_6239;
wire n_4553;
wire n_746;
wire n_6803;
wire n_784;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_7657;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_5867;
wire n_6048;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_6773;
wire n_3833;
wire n_5632;
wire n_865;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_6336;
wire n_2022;
wire n_3814;
wire n_7041;
wire n_1415;
wire n_2592;
wire n_7802;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_1191;
wire n_7557;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_6463;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_6372;
wire n_7176;
wire n_1529;
wire n_5625;
wire n_5778;
wire n_2469;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_7826;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_6254;
wire n_6161;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_908;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_7037;
wire n_4814;
wire n_724;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_959;
wire n_3031;
wire n_7258;
wire n_7432;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_6334;
wire n_1169;
wire n_3385;
wire n_2666;
wire n_6848;
wire n_2171;
wire n_4708;
wire n_6321;
wire n_7765;
wire n_2768;
wire n_2314;
wire n_6794;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_7761;
wire n_7197;
wire n_5489;
wire n_1593;
wire n_6400;
wire n_3767;
wire n_2873;
wire n_2299;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_6705;
wire n_7775;
wire n_2162;
wire n_7619;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_3607;
wire n_4925;
wire n_7548;
wire n_1921;
wire n_1309;
wire n_6534;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_6181;
wire n_3276;
wire n_1177;
wire n_6728;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_6133;
wire n_6528;
wire n_7604;
wire n_7407;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_6670;
wire n_6774;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_6038;
wire n_4818;
wire n_7727;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_2033;
wire n_1591;
wire n_7684;
wire n_7755;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_5932;
wire n_6178;
wire n_1111;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_7787;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_7849;
wire n_5186;
wire n_7367;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_7799;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_5631;
wire n_2467;
wire n_6539;
wire n_1094;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_1209;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_5326;
wire n_1435;
wire n_3394;
wire n_879;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_7738;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_7785;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_7373;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_7874;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_7760;
wire n_4248;
wire n_5915;
wire n_6818;
wire n_5452;
wire n_7226;
wire n_4754;
wire n_7057;
wire n_7685;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6815;
wire n_6753;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_7730;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_6764;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_7706;
wire n_6391;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_6471;
wire n_1844;
wire n_3777;
wire n_6627;
wire n_5761;
wire n_4784;
wire n_7203;
wire n_2999;
wire n_7512;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_7215;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_7694;
wire n_1179;
wire n_6243;
wire n_753;
wire n_6488;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_820;
wire n_1911;
wire n_3616;
wire n_4058;
wire n_2460;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_6867;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_1688;
wire n_6633;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_6574;
wire n_6395;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_7198;
wire n_1557;
wire n_4201;
wire n_6784;
wire n_6168;
wire n_896;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_7249;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_814;
wire n_2707;
wire n_6799;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_1472;
wire n_6149;
wire n_1671;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_1062;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_6450;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_1188;
wire n_6107;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_7759;
wire n_2352;
wire n_7818;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_1110;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_7447;
wire n_866;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_5899;
wire n_7629;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_7601;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_7757;
wire n_5865;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_6679;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_7625;
wire n_5822;
wire n_2564;
wire n_6259;
wire n_4947;
wire n_876;
wire n_7284;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_3450;
wire n_966;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_2217;
wire n_1453;
wire n_6630;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_6279;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_710;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_1168;
wire n_6813;
wire n_5564;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_7106;
wire n_6042;
wire n_7644;
wire n_1853;
wire n_1356;
wire n_6057;
wire n_1787;
wire n_4137;
wire n_7529;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_3972;
wire n_6207;
wire n_5539;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_3308;
wire n_6524;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_1720;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_5261;
wire n_6520;
wire n_7853;
wire n_7648;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_1782;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_1170;
wire n_6425;
wire n_2213;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_7638;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_5534;
wire n_6432;
wire n_1461;
wire n_3204;
wire n_7259;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_7237;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_6388;
wire n_5904;
wire n_4880;
wire n_6760;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_7576;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_6487;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_3647;
wire n_5755;
wire n_825;
wire n_2819;
wire n_5949;
wire n_737;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_7858;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_4535;
wire n_7668;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_792;
wire n_6843;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_7082;
wire n_3084;
wire n_6120;
wire n_1727;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_7689;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_7824;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_7796;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_7034;
wire n_6086;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_7084;
wire n_5845;
wire n_7293;
wire n_1225;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_994;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_1567;
wire n_7520;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_6267;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_1250;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_7163;
wire n_7620;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_2208;
wire n_6847;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_7563;
wire n_6298;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_7361;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_7322;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_5070;
wire n_6377;
wire n_1337;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_1321;
wire n_2296;
wire n_3181;
wire n_6348;
wire n_7713;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_1076;
wire n_1408;
wire n_1761;
wire n_5874;
wire n_730;
wire n_7508;
wire n_7021;
wire n_5270;
wire n_5956;
wire n_7834;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_6078;
wire n_7000;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_1526;
wire n_5823;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_7538;
wire n_712;
wire n_7517;
wire n_1583;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_7077;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_6942;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_6511;
wire n_3721;
wire n_1254;
wire n_6507;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_7319;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_6606;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_269),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_177),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_115),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_116),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_130),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_411),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_515),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_41),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_249),
.Y(n_715)
);

BUFx5_ASAP7_75t_L g716 ( 
.A(n_234),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_205),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_674),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_567),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_642),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_631),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_291),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_329),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_373),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_484),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_595),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_160),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_121),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_370),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_624),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_393),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_51),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_606),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_444),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_32),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_465),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_204),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_506),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_168),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_394),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_179),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_427),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_448),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_6),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_242),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_525),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_348),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_525),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_399),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_98),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_502),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_3),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_281),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_278),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_483),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_309),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_67),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_258),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_220),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_303),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_161),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_114),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_282),
.Y(n_764)
);

CKINVDCx16_ASAP7_75t_R g765 ( 
.A(n_351),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_616),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_326),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_509),
.Y(n_768)
);

BUFx8_ASAP7_75t_SL g769 ( 
.A(n_636),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_463),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_331),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_72),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_349),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_533),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_628),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_361),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_188),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_259),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_520),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_193),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_243),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_200),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_143),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_54),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_42),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_130),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_101),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_377),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_66),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_311),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_593),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_144),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_454),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_204),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_564),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_135),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_421),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_31),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_99),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_386),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_227),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_367),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_697),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_277),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_338),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_471),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_156),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_645),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_484),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_1),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_391),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_138),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_194),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_697),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_701),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_643),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_512),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_257),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_8),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_412),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_55),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_420),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_339),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_453),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_370),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_610),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_645),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_259),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_541),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_322),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_427),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_418),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_467),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_523),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_149),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_549),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_440),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_113),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_140),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_700),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_60),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_13),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_298),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_405),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_128),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_577),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_284),
.Y(n_847)
);

CKINVDCx16_ASAP7_75t_R g848 ( 
.A(n_266),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_179),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_342),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_125),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_510),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_518),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_690),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_511),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_206),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_519),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_596),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_523),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_206),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_596),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_156),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_566),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_302),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_250),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_358),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_557),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_222),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_655),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_349),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_225),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_187),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_0),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_495),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_284),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_147),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_341),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_470),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_388),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_578),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_182),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_540),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_170),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_351),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_414),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_504),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_123),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_314),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_30),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_248),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_418),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_91),
.Y(n_892)
);

BUFx5_ASAP7_75t_L g893 ( 
.A(n_545),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_236),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_331),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_374),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_637),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_287),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_268),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_8),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_701),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_623),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_136),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_243),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_373),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_568),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_542),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_456),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_49),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_183),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_49),
.Y(n_911)
);

CKINVDCx16_ASAP7_75t_R g912 ( 
.A(n_512),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_316),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_252),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_555),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_8),
.Y(n_916)
);

BUFx5_ASAP7_75t_L g917 ( 
.A(n_102),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_508),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_32),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_444),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_586),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_209),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_272),
.Y(n_923)
);

CKINVDCx16_ASAP7_75t_R g924 ( 
.A(n_111),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_393),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_235),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_676),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_41),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_547),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_681),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_475),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_401),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_565),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_111),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_225),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_37),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_452),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_391),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_375),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_25),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_384),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_321),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_650),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_371),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_224),
.Y(n_945)
);

BUFx10_ASAP7_75t_L g946 ( 
.A(n_629),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_157),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_680),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_126),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_375),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_54),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_704),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_254),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_602),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_446),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_623),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_527),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_181),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_578),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_678),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_120),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_176),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_472),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_244),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_453),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_26),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_154),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_71),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_458),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_189),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_93),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_173),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_151),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_76),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_419),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_48),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_463),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_270),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_224),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_706),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_345),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_478),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_85),
.Y(n_983)
);

BUFx10_ASAP7_75t_L g984 ( 
.A(n_226),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_136),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_348),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_434),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_593),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_146),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_627),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_612),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_120),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_506),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_233),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_477),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_328),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_374),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_538),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_503),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_430),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_640),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_272),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_86),
.Y(n_1003)
);

CKINVDCx16_ASAP7_75t_R g1004 ( 
.A(n_78),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_500),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_309),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_467),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_129),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_128),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_289),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_377),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_301),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_77),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_298),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_679),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_585),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_314),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_41),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_403),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_323),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_553),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_449),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_594),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_365),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_278),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_34),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_647),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_310),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_686),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_104),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_429),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_102),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_126),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_587),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_474),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_242),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_288),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_371),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_403),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_489),
.Y(n_1040)
);

CKINVDCx14_ASAP7_75t_R g1041 ( 
.A(n_662),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_594),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_164),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_86),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_240),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_71),
.Y(n_1046)
);

BUFx5_ASAP7_75t_L g1047 ( 
.A(n_534),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_342),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_48),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_197),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_333),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_482),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_271),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_473),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_336),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_335),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_149),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_249),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_455),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_320),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_24),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_559),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_601),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_385),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_280),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_446),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_367),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_44),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_147),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_388),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_143),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_236),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_565),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_95),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_80),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_277),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_386),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_255),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_334),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_198),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_380),
.Y(n_1081)
);

BUFx10_ASAP7_75t_L g1082 ( 
.A(n_279),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_266),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_230),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_694),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_153),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_473),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_358),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_566),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_379),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_507),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_327),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_44),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_123),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_554),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_356),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_189),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_479),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_181),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_558),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_567),
.Y(n_1101)
);

CKINVDCx14_ASAP7_75t_R g1102 ( 
.A(n_661),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_203),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_232),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_705),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_192),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_532),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_412),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_22),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_628),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_219),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_487),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_337),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_579),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_702),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_53),
.Y(n_1116)
);

CKINVDCx14_ASAP7_75t_R g1117 ( 
.A(n_43),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_672),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_581),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_609),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_138),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_214),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_40),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_317),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_700),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_91),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_416),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_241),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_252),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_107),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_574),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_630),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_137),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_271),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_27),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_500),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_146),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_385),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_262),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_209),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_157),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_433),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_10),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_4),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_0),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_630),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_535),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_141),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_536),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_672),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_546),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_592),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_153),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_631),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_100),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_55),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_38),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_413),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_440),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_416),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_665),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_495),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_606),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_64),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_312),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_112),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_552),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_297),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_489),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_199),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_317),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_595),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_562),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_170),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_251),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_129),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_99),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_218),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_618),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_430),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_23),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_541),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_193),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_330),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_94),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_26),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_60),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_57),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_499),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_435),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_380),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_490),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_34),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_73),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_643),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_232),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_398),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_434),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_376),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_80),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_690),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_379),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_476),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_61),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_548),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_14),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_511),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_522),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_150),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_327),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_485),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_382),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_652),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_101),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_656),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_679),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_408),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_162),
.Y(n_1218)
);

CKINVDCx14_ASAP7_75t_R g1219 ( 
.A(n_110),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_211),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_55),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_282),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_34),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_258),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_450),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_452),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_65),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_615),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_479),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_536),
.Y(n_1230)
);

BUFx10_ASAP7_75t_L g1231 ( 
.A(n_670),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_194),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_279),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_113),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_38),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_81),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_237),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_354),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_173),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_51),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_79),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_178),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_560),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_676),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_389),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_626),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_44),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_100),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_442),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_234),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_716),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_716),
.Y(n_1252)
);

INVxp33_ASAP7_75t_L g1253 ( 
.A(n_830),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_974),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1041),
.Y(n_1255)
);

CKINVDCx16_ASAP7_75t_R g1256 ( 
.A(n_1004),
.Y(n_1256)
);

INVxp33_ASAP7_75t_SL g1257 ( 
.A(n_830),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_716),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_716),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_716),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_716),
.Y(n_1261)
);

INVxp33_ASAP7_75t_L g1262 ( 
.A(n_875),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_716),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_716),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1041),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_716),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_716),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_716),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_893),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_893),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_893),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_893),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_893),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_893),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_893),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_893),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_893),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_893),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1102),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1144),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_893),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_917),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_917),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_857),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_1004),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_917),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_1144),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_857),
.Y(n_1288)
);

INVxp33_ASAP7_75t_SL g1289 ( 
.A(n_875),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_917),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1204),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_917),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_1144),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_917),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_917),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_917),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_917),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1102),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_1204),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_917),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_917),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1047),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1144),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1120),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_769),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_714),
.B(n_0),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1047),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1047),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1047),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1047),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1047),
.Y(n_1311)
);

CKINVDCx16_ASAP7_75t_R g1312 ( 
.A(n_712),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1047),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_1144),
.Y(n_1314)
);

INVxp33_ASAP7_75t_L g1315 ( 
.A(n_903),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1047),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_769),
.Y(n_1317)
);

CKINVDCx16_ASAP7_75t_R g1318 ( 
.A(n_712),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1117),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1047),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1144),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_732),
.Y(n_1322)
);

CKINVDCx14_ASAP7_75t_R g1323 ( 
.A(n_1117),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_732),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_732),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1144),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_732),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_732),
.Y(n_1328)
);

CKINVDCx16_ASAP7_75t_R g1329 ( 
.A(n_764),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_974),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1120),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_732),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_732),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_974),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1219),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_739),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_739),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_739),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1219),
.B(n_1),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_739),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_739),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_739),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_903),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_764),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_739),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1062),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1062),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1062),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_819),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1062),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1062),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1062),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1062),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1111),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1111),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_819),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1111),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1111),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1111),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1223),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1111),
.Y(n_1361)
);

INVxp67_ASAP7_75t_SL g1362 ( 
.A(n_1223),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1111),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_772),
.B(n_1),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1226),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1018),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1226),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1226),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1223),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1226),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1018),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1226),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1226),
.Y(n_1373)
);

INVxp33_ASAP7_75t_SL g1374 ( 
.A(n_933),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1226),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_765),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_819),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_976),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_976),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_849),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_933),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_849),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_976),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1049),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_757),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_765),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1049),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1049),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1075),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_805),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_805),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1075),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1075),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_815),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_848),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_807),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_807),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_848),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_807),
.Y(n_1399)
);

CKINVDCx16_ASAP7_75t_R g1400 ( 
.A(n_912),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_808),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_808),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_808),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_849),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_912),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1029),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_868),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_910),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_910),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_910),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_973),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_883),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_924),
.Y(n_1413)
);

INVxp33_ASAP7_75t_SL g1414 ( 
.A(n_1029),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_924),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_973),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1122),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_973),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_975),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_975),
.Y(n_1420)
);

INVxp33_ASAP7_75t_SL g1421 ( 
.A(n_1122),
.Y(n_1421)
);

INVxp33_ASAP7_75t_L g1422 ( 
.A(n_1127),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_975),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_979),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_979),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_979),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1017),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_990),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1031),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_868),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_868),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_925),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_925),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_925),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1063),
.Y(n_1435)
);

INVxp33_ASAP7_75t_SL g1436 ( 
.A(n_1127),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_955),
.Y(n_1437)
);

INVxp67_ASAP7_75t_SL g1438 ( 
.A(n_955),
.Y(n_1438)
);

INVxp33_ASAP7_75t_SL g1439 ( 
.A(n_1131),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1063),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_955),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_982),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_982),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1131),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_982),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1203),
.Y(n_1446)
);

CKINVDCx16_ASAP7_75t_R g1447 ( 
.A(n_1203),
.Y(n_1447)
);

INVxp33_ASAP7_75t_SL g1448 ( 
.A(n_1172),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1010),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1010),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_990),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_707),
.Y(n_1452)
);

INVxp33_ASAP7_75t_L g1453 ( 
.A(n_1172),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_708),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1010),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_990),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1021),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1021),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1021),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1022),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1241),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1022),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1022),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1008),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_817),
.Y(n_1465)
);

INVxp33_ASAP7_75t_SL g1466 ( 
.A(n_733),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1023),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1023),
.Y(n_1468)
);

CKINVDCx14_ASAP7_75t_R g1469 ( 
.A(n_1241),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1023),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1099),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1008),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1140),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1099),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1008),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1099),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_817),
.Y(n_1477)
);

BUFx8_ASAP7_75t_SL g1478 ( 
.A(n_963),
.Y(n_1478)
);

CKINVDCx14_ASAP7_75t_R g1479 ( 
.A(n_1241),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_963),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1115),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1032),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1115),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1115),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_745),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1171),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_709),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1171),
.Y(n_1488)
);

INVxp33_ASAP7_75t_L g1489 ( 
.A(n_714),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1171),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1197),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_710),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1197),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_715),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1032),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1197),
.Y(n_1496)
);

INVxp33_ASAP7_75t_L g1497 ( 
.A(n_753),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1205),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1205),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1205),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1209),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1209),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1209),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_772),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_753),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_789),
.Y(n_1506)
);

INVxp33_ASAP7_75t_SL g1507 ( 
.A(n_758),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_789),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_784),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_772),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1145),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_798),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1240),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1240),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_798),
.Y(n_1515)
);

CKINVDCx16_ASAP7_75t_R g1516 ( 
.A(n_1241),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1240),
.Y(n_1517)
);

INVxp33_ASAP7_75t_L g1518 ( 
.A(n_821),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_821),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_841),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_717),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_841),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_909),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1032),
.Y(n_1524)
);

BUFx10_ASAP7_75t_L g1525 ( 
.A(n_752),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_720),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1056),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_909),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_787),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_916),
.Y(n_1530)
);

INVxp33_ASAP7_75t_L g1531 ( 
.A(n_916),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_936),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1123),
.Y(n_1533)
);

INVxp33_ASAP7_75t_SL g1534 ( 
.A(n_785),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_936),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_787),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_940),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1056),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_940),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_966),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_721),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_966),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1003),
.Y(n_1543)
);

INVxp33_ASAP7_75t_SL g1544 ( 
.A(n_810),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1003),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1026),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1026),
.Y(n_1547)
);

BUFx2_ASAP7_75t_SL g1548 ( 
.A(n_752),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1061),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1061),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1093),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1056),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1069),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_724),
.Y(n_1554)
);

INVxp33_ASAP7_75t_L g1555 ( 
.A(n_1093),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_728),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1116),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_734),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1116),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1143),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1069),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1069),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_737),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_847),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1143),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1156),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1156),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1157),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1157),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1188),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_738),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1188),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1200),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_842),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_740),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_741),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1123),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1200),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1090),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1206),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1206),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_711),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_711),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_742),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_713),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_713),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_718),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1241),
.Y(n_1588)
);

INVxp33_ASAP7_75t_L g1589 ( 
.A(n_718),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1090),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1090),
.Y(n_1591)
);

INVxp33_ASAP7_75t_SL g1592 ( 
.A(n_873),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1100),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_743),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1100),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1100),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1126),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1126),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1126),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1148),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1148),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1148),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_744),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1149),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1149),
.Y(n_1605)
);

INVxp33_ASAP7_75t_SL g1606 ( 
.A(n_889),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1149),
.Y(n_1607)
);

XOR2x2_ASAP7_75t_L g1608 ( 
.A(n_736),
.B(n_2),
.Y(n_1608)
);

INVxp67_ASAP7_75t_SL g1609 ( 
.A(n_1153),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1153),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1153),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1201),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1164),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1162),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_759),
.Y(n_1615)
);

INVxp33_ASAP7_75t_L g1616 ( 
.A(n_719),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1201),
.Y(n_1617)
);

INVxp33_ASAP7_75t_L g1618 ( 
.A(n_719),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1201),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_748),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1218),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1218),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_777),
.B(n_2),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1218),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_722),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_751),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1164),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_755),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_722),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_847),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_760),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_913),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_752),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_900),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_762),
.Y(n_1635)
);

CKINVDCx16_ASAP7_75t_R g1636 ( 
.A(n_759),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_723),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_759),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_763),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_723),
.Y(n_1640)
);

INVxp33_ASAP7_75t_L g1641 ( 
.A(n_725),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1250),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_766),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_725),
.Y(n_1644)
);

CKINVDCx16_ASAP7_75t_R g1645 ( 
.A(n_759),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_726),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_726),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_767),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_727),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_727),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_778),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_913),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_729),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_729),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_730),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_768),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_770),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_730),
.Y(n_1658)
);

CKINVDCx16_ASAP7_75t_R g1659 ( 
.A(n_759),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_731),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_783),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_731),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_735),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_911),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_735),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_746),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_783),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_746),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_747),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_747),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_749),
.B(n_2),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_749),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_780),
.Y(n_1673)
);

CKINVDCx16_ASAP7_75t_R g1674 ( 
.A(n_783),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_781),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_754),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_754),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_782),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_950),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_756),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_788),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_778),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_756),
.Y(n_1683)
);

INVxp33_ASAP7_75t_L g1684 ( 
.A(n_771),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_950),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1162),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1002),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_771),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_778),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_887),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_773),
.Y(n_1691)
);

CKINVDCx16_ASAP7_75t_R g1692 ( 
.A(n_783),
.Y(n_1692)
);

NOR2xp67_ASAP7_75t_L g1693 ( 
.A(n_774),
.B(n_3),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_773),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1303),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1280),
.B(n_887),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1466),
.B(n_1507),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1303),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1360),
.B(n_887),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1303),
.Y(n_1701)
);

XNOR2xp5_ASAP7_75t_L g1702 ( 
.A(n_1608),
.B(n_1193),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1303),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1362),
.B(n_897),
.Y(n_1704)
);

BUFx8_ASAP7_75t_SL g1705 ( 
.A(n_1478),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1369),
.B(n_897),
.Y(n_1706)
);

INVx5_ASAP7_75t_L g1707 ( 
.A(n_1303),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1525),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1382),
.B(n_897),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1504),
.B(n_898),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1464),
.Y(n_1711)
);

BUFx12f_ASAP7_75t_L g1712 ( 
.A(n_1331),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1326),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1510),
.B(n_898),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1326),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1326),
.Y(n_1716)
);

INVx5_ASAP7_75t_L g1717 ( 
.A(n_1326),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1287),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1407),
.B(n_898),
.Y(n_1719)
);

INVx5_ASAP7_75t_L g1720 ( 
.A(n_1326),
.Y(n_1720)
);

INVx5_ASAP7_75t_L g1721 ( 
.A(n_1464),
.Y(n_1721)
);

XNOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1608),
.B(n_928),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1293),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1380),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1321),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1314),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1321),
.Y(n_1728)
);

BUFx8_ASAP7_75t_L g1729 ( 
.A(n_1615),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1438),
.B(n_962),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1524),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1380),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1517),
.B(n_962),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1404),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1322),
.B(n_775),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1372),
.B(n_962),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1534),
.B(n_777),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1544),
.B(n_969),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1464),
.Y(n_1739)
);

INVx5_ASAP7_75t_L g1740 ( 
.A(n_1464),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1464),
.Y(n_1741)
);

INVx5_ASAP7_75t_L g1742 ( 
.A(n_1527),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1375),
.B(n_969),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1633),
.B(n_969),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1331),
.B(n_783),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1254),
.B(n_1034),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1254),
.B(n_1034),
.Y(n_1747)
);

INVxp33_ASAP7_75t_SL g1748 ( 
.A(n_1319),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1527),
.Y(n_1749)
);

BUFx12f_ASAP7_75t_L g1750 ( 
.A(n_1305),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1651),
.B(n_1034),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1538),
.B(n_1040),
.Y(n_1752)
);

BUFx8_ASAP7_75t_SL g1753 ( 
.A(n_1529),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1319),
.B(n_790),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1553),
.B(n_1040),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1561),
.B(n_1040),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1322),
.B(n_775),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1527),
.Y(n_1758)
);

AND2x6_ASAP7_75t_L g1759 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1579),
.B(n_1609),
.Y(n_1760)
);

BUFx12f_ASAP7_75t_L g1761 ( 
.A(n_1305),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1527),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1592),
.B(n_1125),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1682),
.B(n_1125),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1404),
.B(n_1125),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1471),
.B(n_1163),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1527),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1642),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1606),
.B(n_1163),
.Y(n_1769)
);

BUFx12f_ASAP7_75t_L g1770 ( 
.A(n_1317),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1642),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1323),
.B(n_1163),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1689),
.B(n_1690),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1548),
.B(n_776),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1430),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1431),
.Y(n_1776)
);

INVx5_ASAP7_75t_L g1777 ( 
.A(n_1642),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1548),
.B(n_776),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1614),
.B(n_951),
.Y(n_1779)
);

BUFx12f_ASAP7_75t_L g1780 ( 
.A(n_1317),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1471),
.B(n_779),
.Y(n_1781)
);

INVx5_ASAP7_75t_L g1782 ( 
.A(n_1642),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1686),
.B(n_968),
.Y(n_1783)
);

BUFx8_ASAP7_75t_SL g1784 ( 
.A(n_1536),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1339),
.B(n_983),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_SL g1786 ( 
.A(n_1255),
.B(n_790),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1474),
.B(n_779),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1474),
.B(n_786),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1432),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1433),
.B(n_786),
.Y(n_1790)
);

BUFx8_ASAP7_75t_L g1791 ( 
.A(n_1615),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1642),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1434),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1437),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1257),
.B(n_1013),
.Y(n_1795)
);

BUFx8_ASAP7_75t_SL g1796 ( 
.A(n_1564),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1644),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1469),
.B(n_1044),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1644),
.Y(n_1799)
);

INVx5_ASAP7_75t_L g1800 ( 
.A(n_1644),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1441),
.B(n_792),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1442),
.B(n_792),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1644),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1443),
.B(n_793),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1289),
.B(n_1374),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1445),
.Y(n_1806)
);

BUFx12f_ASAP7_75t_L g1807 ( 
.A(n_1284),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1449),
.B(n_793),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1450),
.Y(n_1809)
);

CKINVDCx16_ASAP7_75t_R g1810 ( 
.A(n_1265),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1644),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1349),
.Y(n_1812)
);

BUFx12f_ASAP7_75t_L g1813 ( 
.A(n_1284),
.Y(n_1813)
);

INVx5_ASAP7_75t_L g1814 ( 
.A(n_1268),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1414),
.B(n_1046),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1349),
.Y(n_1816)
);

INVx5_ASAP7_75t_L g1817 ( 
.A(n_1268),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1356),
.Y(n_1818)
);

BUFx8_ASAP7_75t_SL g1819 ( 
.A(n_1630),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1376),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1455),
.Y(n_1821)
);

BUFx12f_ASAP7_75t_L g1822 ( 
.A(n_1288),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1457),
.B(n_796),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1356),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1377),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1482),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1458),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1421),
.B(n_1068),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1459),
.B(n_796),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1376),
.Y(n_1830)
);

BUFx12f_ASAP7_75t_L g1831 ( 
.A(n_1288),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1436),
.B(n_1109),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1479),
.B(n_1135),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1460),
.B(n_802),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1462),
.B(n_802),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1439),
.B(n_1181),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1463),
.B(n_809),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1448),
.B(n_1186),
.Y(n_1838)
);

BUFx8_ASAP7_75t_L g1839 ( 
.A(n_1577),
.Y(n_1839)
);

BUFx12f_ASAP7_75t_L g1840 ( 
.A(n_1386),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1377),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1378),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1378),
.Y(n_1843)
);

BUFx12f_ASAP7_75t_L g1844 ( 
.A(n_1386),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1279),
.B(n_790),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1638),
.B(n_1187),
.Y(n_1846)
);

BUFx8_ASAP7_75t_SL g1847 ( 
.A(n_1632),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1387),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1525),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1638),
.B(n_1221),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1467),
.B(n_809),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1387),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1399),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1468),
.B(n_812),
.Y(n_1854)
);

BUFx12f_ASAP7_75t_L g1855 ( 
.A(n_1390),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1399),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1298),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1470),
.B(n_1476),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1481),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1483),
.B(n_812),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1304),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1511),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1390),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1661),
.B(n_1227),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1484),
.B(n_816),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1324),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1525),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1486),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1324),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1488),
.B(n_816),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1490),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1451),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1491),
.B(n_1493),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1451),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1456),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1661),
.B(n_1235),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1456),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1496),
.Y(n_1878)
);

CKINVDCx6p67_ASAP7_75t_R g1879 ( 
.A(n_1335),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1498),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1667),
.B(n_1236),
.Y(n_1881)
);

INVx5_ASAP7_75t_L g1882 ( 
.A(n_1482),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1499),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1667),
.B(n_1247),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1500),
.B(n_791),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1501),
.B(n_795),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1502),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1503),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1325),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1325),
.B(n_820),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1489),
.B(n_820),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1327),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1636),
.B(n_790),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1327),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1269),
.B(n_797),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1328),
.B(n_825),
.Y(n_1896)
);

CKINVDCx11_ASAP7_75t_R g1897 ( 
.A(n_1652),
.Y(n_1897)
);

BUFx8_ASAP7_75t_SL g1898 ( 
.A(n_1679),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1452),
.B(n_774),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1328),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1270),
.B(n_799),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1332),
.Y(n_1902)
);

AND2x6_ASAP7_75t_L g1903 ( 
.A(n_1251),
.B(n_825),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1332),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1333),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1333),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1336),
.Y(n_1907)
);

BUFx12f_ASAP7_75t_L g1908 ( 
.A(n_1391),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1336),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1337),
.B(n_831),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1391),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1395),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1475),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1475),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1337),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1338),
.B(n_831),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1271),
.B(n_800),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1338),
.Y(n_1918)
);

AND2x6_ASAP7_75t_L g1919 ( 
.A(n_1252),
.B(n_832),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1340),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1495),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1485),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1340),
.B(n_832),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1452),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1341),
.B(n_833),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1497),
.B(n_833),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1454),
.B(n_1176),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1518),
.B(n_1531),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1495),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1272),
.B(n_801),
.Y(n_1930)
);

BUFx12f_ASAP7_75t_L g1931 ( 
.A(n_1395),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1341),
.Y(n_1932)
);

INVx5_ASAP7_75t_L g1933 ( 
.A(n_1482),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1342),
.Y(n_1934)
);

INVx5_ASAP7_75t_L g1935 ( 
.A(n_1552),
.Y(n_1935)
);

BUFx12f_ASAP7_75t_L g1936 ( 
.A(n_1398),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1398),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1555),
.B(n_836),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1342),
.B(n_836),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1405),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1552),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1273),
.B(n_804),
.Y(n_1942)
);

INVx5_ASAP7_75t_L g1943 ( 
.A(n_1562),
.Y(n_1943)
);

BUFx8_ASAP7_75t_L g1944 ( 
.A(n_1577),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1345),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1562),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1601),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1589),
.B(n_840),
.Y(n_1949)
);

INVx5_ASAP7_75t_L g1950 ( 
.A(n_1601),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1274),
.B(n_806),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1616),
.B(n_840),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1405),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1346),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1347),
.Y(n_1955)
);

INVx5_ASAP7_75t_L g1956 ( 
.A(n_1604),
.Y(n_1956)
);

CKINVDCx20_ASAP7_75t_R g1957 ( 
.A(n_1685),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1509),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1604),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1413),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1454),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1275),
.B(n_811),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1607),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1607),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1347),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1618),
.B(n_843),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1487),
.B(n_1176),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1645),
.B(n_790),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1348),
.B(n_843),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1348),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1350),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1610),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1350),
.B(n_845),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1351),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1610),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1621),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1351),
.B(n_845),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1574),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1352),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1352),
.Y(n_1980)
);

AND2x6_ASAP7_75t_L g1981 ( 
.A(n_1258),
.B(n_846),
.Y(n_1981)
);

NOR2x1_ASAP7_75t_L g1982 ( 
.A(n_1353),
.B(n_846),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1276),
.B(n_813),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1413),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1353),
.B(n_851),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1487),
.B(n_814),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1621),
.Y(n_1987)
);

INVx5_ASAP7_75t_L g1988 ( 
.A(n_1624),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1492),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1277),
.B(n_818),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1354),
.Y(n_1991)
);

INVx5_ASAP7_75t_L g1992 ( 
.A(n_1624),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1278),
.B(n_1281),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1282),
.B(n_822),
.Y(n_1994)
);

INVx5_ASAP7_75t_L g1995 ( 
.A(n_1646),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1492),
.B(n_823),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1354),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1494),
.B(n_826),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1355),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1355),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1357),
.B(n_1358),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1283),
.B(n_827),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1357),
.Y(n_2003)
);

INVx5_ASAP7_75t_L g2004 ( 
.A(n_1646),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1358),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1359),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1359),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1494),
.B(n_828),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1361),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1415),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1361),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1654),
.Y(n_2012)
);

BUFx8_ASAP7_75t_L g2013 ( 
.A(n_1613),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1363),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1363),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1365),
.Y(n_2016)
);

INVx5_ASAP7_75t_L g2017 ( 
.A(n_1654),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1521),
.B(n_829),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1461),
.B(n_824),
.Y(n_2019)
);

AND2x2_ASAP7_75t_SL g2020 ( 
.A(n_1623),
.B(n_851),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1365),
.Y(n_2021)
);

INVx5_ASAP7_75t_L g2022 ( 
.A(n_1680),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1367),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1367),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1368),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1286),
.B(n_834),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1290),
.B(n_835),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1521),
.B(n_838),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1368),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1370),
.Y(n_2030)
);

INVx5_ASAP7_75t_L g2031 ( 
.A(n_1680),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1526),
.B(n_839),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1370),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1526),
.B(n_844),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1373),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1634),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1415),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1373),
.B(n_855),
.Y(n_2038)
);

BUFx12f_ASAP7_75t_L g2039 ( 
.A(n_1435),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1379),
.Y(n_2040)
);

INVx4_ASAP7_75t_L g2041 ( 
.A(n_1258),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1505),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1259),
.B(n_855),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1259),
.B(n_860),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1260),
.Y(n_2045)
);

INVx4_ASAP7_75t_L g2046 ( 
.A(n_1260),
.Y(n_2046)
);

INVx5_ASAP7_75t_L g2047 ( 
.A(n_1516),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1379),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1541),
.B(n_852),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1383),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1541),
.B(n_853),
.Y(n_2051)
);

BUFx8_ASAP7_75t_L g2052 ( 
.A(n_1613),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1383),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1554),
.B(n_854),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1659),
.B(n_824),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1695),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1816),
.Y(n_2057)
);

AND2x2_ASAP7_75t_SL g2058 ( 
.A(n_2020),
.B(n_1364),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_2043),
.B(n_1396),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1695),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1718),
.B(n_1554),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1816),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1946),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1725),
.Y(n_2064)
);

CKINVDCx8_ASAP7_75t_R g2065 ( 
.A(n_1810),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1695),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_2043),
.B(n_1396),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1928),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1816),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1816),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1816),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1723),
.B(n_1556),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1928),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1759),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1818),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1726),
.B(n_1384),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1818),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1946),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1946),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1726),
.B(n_1384),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2001),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1710),
.B(n_1388),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2001),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2001),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_2043),
.B(n_1397),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1900),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1708),
.B(n_1588),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1818),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1900),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1818),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1725),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1710),
.B(n_1388),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1695),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1862),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2044),
.B(n_1397),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1714),
.B(n_1389),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1695),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2020),
.A2(n_1193),
.B1(n_1042),
.B2(n_1057),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1907),
.Y(n_2099)
);

AND3x1_ASAP7_75t_L g2100 ( 
.A(n_1805),
.B(n_1477),
.C(n_1465),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1907),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1818),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1701),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1701),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1920),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1714),
.B(n_1389),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1724),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1825),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1727),
.B(n_1556),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1825),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_SL g2111 ( 
.A1(n_1702),
.A2(n_1042),
.B1(n_1057),
.B2(n_1002),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1701),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1920),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1760),
.B(n_1736),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1955),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1825),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1733),
.B(n_1392),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1733),
.B(n_1392),
.Y(n_2118)
);

NAND2x1p5_ASAP7_75t_L g2119 ( 
.A(n_2044),
.B(n_1671),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_1724),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1701),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2044),
.B(n_1401),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1955),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1979),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_1890),
.B(n_1401),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1774),
.B(n_1393),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1753),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1825),
.Y(n_2128)
);

AND2x6_ASAP7_75t_L g2129 ( 
.A(n_1736),
.B(n_1261),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1825),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1979),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1701),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1715),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1760),
.B(n_1558),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_1715),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1760),
.B(n_1558),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_1890),
.B(n_1402),
.Y(n_2137)
);

NAND2xp33_ASAP7_75t_L g2138 ( 
.A(n_1846),
.B(n_1563),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_1732),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1991),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1841),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1841),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1841),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1715),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_1732),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1991),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1736),
.B(n_1563),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1841),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_SL g2149 ( 
.A1(n_1702),
.A2(n_1059),
.B1(n_1064),
.B2(n_1058),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_1986),
.B(n_1571),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1997),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1728),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1997),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2011),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1890),
.B(n_1402),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1774),
.B(n_1393),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1728),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1889),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1778),
.B(n_1403),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1896),
.B(n_1403),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1896),
.B(n_1408),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2011),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2024),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1896),
.B(n_1408),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2024),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1743),
.B(n_1696),
.Y(n_2166)
);

AND2x6_ASAP7_75t_L g2167 ( 
.A(n_1743),
.B(n_1261),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1841),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1715),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1743),
.B(n_1571),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2035),
.Y(n_2171)
);

BUFx2_ASAP7_75t_L g2172 ( 
.A(n_1734),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2035),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2045),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2045),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1778),
.B(n_1409),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1696),
.B(n_1575),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1892),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1715),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1744),
.B(n_1409),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1894),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1902),
.Y(n_2182)
);

OA21x2_ASAP7_75t_L g2183 ( 
.A1(n_1904),
.A2(n_1264),
.B(n_1263),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1716),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1785),
.A2(n_1737),
.B1(n_1783),
.B2(n_1779),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1842),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1996),
.B(n_1575),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1905),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1915),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1974),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2015),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1842),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1759),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1842),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1759),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1842),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1744),
.B(n_1410),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1842),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1759),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1734),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1759),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1759),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1716),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1843),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_1883),
.Y(n_2205)
);

INVx4_ASAP7_75t_L g2206 ( 
.A(n_1814),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1993),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1716),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1843),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1866),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1866),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_1708),
.B(n_1674),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1716),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1843),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1910),
.B(n_1410),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_SL g2216 ( 
.A(n_2019),
.B(n_1312),
.Y(n_2216)
);

CKINVDCx6p67_ASAP7_75t_R g2217 ( 
.A(n_2047),
.Y(n_2217)
);

AND2x6_ASAP7_75t_L g2218 ( 
.A(n_1696),
.B(n_1263),
.Y(n_2218)
);

BUFx8_ASAP7_75t_L g2219 ( 
.A(n_1857),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1843),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_1910),
.B(n_1411),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1843),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1866),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1773),
.B(n_1576),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_1849),
.B(n_1692),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1716),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1751),
.B(n_1411),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_1814),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1869),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1852),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1739),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_1903),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_1751),
.B(n_1416),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1699),
.B(n_1576),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_1891),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1700),
.B(n_1416),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_SL g2237 ( 
.A(n_2047),
.B(n_1318),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1891),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1849),
.B(n_1584),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1869),
.Y(n_2240)
);

INVxp67_ASAP7_75t_SL g2241 ( 
.A(n_1739),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1998),
.B(n_1584),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1699),
.B(n_1594),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_1739),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1852),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1869),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_1700),
.B(n_1418),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1852),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1852),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1852),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1753),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1934),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1704),
.B(n_1418),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1934),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1910),
.B(n_1419),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1934),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1954),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1954),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1704),
.B(n_1419),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1873),
.B(n_1420),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1853),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1853),
.Y(n_2262)
);

OA21x2_ASAP7_75t_L g2263 ( 
.A1(n_1895),
.A2(n_1266),
.B(n_1264),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_1883),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1954),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1873),
.B(n_1420),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1999),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1999),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2041),
.B(n_1594),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2041),
.B(n_1603),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2041),
.B(n_1603),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1999),
.Y(n_2272)
);

BUFx2_ASAP7_75t_L g2273 ( 
.A(n_2010),
.Y(n_2273)
);

OA21x2_ASAP7_75t_L g2274 ( 
.A1(n_1901),
.A2(n_1930),
.B(n_1917),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1853),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2046),
.B(n_1620),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2000),
.Y(n_2277)
);

OR2x6_ASAP7_75t_L g2278 ( 
.A(n_1840),
.B(n_1306),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_1795),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_1903),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2016),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1752),
.B(n_1423),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1889),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2016),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_1916),
.B(n_1423),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2008),
.B(n_1620),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1739),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2016),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1739),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1906),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1758),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_1758),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2033),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2000),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1906),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_1815),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2033),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_1916),
.B(n_1424),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1853),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1758),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2018),
.B(n_1626),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1853),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1758),
.Y(n_2303)
);

NAND2x1_ASAP7_75t_L g2304 ( 
.A(n_1903),
.B(n_1266),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_SL g2305 ( 
.A1(n_1828),
.A2(n_1059),
.B1(n_1064),
.B2(n_1058),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_1916),
.B(n_1424),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2046),
.B(n_1626),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_2000),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_1903),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1752),
.B(n_1425),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1856),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2000),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1758),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1856),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1856),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2046),
.B(n_1628),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2033),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1923),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1856),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1768),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_1768),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2000),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1752),
.B(n_1628),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1923),
.Y(n_2324)
);

HB1xp67_ASAP7_75t_L g2325 ( 
.A(n_1926),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_1755),
.B(n_1425),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2003),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1923),
.Y(n_2328)
);

OR2x6_ASAP7_75t_L g2329 ( 
.A(n_1840),
.B(n_1306),
.Y(n_2329)
);

AND2x6_ASAP7_75t_L g2330 ( 
.A(n_1755),
.B(n_1267),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1925),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_1755),
.B(n_1426),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1856),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_2003),
.Y(n_2334)
);

OA21x2_ASAP7_75t_L g2335 ( 
.A1(n_1942),
.A2(n_1292),
.B(n_1267),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_1784),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2003),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_1925),
.B(n_1426),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2003),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_1756),
.B(n_1428),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_1925),
.B(n_1939),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1939),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1939),
.Y(n_2343)
);

OA21x2_ASAP7_75t_L g2344 ( 
.A1(n_1951),
.A2(n_1294),
.B(n_1292),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_1832),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_1969),
.B(n_1428),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1969),
.Y(n_2347)
);

OA21x2_ASAP7_75t_L g2348 ( 
.A1(n_1962),
.A2(n_1295),
.B(n_1294),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1872),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_1768),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_1969),
.B(n_1472),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1973),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1872),
.Y(n_2353)
);

INVx4_ASAP7_75t_L g2354 ( 
.A(n_1814),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1872),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1872),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1973),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2010),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1973),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2003),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2005),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1977),
.Y(n_2362)
);

BUFx2_ASAP7_75t_L g2363 ( 
.A(n_1922),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_1768),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2051),
.B(n_2028),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1872),
.Y(n_2366)
);

BUFx2_ASAP7_75t_L g2367 ( 
.A(n_1926),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1977),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1977),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1985),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1874),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_1768),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1756),
.B(n_1631),
.Y(n_2373)
);

INVx3_ASAP7_75t_L g2374 ( 
.A(n_2005),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1985),
.Y(n_2375)
);

XNOR2xp5_ASAP7_75t_L g2376 ( 
.A(n_1722),
.B(n_1687),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1874),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1985),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1874),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2038),
.Y(n_2380)
);

BUFx8_ASAP7_75t_L g2381 ( 
.A(n_1861),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1756),
.B(n_1631),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_1781),
.B(n_1472),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_1771),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1874),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2038),
.B(n_1590),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_1781),
.B(n_1590),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_1771),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2038),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1874),
.Y(n_2390)
);

INVx4_ASAP7_75t_L g2391 ( 
.A(n_1814),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1875),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1826),
.Y(n_2393)
);

HB1xp67_ASAP7_75t_L g2394 ( 
.A(n_1938),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1731),
.B(n_1635),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2005),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1826),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_1771),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1983),
.B(n_1635),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1875),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1875),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1826),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_1735),
.B(n_1591),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_1867),
.B(n_2047),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_1990),
.B(n_1639),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1741),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_2005),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_1909),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1741),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_1787),
.B(n_1591),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1909),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1757),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2032),
.B(n_1639),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1982),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_2005),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1811),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2007),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1875),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_2007),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1811),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1811),
.Y(n_2421)
);

NAND2xp33_ASAP7_75t_L g2422 ( 
.A(n_1850),
.B(n_1643),
.Y(n_2422)
);

CKINVDCx11_ASAP7_75t_R g2423 ( 
.A(n_1897),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1749),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_1787),
.B(n_1593),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_1771),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1749),
.Y(n_2427)
);

BUFx6f_ASAP7_75t_L g2428 ( 
.A(n_1771),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2034),
.B(n_1643),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1749),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1762),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_1792),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_1875),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_1784),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1792),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_1994),
.B(n_1648),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_1796),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1762),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2002),
.B(n_1648),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1762),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1767),
.Y(n_2441)
);

BUFx8_ASAP7_75t_L g2442 ( 
.A(n_1807),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_1938),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_1949),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1767),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_1801),
.B(n_1593),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1877),
.Y(n_2447)
);

INVx3_ASAP7_75t_L g2448 ( 
.A(n_2007),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1767),
.Y(n_2449)
);

INVx3_ASAP7_75t_L g2450 ( 
.A(n_2007),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2049),
.B(n_1656),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1877),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1877),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1877),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_2007),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_1918),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_1918),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_1932),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_1788),
.B(n_1595),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_1792),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1877),
.Y(n_2461)
);

XOR2xp5_ASAP7_75t_L g2462 ( 
.A(n_1722),
.B(n_1385),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_1913),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_1913),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1913),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_1949),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2026),
.B(n_1656),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_1867),
.B(n_1657),
.Y(n_2468)
);

BUFx6f_ASAP7_75t_L g2469 ( 
.A(n_1792),
.Y(n_2469)
);

BUFx6f_ASAP7_75t_L g2470 ( 
.A(n_1792),
.Y(n_2470)
);

AND2x6_ASAP7_75t_L g2471 ( 
.A(n_1765),
.B(n_1295),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_1788),
.B(n_1595),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1913),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_1864),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_1858),
.B(n_1596),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2027),
.B(n_1657),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2047),
.B(n_1673),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_1913),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_1797),
.Y(n_2479)
);

BUFx6f_ASAP7_75t_L g2480 ( 
.A(n_1797),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1797),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2279),
.B(n_2296),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2183),
.Y(n_2483)
);

OAI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2185),
.A2(n_1845),
.B1(n_1786),
.B2(n_1958),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_2185),
.B(n_2047),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2183),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2318),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2471),
.Y(n_2488)
);

AND2x2_ASAP7_75t_SL g2489 ( 
.A(n_2058),
.B(n_1763),
.Y(n_2489)
);

NAND2xp33_ASAP7_75t_R g2490 ( 
.A(n_2273),
.B(n_1924),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2318),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2324),
.Y(n_2492)
);

AO21x2_ASAP7_75t_L g2493 ( 
.A1(n_2166),
.A2(n_2054),
.B(n_1881),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2074),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2183),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2324),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2328),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2183),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2328),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2064),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2367),
.B(n_1958),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2367),
.B(n_1978),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2331),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2443),
.B(n_1978),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2365),
.B(n_1903),
.Y(n_2505)
);

OAI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_2207),
.A2(n_2036),
.B1(n_1884),
.B2(n_1876),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2064),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2345),
.B(n_1748),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2443),
.B(n_2036),
.Y(n_2509)
);

INVxp67_ASAP7_75t_SL g2510 ( 
.A(n_2114),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2064),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2094),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2091),
.Y(n_2513)
);

INVx2_ASAP7_75t_SL g2514 ( 
.A(n_2383),
.Y(n_2514)
);

NOR2x1p5_ASAP7_75t_L g2515 ( 
.A(n_2323),
.B(n_1712),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2331),
.Y(n_2516)
);

NAND2xp33_ASAP7_75t_SL g2517 ( 
.A(n_2212),
.B(n_1924),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2091),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2207),
.B(n_1903),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2091),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2341),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2152),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2059),
.Y(n_2523)
);

HB1xp67_ASAP7_75t_L g2524 ( 
.A(n_2068),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2076),
.B(n_2080),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2373),
.B(n_2382),
.Y(n_2526)
);

INVx4_ASAP7_75t_L g2527 ( 
.A(n_2129),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2383),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2342),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2224),
.B(n_1697),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2134),
.B(n_1729),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2342),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2076),
.B(n_2080),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2343),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2282),
.B(n_1765),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2150),
.B(n_1748),
.Y(n_2536)
);

OAI21xp33_ASAP7_75t_SL g2537 ( 
.A1(n_2058),
.A2(n_1769),
.B(n_1738),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2059),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2282),
.B(n_1919),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2059),
.Y(n_2540)
);

OR2x2_ASAP7_75t_L g2541 ( 
.A(n_2234),
.B(n_1533),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2136),
.B(n_1729),
.Y(n_2542)
);

NAND3xp33_ASAP7_75t_L g2543 ( 
.A(n_2243),
.B(n_1927),
.C(n_1899),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2343),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2347),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2423),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2347),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2187),
.B(n_1961),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2059),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2352),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2352),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2067),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2357),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2357),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2058),
.A2(n_1981),
.B1(n_1919),
.B2(n_1967),
.Y(n_2555)
);

BUFx10_ASAP7_75t_L g2556 ( 
.A(n_2242),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2067),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_2074),
.Y(n_2558)
);

NAND3xp33_ASAP7_75t_L g2559 ( 
.A(n_2147),
.B(n_1838),
.C(n_1836),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2286),
.B(n_1961),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2301),
.B(n_1989),
.Y(n_2561)
);

OAI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2170),
.A2(n_2177),
.B1(n_2216),
.B2(n_2119),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2359),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2067),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2413),
.B(n_1989),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2067),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2310),
.B(n_1919),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2152),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2152),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2157),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2157),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2341),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2429),
.B(n_1729),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2387),
.Y(n_2574)
);

INVx4_ASAP7_75t_L g2575 ( 
.A(n_2129),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2451),
.B(n_1791),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2157),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2359),
.Y(n_2578)
);

INVx4_ASAP7_75t_L g2579 ( 
.A(n_2129),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_2387),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2310),
.B(n_1919),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2158),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2362),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2158),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2326),
.B(n_1919),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2362),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2158),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2283),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2474),
.B(n_1791),
.Y(n_2589)
);

INVx2_ASAP7_75t_SL g2590 ( 
.A(n_2410),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2326),
.B(n_1919),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2341),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2332),
.A2(n_2340),
.B1(n_2156),
.B2(n_2126),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2474),
.B(n_1791),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2332),
.B(n_1981),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2129),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2283),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2399),
.B(n_1798),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2368),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2368),
.Y(n_2600)
);

NOR2x1p5_ASAP7_75t_L g2601 ( 
.A(n_2217),
.B(n_1712),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2405),
.B(n_1329),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2283),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2369),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2369),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2370),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2290),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2370),
.Y(n_2608)
);

AND3x2_ASAP7_75t_L g2609 ( 
.A(n_2237),
.B(n_1244),
.C(n_1912),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2290),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2375),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2340),
.B(n_1981),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2074),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2375),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2129),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_2085),
.A2(n_1981),
.B1(n_1766),
.B2(n_1765),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2290),
.Y(n_2617)
);

NAND3xp33_ASAP7_75t_L g2618 ( 
.A(n_2073),
.B(n_1675),
.C(n_1673),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2378),
.Y(n_2619)
);

AOI22x1_ASAP7_75t_L g2620 ( 
.A1(n_2193),
.A2(n_2195),
.B1(n_2201),
.B2(n_2199),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2273),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2180),
.B(n_1981),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2378),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2380),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2180),
.B(n_2197),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_SL g2626 ( 
.A(n_2436),
.B(n_1833),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_2410),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2341),
.Y(n_2628)
);

AND3x2_ASAP7_75t_L g2629 ( 
.A(n_2358),
.B(n_1244),
.C(n_1940),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2085),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2380),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2205),
.B(n_2264),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2363),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2439),
.B(n_1344),
.Y(n_2634)
);

INVx2_ASAP7_75t_SL g2635 ( 
.A(n_2425),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2467),
.B(n_1400),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2389),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2389),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2363),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2063),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2063),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2295),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2078),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2197),
.B(n_2227),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2295),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2078),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2079),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2236),
.B(n_1766),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2079),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2295),
.Y(n_2650)
);

NAND2xp33_ASAP7_75t_L g2651 ( 
.A(n_2330),
.B(n_1981),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2408),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2476),
.B(n_1447),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2085),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2269),
.B(n_1256),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2127),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2408),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2270),
.B(n_1285),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2471),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2408),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2081),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2411),
.Y(n_2662)
);

INVx3_ASAP7_75t_L g2663 ( 
.A(n_2085),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_2251),
.Y(n_2664)
);

NAND3xp33_ASAP7_75t_L g2665 ( 
.A(n_2235),
.B(n_1678),
.C(n_1675),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2411),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2227),
.B(n_1772),
.Y(n_2667)
);

NAND2xp33_ASAP7_75t_L g2668 ( 
.A(n_2330),
.B(n_1709),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2095),
.Y(n_2669)
);

BUFx10_ASAP7_75t_L g2670 ( 
.A(n_2129),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2081),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2233),
.B(n_1764),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2471),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2238),
.B(n_1627),
.Y(n_2674)
);

INVx8_ASAP7_75t_L g2675 ( 
.A(n_2330),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2083),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2411),
.Y(n_2677)
);

BUFx3_ASAP7_75t_L g2678 ( 
.A(n_2471),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2456),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2233),
.B(n_1711),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2456),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2095),
.A2(n_1766),
.B1(n_1747),
.B2(n_1746),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2083),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2084),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2456),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2457),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2084),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_2271),
.B(n_1291),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2425),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2457),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2276),
.B(n_1299),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2082),
.B(n_1711),
.Y(n_2692)
);

INVx2_ASAP7_75t_SL g2693 ( 
.A(n_2459),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2459),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2457),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2095),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2458),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2458),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2095),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2122),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2122),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_L g2702 ( 
.A(n_2307),
.B(n_1435),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2458),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2082),
.B(n_1711),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2122),
.Y(n_2705)
);

BUFx10_ASAP7_75t_L g2706 ( 
.A(n_2129),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2122),
.Y(n_2707)
);

INVx4_ASAP7_75t_L g2708 ( 
.A(n_2167),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2125),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2092),
.B(n_1803),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2092),
.B(n_1803),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2174),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2174),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2210),
.Y(n_2714)
);

INVx2_ASAP7_75t_SL g2715 ( 
.A(n_2472),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2330),
.A2(n_1747),
.B1(n_1746),
.B2(n_1801),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2096),
.B(n_1803),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2096),
.B(n_1746),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2236),
.B(n_1747),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2210),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2211),
.Y(n_2721)
);

BUFx6f_ASAP7_75t_SL g2722 ( 
.A(n_2278),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2167),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2175),
.Y(n_2724)
);

CKINVDCx6p67_ASAP7_75t_R g2725 ( 
.A(n_2278),
.Y(n_2725)
);

INVx2_ASAP7_75t_SL g2726 ( 
.A(n_2472),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2316),
.B(n_1893),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2395),
.B(n_1440),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2167),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2125),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2125),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2211),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2325),
.B(n_1968),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2125),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2137),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2223),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2223),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2336),
.Y(n_2738)
);

INVx3_ASAP7_75t_L g2739 ( 
.A(n_2137),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2137),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2137),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2358),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2394),
.B(n_2055),
.Y(n_2743)
);

INVx4_ASAP7_75t_L g2744 ( 
.A(n_2167),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2155),
.Y(n_2745)
);

NAND2xp33_ASAP7_75t_L g2746 ( 
.A(n_2330),
.B(n_1719),
.Y(n_2746)
);

INVx4_ASAP7_75t_L g2747 ( 
.A(n_2167),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2155),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_2061),
.B(n_1440),
.Y(n_2749)
);

AND3x2_ASAP7_75t_L g2750 ( 
.A(n_2172),
.B(n_1984),
.C(n_1960),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2155),
.Y(n_2751)
);

INVxp33_ASAP7_75t_L g2752 ( 
.A(n_2462),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2155),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2229),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2106),
.B(n_1730),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2444),
.B(n_2466),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2160),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2160),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2126),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2160),
.Y(n_2760)
);

AND2x6_ASAP7_75t_L g2761 ( 
.A(n_2193),
.B(n_860),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2106),
.B(n_1706),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2247),
.B(n_1952),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2117),
.B(n_1885),
.Y(n_2764)
);

NOR2x1p5_ASAP7_75t_L g2765 ( 
.A(n_2217),
.B(n_1844),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2229),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2240),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2072),
.B(n_1446),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2160),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2175),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2240),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2246),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2246),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2252),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2172),
.Y(n_2775)
);

INVx2_ASAP7_75t_SL g2776 ( 
.A(n_2156),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2109),
.B(n_1446),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2252),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2200),
.B(n_1820),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2471),
.Y(n_2780)
);

NAND2xp33_ASAP7_75t_L g2781 ( 
.A(n_2330),
.B(n_1830),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2254),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_SL g2783 ( 
.A1(n_2305),
.A2(n_1412),
.B1(n_1427),
.B2(n_1394),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2254),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2256),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2256),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2257),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2257),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2167),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2117),
.B(n_2118),
.Y(n_2790)
);

BUFx10_ASAP7_75t_L g2791 ( 
.A(n_2167),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2258),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2258),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2138),
.B(n_1681),
.C(n_1678),
.Y(n_2794)
);

NAND3xp33_ASAP7_75t_L g2795 ( 
.A(n_2422),
.B(n_1681),
.C(n_1886),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2265),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2247),
.B(n_2253),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2253),
.B(n_1952),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2330),
.A2(n_1804),
.B1(n_1808),
.B2(n_1801),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_2434),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2265),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2267),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2205),
.B(n_1863),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2259),
.B(n_1966),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2200),
.B(n_1911),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2267),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2268),
.Y(n_2807)
);

INVx3_ASAP7_75t_L g2808 ( 
.A(n_2161),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2268),
.Y(n_2809)
);

INVxp67_ASAP7_75t_SL g2810 ( 
.A(n_2277),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2272),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2272),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2119),
.A2(n_2397),
.B1(n_2402),
.B2(n_2393),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2205),
.B(n_1937),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2264),
.B(n_1953),
.Y(n_2815)
);

INVx1_ASAP7_75t_SL g2816 ( 
.A(n_2462),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2264),
.B(n_1754),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2239),
.B(n_1745),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_2471),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2281),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2281),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2284),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2284),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2159),
.B(n_1966),
.Y(n_2824)
);

BUFx10_ASAP7_75t_L g2825 ( 
.A(n_2218),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2288),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2159),
.B(n_1858),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2288),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2293),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2118),
.B(n_1858),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2293),
.Y(n_2831)
);

INVx3_ASAP7_75t_L g2832 ( 
.A(n_2161),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2297),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2161),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2161),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2164),
.Y(n_2836)
);

INVx5_ASAP7_75t_L g2837 ( 
.A(n_2218),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2259),
.B(n_2176),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_2176),
.B(n_2037),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2164),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2164),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2297),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2471),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_SL g2844 ( 
.A1(n_2305),
.A2(n_1473),
.B1(n_1429),
.B2(n_1106),
.Y(n_2844)
);

AOI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2218),
.A2(n_1808),
.B1(n_1823),
.B2(n_1804),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2317),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2317),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2119),
.A2(n_1480),
.B1(n_1693),
.B2(n_1775),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2164),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2215),
.Y(n_2850)
);

CKINVDCx11_ASAP7_75t_R g2851 ( 
.A(n_2065),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2215),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2215),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2475),
.B(n_1790),
.Y(n_2854)
);

NAND3xp33_ASAP7_75t_L g2855 ( 
.A(n_2098),
.B(n_1664),
.C(n_1371),
.Y(n_2855)
);

INVx3_ASAP7_75t_L g2856 ( 
.A(n_2215),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2086),
.B(n_1703),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2446),
.A2(n_1808),
.B1(n_1823),
.B2(n_1804),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2221),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2221),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2412),
.B(n_2039),
.Y(n_2861)
);

INVx4_ASAP7_75t_L g2862 ( 
.A(n_2218),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2475),
.B(n_1790),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2221),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2437),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2221),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2255),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2412),
.B(n_1844),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2255),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2255),
.Y(n_2870)
);

BUFx10_ASAP7_75t_L g2871 ( 
.A(n_2218),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2218),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2255),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2285),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2285),
.Y(n_2875)
);

OAI21xp33_ASAP7_75t_SL g2876 ( 
.A1(n_2098),
.A2(n_1671),
.B(n_1802),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2285),
.Y(n_2877)
);

BUFx6f_ASAP7_75t_L g2878 ( 
.A(n_2218),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2285),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2298),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2298),
.Y(n_2881)
);

INVx4_ASAP7_75t_L g2882 ( 
.A(n_2232),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2298),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2468),
.B(n_1855),
.Y(n_2884)
);

BUFx10_ASAP7_75t_L g2885 ( 
.A(n_2195),
.Y(n_2885)
);

INVx3_ASAP7_75t_L g2886 ( 
.A(n_2298),
.Y(n_2886)
);

AOI21x1_ASAP7_75t_L g2887 ( 
.A1(n_2406),
.A2(n_1945),
.B(n_1932),
.Y(n_2887)
);

AOI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_2306),
.A2(n_1829),
.B1(n_1837),
.B2(n_1823),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2306),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2280),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2306),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2225),
.B(n_2087),
.Y(n_2892)
);

BUFx6f_ASAP7_75t_L g2893 ( 
.A(n_2280),
.Y(n_2893)
);

NAND2xp33_ASAP7_75t_L g2894 ( 
.A(n_2199),
.B(n_1776),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2086),
.B(n_1703),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2306),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2338),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2338),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2338),
.Y(n_2899)
);

CKINVDCx5p33_ASAP7_75t_R g2900 ( 
.A(n_2065),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2338),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_SL g2902 ( 
.A(n_2414),
.B(n_1855),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2346),
.Y(n_2903)
);

BUFx3_ASAP7_75t_L g2904 ( 
.A(n_2280),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2346),
.Y(n_2905)
);

INVx2_ASAP7_75t_SL g2906 ( 
.A(n_2260),
.Y(n_2906)
);

BUFx10_ASAP7_75t_L g2907 ( 
.A(n_2201),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2346),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2346),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2351),
.Y(n_2910)
);

BUFx2_ASAP7_75t_L g2911 ( 
.A(n_2219),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2351),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2089),
.B(n_2099),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2351),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2351),
.Y(n_2915)
);

INVx1_ASAP7_75t_SL g2916 ( 
.A(n_2376),
.Y(n_2916)
);

INVx3_ASAP7_75t_L g2917 ( 
.A(n_2386),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2386),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2414),
.B(n_2037),
.Y(n_2919)
);

NAND2xp33_ASAP7_75t_SL g2920 ( 
.A(n_2404),
.B(n_1088),
.Y(n_2920)
);

NOR2x1p5_ASAP7_75t_L g2921 ( 
.A(n_2442),
.B(n_1908),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2446),
.B(n_2039),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2260),
.Y(n_2923)
);

OAI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2537),
.A2(n_2202),
.B(n_2263),
.Y(n_2924)
);

OR2x6_ASAP7_75t_L g2925 ( 
.A(n_2675),
.B(n_2278),
.Y(n_2925)
);

INVx1_ASAP7_75t_SL g2926 ( 
.A(n_2633),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2772),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2525),
.B(n_2266),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2482),
.B(n_2107),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2640),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2772),
.Y(n_2931)
);

BUFx2_ASAP7_75t_L g2932 ( 
.A(n_2742),
.Y(n_2932)
);

CKINVDCx20_ASAP7_75t_R g2933 ( 
.A(n_2851),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2537),
.A2(n_2202),
.B(n_2263),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2772),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2640),
.Y(n_2936)
);

INVx2_ASAP7_75t_SL g2937 ( 
.A(n_2525),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2641),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2641),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_SL g2940 ( 
.A(n_2556),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2622),
.A2(n_2335),
.B(n_2263),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2773),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2643),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2510),
.B(n_2089),
.Y(n_2944)
);

XOR2xp5_ASAP7_75t_L g2945 ( 
.A(n_2783),
.B(n_2376),
.Y(n_2945)
);

INVxp33_ASAP7_75t_L g2946 ( 
.A(n_2512),
.Y(n_2946)
);

CKINVDCx20_ASAP7_75t_R g2947 ( 
.A(n_2900),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2643),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2773),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2837),
.A2(n_2232),
.B(n_2304),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2646),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2646),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2647),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2647),
.Y(n_2954)
);

XOR2xp5_ASAP7_75t_L g2955 ( 
.A(n_2656),
.B(n_1957),
.Y(n_2955)
);

INVxp33_ASAP7_75t_L g2956 ( 
.A(n_2674),
.Y(n_2956)
);

INVx1_ASAP7_75t_SL g2957 ( 
.A(n_2639),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2763),
.B(n_2120),
.Y(n_2958)
);

NAND2x1p5_ASAP7_75t_L g2959 ( 
.A(n_2488),
.B(n_2309),
.Y(n_2959)
);

XOR2xp5_ASAP7_75t_L g2960 ( 
.A(n_2664),
.B(n_1957),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2764),
.B(n_2099),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2649),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2649),
.Y(n_2963)
);

XOR2xp5_ASAP7_75t_L g2964 ( 
.A(n_2738),
.B(n_2111),
.Y(n_2964)
);

NAND2xp33_ASAP7_75t_SL g2965 ( 
.A(n_2494),
.B(n_2477),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2661),
.Y(n_2966)
);

INVx2_ASAP7_75t_SL g2967 ( 
.A(n_2797),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2773),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2536),
.B(n_2548),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2521),
.Y(n_2970)
);

XOR2xp5_ASAP7_75t_L g2971 ( 
.A(n_2800),
.B(n_2111),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2661),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2838),
.B(n_2797),
.Y(n_2973)
);

XNOR2xp5_ASAP7_75t_L g2974 ( 
.A(n_2916),
.B(n_2149),
.Y(n_2974)
);

INVx2_ASAP7_75t_SL g2975 ( 
.A(n_2838),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2782),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2560),
.B(n_2139),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2671),
.Y(n_2978)
);

XNOR2xp5_ASAP7_75t_L g2979 ( 
.A(n_2816),
.B(n_2149),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2671),
.Y(n_2980)
);

XOR2xp5_ASAP7_75t_L g2981 ( 
.A(n_2865),
.B(n_2100),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_SL g2982 ( 
.A(n_2565),
.B(n_2442),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2676),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2676),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2533),
.B(n_2101),
.Y(n_2985)
);

CKINVDCx16_ASAP7_75t_R g2986 ( 
.A(n_2490),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2683),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2683),
.Y(n_2988)
);

OR2x6_ASAP7_75t_L g2989 ( 
.A(n_2675),
.B(n_2278),
.Y(n_2989)
);

NAND2xp33_ASAP7_75t_R g2990 ( 
.A(n_2742),
.B(n_2775),
.Y(n_2990)
);

NAND2x1p5_ASAP7_75t_L g2991 ( 
.A(n_2488),
.B(n_2309),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2684),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2684),
.Y(n_2993)
);

XNOR2x1_ASAP7_75t_L g2994 ( 
.A(n_2484),
.B(n_1381),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2687),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2782),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2687),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2487),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2487),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2837),
.B(n_2232),
.Y(n_3000)
);

AND2x4_ASAP7_75t_L g3001 ( 
.A(n_2632),
.B(n_2446),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2837),
.B(n_2232),
.Y(n_3002)
);

CKINVDCx5p33_ASAP7_75t_R g3003 ( 
.A(n_2546),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2763),
.B(n_2798),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2667),
.B(n_2101),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2491),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2632),
.B(n_2446),
.Y(n_3007)
);

NOR2xp67_ASAP7_75t_L g3008 ( 
.A(n_2559),
.B(n_1908),
.Y(n_3008)
);

CKINVDCx20_ASAP7_75t_R g3009 ( 
.A(n_2725),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2491),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2556),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2782),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2492),
.Y(n_3013)
);

OR2x6_ASAP7_75t_L g3014 ( 
.A(n_2675),
.B(n_2278),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2784),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2672),
.B(n_2105),
.Y(n_3016)
);

CKINVDCx20_ASAP7_75t_R g3017 ( 
.A(n_2725),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2492),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2496),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2759),
.B(n_2105),
.Y(n_3020)
);

OR2x2_ASAP7_75t_L g3021 ( 
.A(n_2541),
.B(n_2145),
.Y(n_3021)
);

NAND2xp33_ASAP7_75t_SL g3022 ( 
.A(n_2494),
.B(n_2304),
.Y(n_3022)
);

XOR2xp5_ASAP7_75t_L g3023 ( 
.A(n_2752),
.B(n_1796),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2496),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2497),
.Y(n_3025)
);

XNOR2xp5_ASAP7_75t_L g3026 ( 
.A(n_2844),
.B(n_2601),
.Y(n_3026)
);

AND2x4_ASAP7_75t_L g3027 ( 
.A(n_2632),
.B(n_2113),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2798),
.B(n_2266),
.Y(n_3028)
);

BUFx3_ASAP7_75t_L g3029 ( 
.A(n_2632),
.Y(n_3029)
);

BUFx3_ASAP7_75t_L g3030 ( 
.A(n_2775),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2561),
.B(n_2113),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2849),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2541),
.B(n_2115),
.Y(n_3033)
);

CKINVDCx20_ASAP7_75t_R g3034 ( 
.A(n_2621),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2759),
.B(n_2115),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2521),
.B(n_2123),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2497),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2508),
.B(n_2123),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2499),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2499),
.Y(n_3040)
);

INVxp33_ASAP7_75t_SL g3041 ( 
.A(n_2884),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_L g3042 ( 
.A(n_2543),
.B(n_2530),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2503),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2489),
.B(n_2124),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2503),
.Y(n_3045)
);

XOR2xp5_ASAP7_75t_L g3046 ( 
.A(n_2911),
.B(n_1819),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_2521),
.B(n_2124),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2516),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2516),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2776),
.B(n_2131),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2837),
.A2(n_2232),
.B(n_2393),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2804),
.B(n_1253),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2529),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2804),
.B(n_1262),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2784),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2489),
.B(n_2131),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2529),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2532),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2532),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2534),
.Y(n_3060)
);

XNOR2x2_ASAP7_75t_L g3061 ( 
.A(n_2855),
.B(n_736),
.Y(n_3061)
);

NOR2xp67_ASAP7_75t_L g3062 ( 
.A(n_2794),
.B(n_1931),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2534),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2776),
.B(n_2648),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2544),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2784),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2648),
.B(n_1315),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2785),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2785),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2544),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2719),
.B(n_2386),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2545),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2489),
.B(n_2140),
.Y(n_3073)
);

CKINVDCx20_ASAP7_75t_R g3074 ( 
.A(n_2911),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2526),
.B(n_2524),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2545),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2547),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2547),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2550),
.Y(n_3079)
);

XNOR2xp5_ASAP7_75t_L g3080 ( 
.A(n_2601),
.B(n_2329),
.Y(n_3080)
);

CKINVDCx20_ASAP7_75t_R g3081 ( 
.A(n_2517),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2550),
.Y(n_3082)
);

AND2x2_ASAP7_75t_SL g3083 ( 
.A(n_2781),
.B(n_2263),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2551),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2719),
.B(n_2386),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2551),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_SL g3087 ( 
.A(n_2818),
.B(n_2442),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2785),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2602),
.B(n_2140),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2553),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2553),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_L g3092 ( 
.A(n_2501),
.B(n_2146),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2554),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2554),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2755),
.B(n_2146),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2563),
.Y(n_3096)
);

INVx1_ASAP7_75t_SL g3097 ( 
.A(n_2674),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2502),
.B(n_2504),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2535),
.B(n_2151),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_SL g3100 ( 
.A(n_2837),
.B(n_2232),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2786),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2563),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2578),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2578),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2583),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2583),
.Y(n_3106)
);

XOR2xp5_ASAP7_75t_L g3107 ( 
.A(n_2618),
.B(n_1819),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2762),
.B(n_2151),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2786),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2586),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2586),
.Y(n_3111)
);

INVx2_ASAP7_75t_SL g3112 ( 
.A(n_2849),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2786),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2599),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2599),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2600),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2718),
.B(n_2153),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2792),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2600),
.Y(n_3119)
);

XOR2xp5_ASAP7_75t_L g3120 ( 
.A(n_2795),
.B(n_1847),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2792),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2509),
.B(n_2153),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2906),
.B(n_1343),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2604),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2906),
.B(n_2923),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2604),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2605),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_2556),
.B(n_2154),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2605),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2606),
.Y(n_3130)
);

OR2x6_ASAP7_75t_L g3131 ( 
.A(n_2675),
.B(n_2329),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_SL g3132 ( 
.A(n_2556),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2792),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_SL g3134 ( 
.A(n_2722),
.B(n_2442),
.Y(n_3134)
);

AND2x2_ASAP7_75t_SL g3135 ( 
.A(n_2555),
.B(n_2335),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2606),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2608),
.Y(n_3137)
);

AND2x2_ASAP7_75t_L g3138 ( 
.A(n_2923),
.B(n_2514),
.Y(n_3138)
);

INVxp33_ASAP7_75t_L g3139 ( 
.A(n_2779),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2514),
.B(n_1422),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2528),
.B(n_1453),
.Y(n_3141)
);

AND2x4_ASAP7_75t_L g3142 ( 
.A(n_2521),
.B(n_2154),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2793),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2608),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_2572),
.B(n_2162),
.Y(n_3145)
);

CKINVDCx20_ASAP7_75t_R g3146 ( 
.A(n_2920),
.Y(n_3146)
);

AND2x4_ASAP7_75t_L g3147 ( 
.A(n_2572),
.B(n_2162),
.Y(n_3147)
);

CKINVDCx16_ASAP7_75t_R g3148 ( 
.A(n_2722),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2793),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2611),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2611),
.Y(n_3151)
);

INVx2_ASAP7_75t_SL g3152 ( 
.A(n_2849),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2614),
.Y(n_3153)
);

XOR2x2_ASAP7_75t_L g3154 ( 
.A(n_2892),
.B(n_1417),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2728),
.B(n_2749),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2614),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2535),
.B(n_2163),
.Y(n_3157)
);

BUFx6f_ASAP7_75t_L g3158 ( 
.A(n_2494),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2619),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2854),
.B(n_2163),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2619),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2623),
.Y(n_3162)
);

AND2x4_ASAP7_75t_L g3163 ( 
.A(n_2572),
.B(n_2165),
.Y(n_3163)
);

BUFx8_ASAP7_75t_L g3164 ( 
.A(n_2722),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2854),
.B(n_2165),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2623),
.Y(n_3166)
);

AOI21x1_ASAP7_75t_L g3167 ( 
.A1(n_2519),
.A2(n_2402),
.B(n_2397),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2624),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_2863),
.B(n_2171),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2598),
.B(n_2171),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2624),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2631),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2631),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2637),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2637),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_2863),
.B(n_2173),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2638),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2625),
.B(n_2173),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2626),
.B(n_2178),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2793),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2638),
.Y(n_3181)
);

XNOR2xp5_ASAP7_75t_L g3182 ( 
.A(n_2765),
.B(n_2921),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2756),
.B(n_2178),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2528),
.B(n_2574),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_2850),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2801),
.Y(n_3186)
);

XOR2xp5_ASAP7_75t_L g3187 ( 
.A(n_2665),
.B(n_1847),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2714),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2714),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2801),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2876),
.B(n_2181),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2876),
.B(n_2181),
.Y(n_3192)
);

NOR2xp67_ASAP7_75t_L g3193 ( 
.A(n_2805),
.B(n_1931),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_2750),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2720),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2574),
.B(n_1366),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2720),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2721),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2721),
.Y(n_3199)
);

XOR2xp5_ASAP7_75t_L g3200 ( 
.A(n_2634),
.B(n_1898),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2732),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2732),
.Y(n_3202)
);

XOR2xp5_ASAP7_75t_L g3203 ( 
.A(n_2636),
.B(n_1898),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2736),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2736),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2644),
.B(n_2182),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2737),
.Y(n_3207)
);

XNOR2xp5_ASAP7_75t_L g3208 ( 
.A(n_2765),
.B(n_2329),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2790),
.B(n_2182),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2737),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2801),
.Y(n_3211)
);

XOR2xp5_ASAP7_75t_L g3212 ( 
.A(n_2653),
.B(n_1897),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_2580),
.B(n_1879),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2754),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_2593),
.B(n_2335),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2754),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2766),
.Y(n_3217)
);

OAI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_2505),
.A2(n_2344),
.B(n_2335),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_2593),
.B(n_2344),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2580),
.B(n_2188),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2766),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2590),
.B(n_2344),
.Y(n_3222)
);

AND2x4_ASAP7_75t_L g3223 ( 
.A(n_2572),
.B(n_2309),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2485),
.B(n_2188),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2807),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2767),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2767),
.Y(n_3227)
);

CKINVDCx5p33_ASAP7_75t_R g3228 ( 
.A(n_2722),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2771),
.Y(n_3229)
);

AND2x6_ASAP7_75t_L g3230 ( 
.A(n_2615),
.B(n_2723),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_2691),
.B(n_2189),
.Y(n_3231)
);

XNOR2x2_ASAP7_75t_L g3232 ( 
.A(n_2573),
.B(n_919),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_2702),
.B(n_2562),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_L g3234 ( 
.A(n_2506),
.B(n_2189),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2771),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2774),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2774),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2778),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2778),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2807),
.Y(n_3240)
);

NAND2xp33_ASAP7_75t_R g3241 ( 
.A(n_2629),
.B(n_2329),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2787),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2787),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2837),
.A2(n_2241),
.B(n_2274),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2788),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2807),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_2590),
.B(n_2344),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_L g3248 ( 
.A(n_2727),
.B(n_2190),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2788),
.Y(n_3249)
);

XOR2x2_ASAP7_75t_L g3250 ( 
.A(n_2609),
.B(n_1444),
.Y(n_3250)
);

NOR2xp67_ASAP7_75t_L g3251 ( 
.A(n_2576),
.B(n_1936),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2627),
.B(n_2190),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2627),
.B(n_2348),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2796),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2635),
.B(n_2348),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2635),
.B(n_2348),
.Y(n_3256)
);

CKINVDCx20_ASAP7_75t_R g3257 ( 
.A(n_2922),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2689),
.B(n_2693),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2796),
.Y(n_3259)
);

XOR2x2_ASAP7_75t_L g3260 ( 
.A(n_2733),
.B(n_2743),
.Y(n_3260)
);

XNOR2xp5_ASAP7_75t_L g3261 ( 
.A(n_2921),
.B(n_2515),
.Y(n_3261)
);

AND2x4_ASAP7_75t_L g3262 ( 
.A(n_2592),
.B(n_2191),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2689),
.B(n_2348),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2802),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2802),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_2693),
.B(n_1879),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2811),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2668),
.A2(n_2274),
.B(n_1817),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_2694),
.B(n_2191),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_2694),
.B(n_1936),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_2715),
.B(n_2329),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_2715),
.B(n_1406),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2806),
.Y(n_3273)
);

CKINVDCx20_ASAP7_75t_R g3274 ( 
.A(n_2861),
.Y(n_3274)
);

INVxp33_ASAP7_75t_SL g3275 ( 
.A(n_2555),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_2850),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2806),
.Y(n_3277)
);

INVxp33_ASAP7_75t_SL g3278 ( 
.A(n_2848),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2809),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2726),
.B(n_2403),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2809),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2812),
.Y(n_3282)
);

NOR2xp67_ASAP7_75t_L g3283 ( 
.A(n_2726),
.B(n_1750),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2811),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2811),
.Y(n_3285)
);

BUFx3_ASAP7_75t_L g3286 ( 
.A(n_2850),
.Y(n_3286)
);

INVxp33_ASAP7_75t_L g3287 ( 
.A(n_2655),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2812),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2820),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_2592),
.B(n_2403),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2820),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2821),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2824),
.B(n_2403),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_2830),
.B(n_2403),
.Y(n_3294)
);

NOR2xp67_ASAP7_75t_L g3295 ( 
.A(n_2531),
.B(n_1750),
.Y(n_3295)
);

OAI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_2539),
.A2(n_2274),
.B(n_2424),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2821),
.Y(n_3297)
);

AND2x4_ASAP7_75t_L g3298 ( 
.A(n_2592),
.B(n_2628),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2682),
.B(n_2274),
.Y(n_3299)
);

INVxp67_ASAP7_75t_SL g3300 ( 
.A(n_2494),
.Y(n_3300)
);

NOR2xp33_ASAP7_75t_L g3301 ( 
.A(n_2768),
.B(n_2416),
.Y(n_3301)
);

XOR2xp5_ASAP7_75t_L g3302 ( 
.A(n_2658),
.B(n_2219),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_2688),
.B(n_1789),
.Y(n_3303)
);

CKINVDCx20_ASAP7_75t_R g3304 ( 
.A(n_2868),
.Y(n_3304)
);

INVxp67_ASAP7_75t_L g3305 ( 
.A(n_2777),
.Y(n_3305)
);

INVx2_ASAP7_75t_SL g3306 ( 
.A(n_2853),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2710),
.B(n_2416),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2822),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2803),
.B(n_1641),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2822),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_SL g3311 ( 
.A(n_2853),
.B(n_1705),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2567),
.A2(n_2427),
.B(n_2424),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2829),
.Y(n_3313)
);

INVx1_ASAP7_75t_SL g3314 ( 
.A(n_2814),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2823),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2829),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2833),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2823),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2823),
.Y(n_3319)
);

XNOR2xp5_ASAP7_75t_L g3320 ( 
.A(n_2515),
.B(n_2219),
.Y(n_3320)
);

HB1xp67_ASAP7_75t_L g3321 ( 
.A(n_2913),
.Y(n_3321)
);

AND2x2_ASAP7_75t_L g3322 ( 
.A(n_2815),
.B(n_1684),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2833),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2842),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_2827),
.B(n_2420),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_2826),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2826),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2842),
.Y(n_3328)
);

NAND2xp33_ASAP7_75t_R g3329 ( 
.A(n_2483),
.B(n_2486),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_2592),
.B(n_1829),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2826),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2846),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_2853),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2846),
.Y(n_3334)
);

INVxp67_ASAP7_75t_SL g3335 ( 
.A(n_2494),
.Y(n_3335)
);

XNOR2xp5_ASAP7_75t_L g3336 ( 
.A(n_2902),
.B(n_2219),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_2628),
.B(n_1829),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2828),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_2493),
.B(n_1837),
.Y(n_3339)
);

INVx4_ASAP7_75t_L g3340 ( 
.A(n_2675),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_2746),
.A2(n_1817),
.B(n_1814),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2828),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2828),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2711),
.B(n_2420),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2831),
.Y(n_3345)
);

INVx2_ASAP7_75t_SL g3346 ( 
.A(n_2867),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2717),
.B(n_2421),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2696),
.B(n_2421),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2831),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2831),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_2493),
.B(n_1837),
.Y(n_3351)
);

OAI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2581),
.A2(n_2430),
.B(n_2427),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2847),
.Y(n_3353)
);

CKINVDCx20_ASAP7_75t_R g3354 ( 
.A(n_2919),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2847),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_L g3356 ( 
.A(n_2696),
.B(n_2430),
.Y(n_3356)
);

XOR2xp5_ASAP7_75t_L g3357 ( 
.A(n_2839),
.B(n_2381),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2847),
.Y(n_3358)
);

CKINVDCx20_ASAP7_75t_R g3359 ( 
.A(n_2589),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_2700),
.B(n_2431),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_2716),
.B(n_1802),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2867),
.Y(n_3362)
);

INVxp33_ASAP7_75t_L g3363 ( 
.A(n_2594),
.Y(n_3363)
);

OAI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_2585),
.A2(n_2438),
.B(n_2431),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_2591),
.A2(n_2440),
.B(n_2438),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_2628),
.B(n_1865),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_SL g3367 ( 
.A(n_2867),
.B(n_1705),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_2628),
.B(n_1865),
.Y(n_3368)
);

AND2x6_ASAP7_75t_L g3369 ( 
.A(n_2615),
.B(n_2723),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_2700),
.B(n_2440),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2712),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_2873),
.Y(n_3372)
);

NAND2xp33_ASAP7_75t_SL g3373 ( 
.A(n_2494),
.B(n_1088),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_2873),
.Y(n_3374)
);

OAI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_2595),
.A2(n_2445),
.B(n_2441),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_2493),
.B(n_1865),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2873),
.Y(n_3377)
);

INVxp67_ASAP7_75t_SL g3378 ( 
.A(n_2558),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2874),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2874),
.Y(n_3380)
);

OAI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_2612),
.A2(n_2445),
.B(n_2441),
.Y(n_3381)
);

CKINVDCx5p33_ASAP7_75t_R g3382 ( 
.A(n_2542),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_2874),
.B(n_1834),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2875),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2875),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2875),
.Y(n_3386)
);

XOR2xp5_ASAP7_75t_L g3387 ( 
.A(n_2858),
.B(n_2381),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2712),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2889),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_3001),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2930),
.Y(n_3391)
);

AND2x2_ASAP7_75t_L g3392 ( 
.A(n_3067),
.B(n_2817),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_3155),
.B(n_2527),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2936),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2927),
.Y(n_3395)
);

INVx3_ASAP7_75t_L g3396 ( 
.A(n_3001),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3052),
.B(n_1834),
.Y(n_3397)
);

BUFx6f_ASAP7_75t_SL g3398 ( 
.A(n_3030),
.Y(n_3398)
);

BUFx3_ASAP7_75t_L g3399 ( 
.A(n_3030),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2938),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2969),
.B(n_2680),
.Y(n_3401)
);

HB1xp67_ASAP7_75t_L g3402 ( 
.A(n_2932),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2969),
.B(n_2692),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3155),
.B(n_3031),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2927),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2931),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3031),
.B(n_3231),
.Y(n_3407)
);

A2O1A1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_3233),
.A2(n_2705),
.B(n_2707),
.C(n_2701),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3231),
.B(n_3004),
.Y(n_3409)
);

AOI22xp33_ASAP7_75t_L g3410 ( 
.A1(n_3233),
.A2(n_2891),
.B1(n_2918),
.B2(n_2889),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_3158),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2931),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3054),
.B(n_1835),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2935),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3178),
.B(n_2704),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2939),
.Y(n_3416)
);

INVx2_ASAP7_75t_SL g3417 ( 
.A(n_2926),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3178),
.B(n_2523),
.Y(n_3418)
);

HB1xp67_ASAP7_75t_L g3419 ( 
.A(n_2990),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2973),
.B(n_2523),
.Y(n_3420)
);

BUFx3_ASAP7_75t_L g3421 ( 
.A(n_3034),
.Y(n_3421)
);

CKINVDCx16_ASAP7_75t_R g3422 ( 
.A(n_2986),
.Y(n_3422)
);

NOR2xp33_ASAP7_75t_L g3423 ( 
.A(n_3139),
.B(n_2701),
.Y(n_3423)
);

NOR2x1p5_ASAP7_75t_L g3424 ( 
.A(n_3003),
.B(n_1761),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2973),
.B(n_2538),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2943),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_3158),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2948),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3278),
.A2(n_2891),
.B1(n_2918),
.B2(n_2889),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2935),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_3298),
.B(n_2527),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3139),
.B(n_2705),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3278),
.A2(n_2918),
.B1(n_2891),
.B2(n_2538),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3038),
.B(n_2540),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3275),
.A2(n_2540),
.B1(n_2552),
.B2(n_2549),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3038),
.B(n_2549),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3275),
.A2(n_2552),
.B1(n_2564),
.B2(n_2557),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2942),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3089),
.B(n_2557),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_2942),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2951),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2952),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2953),
.Y(n_3443)
);

INVxp67_ASAP7_75t_L g3444 ( 
.A(n_2990),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_3298),
.B(n_2527),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3089),
.B(n_2564),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_2947),
.Y(n_3447)
);

BUFx8_ASAP7_75t_L g3448 ( 
.A(n_2940),
.Y(n_3448)
);

AOI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_3042),
.A2(n_2730),
.B1(n_2731),
.B2(n_2566),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3298),
.B(n_2527),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_2949),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2954),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_2962),
.Y(n_3453)
);

BUFx3_ASAP7_75t_L g3454 ( 
.A(n_3034),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_2949),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_3041),
.B(n_2707),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3042),
.B(n_2575),
.Y(n_3457)
);

OR2x6_ASAP7_75t_L g3458 ( 
.A(n_2925),
.B(n_2615),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3321),
.B(n_2566),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3044),
.A2(n_2731),
.B1(n_2734),
.B2(n_2730),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_2961),
.B(n_2734),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_2957),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3028),
.B(n_2735),
.Y(n_3463)
);

AND2x6_ASAP7_75t_SL g3464 ( 
.A(n_3270),
.B(n_1835),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2963),
.Y(n_3465)
);

INVxp67_ASAP7_75t_L g3466 ( 
.A(n_3021),
.Y(n_3466)
);

BUFx6f_ASAP7_75t_L g3467 ( 
.A(n_3158),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_2970),
.B(n_2575),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_2968),
.Y(n_3469)
);

NAND2x1_ASAP7_75t_L g3470 ( 
.A(n_3340),
.B(n_2575),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3028),
.B(n_2735),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2966),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_2968),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3123),
.B(n_1851),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_3041),
.B(n_2859),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3005),
.B(n_2740),
.Y(n_3476)
);

INVx4_ASAP7_75t_L g3477 ( 
.A(n_3158),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2956),
.B(n_2929),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2928),
.B(n_2740),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2928),
.B(n_2741),
.Y(n_3480)
);

NOR3xp33_ASAP7_75t_L g3481 ( 
.A(n_3270),
.B(n_2915),
.C(n_2912),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_2976),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_2970),
.B(n_2575),
.Y(n_3483)
);

NAND3xp33_ASAP7_75t_L g3484 ( 
.A(n_2929),
.B(n_2977),
.C(n_2994),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_2976),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_2956),
.B(n_2859),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_2937),
.B(n_2741),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_2996),
.Y(n_3488)
);

INVxp67_ASAP7_75t_L g3489 ( 
.A(n_3140),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2937),
.B(n_2745),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_2967),
.B(n_2745),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_2970),
.B(n_2579),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2967),
.B(n_2748),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3097),
.B(n_2860),
.Y(n_3494)
);

OAI22xp5_ASAP7_75t_SL g3495 ( 
.A1(n_2945),
.A2(n_1106),
.B1(n_1229),
.B2(n_1189),
.Y(n_3495)
);

INVx8_ASAP7_75t_L g3496 ( 
.A(n_3001),
.Y(n_3496)
);

INVxp67_ASAP7_75t_L g3497 ( 
.A(n_3141),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3196),
.B(n_1851),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_2975),
.B(n_2748),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3373),
.A2(n_2758),
.B1(n_2760),
.B2(n_2753),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2972),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_2977),
.B(n_2860),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3044),
.B(n_2579),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_2996),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_2975),
.B(n_2753),
.Y(n_3505)
);

NAND2xp33_ASAP7_75t_L g3506 ( 
.A(n_3230),
.B(n_2558),
.Y(n_3506)
);

OAI22xp5_ASAP7_75t_L g3507 ( 
.A1(n_3056),
.A2(n_2904),
.B1(n_2890),
.B2(n_2558),
.Y(n_3507)
);

INVxp67_ASAP7_75t_L g3508 ( 
.A(n_3272),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_2958),
.B(n_1854),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3016),
.B(n_2758),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3095),
.B(n_3108),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_SL g3512 ( 
.A(n_3056),
.B(n_2579),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2978),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3206),
.B(n_2760),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3209),
.B(n_2834),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3064),
.B(n_3160),
.Y(n_3516)
);

INVxp33_ASAP7_75t_SL g3517 ( 
.A(n_2955),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3073),
.B(n_2579),
.Y(n_3518)
);

INVxp33_ASAP7_75t_L g3519 ( 
.A(n_2946),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3160),
.B(n_2834),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_3073),
.B(n_2596),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3012),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3012),
.Y(n_3523)
);

NOR3x1_ASAP7_75t_L g3524 ( 
.A(n_3303),
.B(n_863),
.C(n_861),
.Y(n_3524)
);

BUFx8_ASAP7_75t_L g3525 ( 
.A(n_2940),
.Y(n_3525)
);

OAI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_2982),
.A2(n_3087),
.B1(n_3287),
.B2(n_3382),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3165),
.B(n_2836),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3033),
.B(n_2864),
.Y(n_3528)
);

OAI22xp33_ASAP7_75t_L g3529 ( 
.A1(n_3287),
.A2(n_2858),
.B1(n_2841),
.B2(n_2836),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3165),
.B(n_2841),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3169),
.B(n_2896),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3033),
.B(n_2864),
.Y(n_3532)
);

INVx4_ASAP7_75t_L g3533 ( 
.A(n_3007),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3015),
.Y(n_3534)
);

AOI22xp33_ASAP7_75t_L g3535 ( 
.A1(n_3071),
.A2(n_2908),
.B1(n_2910),
.B2(n_2896),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_3294),
.B(n_2596),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3071),
.A2(n_2910),
.B1(n_2908),
.B2(n_2869),
.Y(n_3537)
);

INVxp67_ASAP7_75t_SL g3538 ( 
.A(n_3329),
.Y(n_3538)
);

OR2x2_ASAP7_75t_L g3539 ( 
.A(n_3154),
.B(n_2994),
.Y(n_3539)
);

OAI221xp5_ASAP7_75t_L g3540 ( 
.A1(n_3154),
.A2(n_2888),
.B1(n_2616),
.B2(n_2845),
.C(n_2799),
.Y(n_3540)
);

A2O1A1Ixp33_ASAP7_75t_L g3541 ( 
.A1(n_3191),
.A2(n_2869),
.B(n_2870),
.C(n_2866),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3294),
.B(n_2596),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3290),
.B(n_2596),
.Y(n_3543)
);

INVx5_ASAP7_75t_L g3544 ( 
.A(n_3230),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3015),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_2980),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3169),
.B(n_2866),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3085),
.A2(n_2877),
.B1(n_2879),
.B2(n_2870),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3176),
.B(n_2877),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2983),
.Y(n_3550)
);

INVx2_ASAP7_75t_SL g3551 ( 
.A(n_3213),
.Y(n_3551)
);

AOI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3085),
.A2(n_2880),
.B1(n_2881),
.B2(n_2879),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_SL g3553 ( 
.A(n_3290),
.B(n_2708),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3290),
.B(n_3262),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3176),
.B(n_2880),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_3309),
.B(n_2912),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3262),
.B(n_2708),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_3262),
.B(n_2708),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_2984),
.Y(n_3559)
);

INVx2_ASAP7_75t_SL g3560 ( 
.A(n_3266),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_2987),
.Y(n_3561)
);

BUFx2_ASAP7_75t_L g3562 ( 
.A(n_2947),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3269),
.B(n_2881),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3269),
.B(n_2883),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3280),
.B(n_2883),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3280),
.B(n_2899),
.Y(n_3566)
);

AND2x4_ASAP7_75t_L g3567 ( 
.A(n_3029),
.B(n_2899),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_2988),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_2992),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_2985),
.B(n_2901),
.Y(n_3570)
);

AND2x4_ASAP7_75t_L g3571 ( 
.A(n_3029),
.B(n_2901),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_SL g3572 ( 
.A(n_3007),
.B(n_3075),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_2993),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_SL g3574 ( 
.A(n_3032),
.B(n_2708),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_3293),
.A2(n_3192),
.B1(n_3191),
.B2(n_3361),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3322),
.B(n_1854),
.Y(n_3576)
);

BUFx12f_ASAP7_75t_SL g3577 ( 
.A(n_2925),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3099),
.B(n_2905),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2995),
.Y(n_3579)
);

NOR2xp67_ASAP7_75t_L g3580 ( 
.A(n_3003),
.B(n_1761),
.Y(n_3580)
);

BUFx3_ASAP7_75t_L g3581 ( 
.A(n_3164),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3099),
.B(n_2905),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3055),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3157),
.B(n_1860),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_3032),
.B(n_2744),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3157),
.B(n_2915),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3179),
.B(n_2630),
.Y(n_3587)
);

AOI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3373),
.A2(n_3098),
.B1(n_3293),
.B2(n_3260),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_2946),
.B(n_2630),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_2997),
.Y(n_3590)
);

INVx2_ASAP7_75t_SL g3591 ( 
.A(n_3260),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_SL g3592 ( 
.A(n_3112),
.B(n_2744),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3192),
.A2(n_2898),
.B(n_2903),
.C(n_2897),
.Y(n_3593)
);

OAI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3224),
.A2(n_2904),
.B1(n_2890),
.B2(n_2558),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3112),
.B(n_2744),
.Y(n_3595)
);

INVxp67_ASAP7_75t_L g3596 ( 
.A(n_3075),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3055),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2998),
.Y(n_3598)
);

AOI22xp33_ASAP7_75t_L g3599 ( 
.A1(n_3007),
.A2(n_2630),
.B1(n_2663),
.B2(n_2654),
.Y(n_3599)
);

AND2x2_ASAP7_75t_SL g3600 ( 
.A(n_3135),
.B(n_2615),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3179),
.B(n_2630),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3258),
.B(n_2654),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3066),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3125),
.B(n_2654),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_2999),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3006),
.Y(n_3606)
);

INVx3_ASAP7_75t_L g3607 ( 
.A(n_3223),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3138),
.B(n_2654),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3268),
.A2(n_2747),
.B(n_2744),
.Y(n_3609)
);

NAND2xp33_ASAP7_75t_SL g3610 ( 
.A(n_2940),
.B(n_2558),
.Y(n_3610)
);

AOI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3098),
.A2(n_2669),
.B1(n_2699),
.B2(n_2663),
.Y(n_3611)
);

AOI22xp33_ASAP7_75t_L g3612 ( 
.A1(n_3061),
.A2(n_2669),
.B1(n_2699),
.B2(n_2663),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3184),
.B(n_2663),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3170),
.B(n_2669),
.Y(n_3614)
);

OAI21xp33_ASAP7_75t_L g3615 ( 
.A1(n_3183),
.A2(n_1229),
.B(n_1189),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_3305),
.B(n_2669),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_SL g3617 ( 
.A(n_2933),
.B(n_2381),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3061),
.A2(n_2709),
.B1(n_2739),
.B2(n_2699),
.Y(n_3618)
);

INVx2_ASAP7_75t_SL g3619 ( 
.A(n_3232),
.Y(n_3619)
);

NAND3xp33_ASAP7_75t_L g3620 ( 
.A(n_3183),
.B(n_1944),
.C(n_1839),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3170),
.B(n_2699),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3010),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_SL g3623 ( 
.A(n_3152),
.B(n_2747),
.Y(n_3623)
);

BUFx3_ASAP7_75t_L g3624 ( 
.A(n_3164),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3066),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3248),
.B(n_2709),
.Y(n_3626)
);

AOI22xp5_ASAP7_75t_L g3627 ( 
.A1(n_3271),
.A2(n_2739),
.B1(n_2751),
.B2(n_2709),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3248),
.B(n_2709),
.Y(n_3628)
);

HB1xp67_ASAP7_75t_L g3629 ( 
.A(n_3027),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_3314),
.B(n_2739),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3234),
.B(n_2739),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3234),
.B(n_2751),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3117),
.B(n_2751),
.Y(n_3633)
);

NOR2x1p5_ASAP7_75t_L g3634 ( 
.A(n_3382),
.B(n_1770),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3027),
.B(n_2751),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3068),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3224),
.B(n_2757),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3068),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3069),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3383),
.B(n_2757),
.Y(n_3640)
);

INVx2_ASAP7_75t_SL g3641 ( 
.A(n_3232),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_L g3642 ( 
.A(n_2974),
.B(n_2757),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3383),
.B(n_2757),
.Y(n_3643)
);

NOR3xp33_ASAP7_75t_L g3644 ( 
.A(n_3271),
.B(n_2808),
.C(n_2769),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3013),
.Y(n_3645)
);

NOR2xp67_ASAP7_75t_L g3646 ( 
.A(n_3283),
.B(n_1770),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3152),
.B(n_2747),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3244),
.A2(n_2862),
.B(n_2747),
.Y(n_3648)
);

AOI221xp5_ASAP7_75t_L g3649 ( 
.A1(n_2979),
.A2(n_1194),
.B1(n_919),
.B2(n_794),
.C(n_850),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_L g3650 ( 
.A(n_3220),
.B(n_2808),
.Y(n_3650)
);

INVx4_ASAP7_75t_L g3651 ( 
.A(n_3223),
.Y(n_3651)
);

AND2x6_ASAP7_75t_SL g3652 ( 
.A(n_2925),
.B(n_1860),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_SL g3653 ( 
.A(n_3185),
.B(n_2862),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3252),
.B(n_2769),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3018),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3092),
.B(n_2769),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_2933),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3019),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3128),
.B(n_2769),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3024),
.Y(n_3660)
);

AND2x4_ASAP7_75t_L g3661 ( 
.A(n_3027),
.B(n_2808),
.Y(n_3661)
);

BUFx3_ASAP7_75t_L g3662 ( 
.A(n_3164),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_3230),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3092),
.B(n_3122),
.Y(n_3664)
);

BUFx2_ASAP7_75t_L g3665 ( 
.A(n_3074),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3185),
.B(n_2862),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_SL g3667 ( 
.A(n_3306),
.B(n_2862),
.Y(n_3667)
);

INVx2_ASAP7_75t_SL g3668 ( 
.A(n_3250),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3025),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3276),
.A2(n_2808),
.B1(n_2835),
.B2(n_2832),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3069),
.Y(n_3671)
);

O2A1O1Ixp5_ASAP7_75t_L g3672 ( 
.A1(n_2965),
.A2(n_2813),
.B(n_2713),
.C(n_2724),
.Y(n_3672)
);

NAND2xp33_ASAP7_75t_L g3673 ( 
.A(n_3230),
.B(n_2558),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3022),
.A2(n_2651),
.B(n_2882),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3088),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3088),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3101),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_3306),
.B(n_2615),
.Y(n_3678)
);

NOR2xp67_ASAP7_75t_L g3679 ( 
.A(n_3193),
.B(n_1780),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3128),
.B(n_2832),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3037),
.B(n_2832),
.Y(n_3681)
);

BUFx6f_ASAP7_75t_L g3682 ( 
.A(n_3230),
.Y(n_3682)
);

INVx2_ASAP7_75t_SL g3683 ( 
.A(n_3250),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3122),
.B(n_1870),
.Y(n_3684)
);

INVx4_ASAP7_75t_L g3685 ( 
.A(n_3223),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3039),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3040),
.B(n_2832),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3333),
.B(n_2615),
.Y(n_3688)
);

HB1xp67_ASAP7_75t_L g3689 ( 
.A(n_3020),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3043),
.B(n_2835),
.Y(n_3690)
);

OR2x6_ASAP7_75t_L g3691 ( 
.A(n_2925),
.B(n_2723),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3045),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3333),
.B(n_2723),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3101),
.Y(n_3694)
);

AND2x2_ASAP7_75t_SL g3695 ( 
.A(n_3135),
.B(n_2723),
.Y(n_3695)
);

OAI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_3363),
.A2(n_2914),
.B1(n_2917),
.B2(n_2909),
.Y(n_3696)
);

BUFx2_ASAP7_75t_L g3697 ( 
.A(n_3074),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3276),
.A2(n_2835),
.B1(n_2852),
.B2(n_2840),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3035),
.B(n_2835),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3048),
.B(n_2840),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3049),
.B(n_2840),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3053),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3109),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3057),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3050),
.B(n_2840),
.Y(n_3705)
);

INVxp67_ASAP7_75t_L g3706 ( 
.A(n_2960),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3058),
.B(n_2852),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3059),
.B(n_2852),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3346),
.B(n_2723),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_3346),
.B(n_2729),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3374),
.B(n_2729),
.Y(n_3711)
);

BUFx3_ASAP7_75t_L g3712 ( 
.A(n_3009),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3109),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3113),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3363),
.B(n_1870),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3060),
.B(n_2852),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_SL g3717 ( 
.A(n_3286),
.B(n_2886),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3146),
.B(n_2856),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3063),
.B(n_2856),
.Y(n_3719)
);

INVx2_ASAP7_75t_SL g3720 ( 
.A(n_3194),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_L g3721 ( 
.A1(n_3286),
.A2(n_2856),
.B1(n_2897),
.B2(n_2886),
.Y(n_3721)
);

INVx2_ASAP7_75t_SL g3722 ( 
.A(n_3274),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3065),
.B(n_2856),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_3146),
.B(n_2886),
.Y(n_3724)
);

AOI22xp33_ASAP7_75t_L g3725 ( 
.A1(n_3339),
.A2(n_2886),
.B1(n_2898),
.B2(n_2897),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3113),
.Y(n_3726)
);

O2A1O1Ixp33_ASAP7_75t_L g3727 ( 
.A1(n_2944),
.A2(n_2894),
.B(n_2895),
.C(n_2857),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3118),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3118),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3070),
.B(n_2897),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3072),
.B(n_2898),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3076),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3230),
.Y(n_3733)
);

OAI221xp5_ASAP7_75t_L g3734 ( 
.A1(n_3026),
.A2(n_794),
.B1(n_803),
.B2(n_761),
.C(n_750),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_3011),
.B(n_2898),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3121),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3011),
.B(n_1793),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3008),
.B(n_1794),
.Y(n_3738)
);

INVx2_ASAP7_75t_SL g3739 ( 
.A(n_3274),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3121),
.Y(n_3740)
);

INVx4_ASAP7_75t_L g3741 ( 
.A(n_3369),
.Y(n_3741)
);

NAND2xp33_ASAP7_75t_L g3742 ( 
.A(n_3369),
.B(n_2613),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3077),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3022),
.A2(n_2882),
.B(n_2613),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3304),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3078),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3133),
.Y(n_3747)
);

OAI22xp5_ASAP7_75t_SL g3748 ( 
.A1(n_2964),
.A2(n_1813),
.B1(n_1822),
.B2(n_1807),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3079),
.B(n_2903),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_SL g3750 ( 
.A(n_3374),
.B(n_2729),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3339),
.A2(n_2903),
.B1(n_2914),
.B2(n_2909),
.Y(n_3751)
);

NAND3xp33_ASAP7_75t_L g3752 ( 
.A(n_3301),
.B(n_1944),
.C(n_1839),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3133),
.Y(n_3753)
);

NOR2xp33_ASAP7_75t_L g3754 ( 
.A(n_3082),
.B(n_3084),
.Y(n_3754)
);

AND2x6_ASAP7_75t_L g3755 ( 
.A(n_3215),
.B(n_2729),
.Y(n_3755)
);

BUFx5_ASAP7_75t_L g3756 ( 
.A(n_3369),
.Y(n_3756)
);

NOR2xp33_ASAP7_75t_L g3757 ( 
.A(n_3086),
.B(n_2903),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3090),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3091),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3093),
.B(n_2909),
.Y(n_3760)
);

OR2x2_ASAP7_75t_L g3761 ( 
.A(n_3212),
.B(n_2712),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3094),
.B(n_2909),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3096),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3102),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3103),
.B(n_2914),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3104),
.B(n_2914),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3143),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3105),
.B(n_2917),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3143),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3106),
.B(n_2917),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3149),
.Y(n_3771)
);

INVxp67_ASAP7_75t_L g3772 ( 
.A(n_3301),
.Y(n_3772)
);

BUFx2_ASAP7_75t_L g3773 ( 
.A(n_3257),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3304),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_SL g3775 ( 
.A(n_3134),
.B(n_2381),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3110),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3111),
.B(n_2917),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3114),
.B(n_2713),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3115),
.B(n_2713),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3116),
.B(n_2890),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3036),
.B(n_2729),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3351),
.A2(n_2761),
.B1(n_2770),
.B2(n_2724),
.Y(n_3782)
);

NOR2xp33_ASAP7_75t_L g3783 ( 
.A(n_3119),
.B(n_2724),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_SL g3784 ( 
.A(n_3036),
.B(n_2729),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3124),
.B(n_2904),
.Y(n_3785)
);

INVxp33_ASAP7_75t_SL g3786 ( 
.A(n_3023),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3126),
.B(n_2770),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_SL g3788 ( 
.A(n_3484),
.B(n_3251),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3506),
.A2(n_3335),
.B(n_3300),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3395),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3673),
.A2(n_3742),
.B(n_3609),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3407),
.B(n_3127),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3404),
.B(n_3409),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3674),
.A2(n_3378),
.B(n_3299),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3539),
.B(n_3257),
.Y(n_3795)
);

BUFx3_ASAP7_75t_L g3796 ( 
.A(n_3399),
.Y(n_3796)
);

OAI22xp5_ASAP7_75t_L g3797 ( 
.A1(n_3664),
.A2(n_3129),
.B1(n_3136),
.B2(n_3130),
.Y(n_3797)
);

OAI21xp33_ASAP7_75t_L g3798 ( 
.A1(n_3615),
.A2(n_2971),
.B(n_3311),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3664),
.B(n_3354),
.Y(n_3799)
);

INVxp67_ASAP7_75t_L g3800 ( 
.A(n_3462),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3619),
.A2(n_3295),
.B(n_3144),
.C(n_3150),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3401),
.B(n_3137),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3444),
.B(n_3354),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3395),
.Y(n_3804)
);

OAI22xp5_ASAP7_75t_L g3805 ( 
.A1(n_3540),
.A2(n_3151),
.B1(n_3156),
.B2(n_3153),
.Y(n_3805)
);

OAI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3511),
.A2(n_3159),
.B1(n_3162),
.B2(n_3161),
.Y(n_3806)
);

A2O1A1Ixp33_ASAP7_75t_L g3807 ( 
.A1(n_3502),
.A2(n_2965),
.B(n_3325),
.C(n_3062),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3648),
.A2(n_3083),
.B(n_2882),
.Y(n_3808)
);

OAI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3575),
.A2(n_3166),
.B1(n_3171),
.B2(n_3168),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3393),
.A2(n_3083),
.B(n_2882),
.Y(n_3810)
);

OAI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3403),
.A2(n_3376),
.B(n_3351),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3415),
.B(n_3172),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3528),
.B(n_3173),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3528),
.B(n_3174),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3532),
.B(n_3175),
.Y(n_3815)
);

OAI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3502),
.A2(n_3181),
.B1(n_3177),
.B2(n_3188),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3391),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3621),
.A2(n_3325),
.B(n_3356),
.C(n_3348),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3532),
.B(n_3189),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3393),
.A2(n_3344),
.B(n_3307),
.Y(n_3820)
);

BUFx2_ASAP7_75t_L g3821 ( 
.A(n_3417),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3772),
.B(n_3195),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3516),
.B(n_3197),
.Y(n_3823)
);

BUFx12f_ASAP7_75t_L g3824 ( 
.A(n_3448),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3596),
.B(n_3478),
.Y(n_3825)
);

OAI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_3538),
.A2(n_3199),
.B1(n_3201),
.B2(n_3198),
.Y(n_3826)
);

O2A1O1Ixp33_ASAP7_75t_L g3827 ( 
.A1(n_3641),
.A2(n_3734),
.B(n_3591),
.C(n_3478),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3744),
.A2(n_3347),
.B(n_3218),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3503),
.A2(n_3340),
.B(n_3312),
.Y(n_3829)
);

NOR2xp67_ASAP7_75t_L g3830 ( 
.A(n_3620),
.B(n_3182),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3503),
.A2(n_3340),
.B(n_3352),
.Y(n_3831)
);

AND2x4_ASAP7_75t_L g3832 ( 
.A(n_3533),
.B(n_2989),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3684),
.B(n_3215),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3512),
.A2(n_3365),
.B(n_3364),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3689),
.B(n_3219),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3642),
.B(n_3336),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3405),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3509),
.B(n_3219),
.Y(n_3838)
);

NOR3xp33_ASAP7_75t_SL g3839 ( 
.A(n_3526),
.B(n_3241),
.C(n_3228),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3512),
.A2(n_3381),
.B(n_3375),
.Y(n_3840)
);

O2A1O1Ixp33_ASAP7_75t_SL g3841 ( 
.A1(n_3408),
.A2(n_2934),
.B(n_2924),
.C(n_3202),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3518),
.A2(n_3296),
.B(n_2613),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3584),
.B(n_3204),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_SL g3844 ( 
.A(n_3642),
.B(n_3367),
.Y(n_3844)
);

O2A1O1Ixp33_ASAP7_75t_L g3845 ( 
.A1(n_3419),
.A2(n_3207),
.B(n_3210),
.C(n_3205),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3456),
.B(n_3148),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3588),
.B(n_3359),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3518),
.A2(n_2613),
.B(n_3341),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3498),
.B(n_3214),
.Y(n_3849)
);

BUFx3_ASAP7_75t_L g3850 ( 
.A(n_3399),
.Y(n_3850)
);

OAI321xp33_ASAP7_75t_L g3851 ( 
.A1(n_3495),
.A2(n_867),
.A3(n_861),
.B1(n_870),
.B2(n_864),
.C(n_863),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3521),
.A2(n_2613),
.B(n_2893),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3519),
.B(n_3359),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3405),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3394),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3400),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3521),
.A2(n_2613),
.B(n_2893),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3457),
.A2(n_2893),
.B(n_2872),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3423),
.B(n_3432),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3576),
.B(n_3228),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_SL g3861 ( 
.A(n_3456),
.B(n_3320),
.Y(n_3861)
);

OAI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3656),
.A2(n_3376),
.B(n_2941),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3475),
.B(n_3080),
.Y(n_3863)
);

AND2x4_ASAP7_75t_L g3864 ( 
.A(n_3533),
.B(n_2989),
.Y(n_3864)
);

OAI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3656),
.A2(n_3356),
.B(n_3348),
.Y(n_3865)
);

AOI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3668),
.A2(n_3081),
.B1(n_2981),
.B2(n_3200),
.Y(n_3866)
);

INVxp67_ASAP7_75t_L g3867 ( 
.A(n_3402),
.Y(n_3867)
);

AOI21xp33_ASAP7_75t_L g3868 ( 
.A1(n_3631),
.A2(n_3632),
.B(n_3621),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_L g3869 ( 
.A(n_3475),
.B(n_3203),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3593),
.A2(n_3370),
.B(n_3360),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3416),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3754),
.A2(n_3217),
.B1(n_3221),
.B2(n_3216),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3423),
.B(n_3226),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_L g3874 ( 
.A(n_3683),
.B(n_3081),
.Y(n_3874)
);

AOI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3718),
.A2(n_3187),
.B1(n_3107),
.B2(n_3387),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3397),
.B(n_3330),
.Y(n_3876)
);

OAI321xp33_ASAP7_75t_L g3877 ( 
.A1(n_3649),
.A2(n_879),
.A3(n_864),
.B1(n_882),
.B2(n_870),
.C(n_867),
.Y(n_3877)
);

A2O1A1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_3616),
.A2(n_3481),
.B(n_3654),
.C(n_3650),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3457),
.A2(n_2893),
.B(n_2872),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3426),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3594),
.A2(n_2893),
.B(n_2872),
.Y(n_3881)
);

O2A1O1Ixp33_ASAP7_75t_L g3882 ( 
.A1(n_3489),
.A2(n_3227),
.B(n_3235),
.C(n_3229),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3413),
.B(n_3330),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3544),
.A2(n_3507),
.B(n_3536),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3428),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3544),
.A2(n_2893),
.B(n_2872),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3432),
.B(n_3236),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3474),
.B(n_3330),
.Y(n_3888)
);

A2O1A1Ixp33_ASAP7_75t_L g3889 ( 
.A1(n_3616),
.A2(n_3370),
.B(n_3360),
.C(n_3238),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3434),
.B(n_3436),
.Y(n_3890)
);

AND2x4_ASAP7_75t_L g3891 ( 
.A(n_3651),
.B(n_2989),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3422),
.B(n_3208),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3544),
.A2(n_2872),
.B(n_2789),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_3421),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_3427),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3439),
.B(n_3237),
.Y(n_3896)
);

A2O1A1Ixp33_ASAP7_75t_L g3897 ( 
.A1(n_3650),
.A2(n_3242),
.B(n_3243),
.C(n_3239),
.Y(n_3897)
);

NAND2x1p5_ASAP7_75t_L g3898 ( 
.A(n_3544),
.B(n_3384),
.Y(n_3898)
);

INVx4_ASAP7_75t_L g3899 ( 
.A(n_3496),
.Y(n_3899)
);

AOI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_3536),
.A2(n_2872),
.B(n_2789),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3542),
.A2(n_2878),
.B(n_2789),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3542),
.A2(n_2878),
.B(n_2789),
.Y(n_3902)
);

NOR2xp33_ASAP7_75t_L g3903 ( 
.A(n_3508),
.B(n_3120),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3514),
.A2(n_2878),
.B(n_2789),
.Y(n_3904)
);

OAI21xp33_ASAP7_75t_L g3905 ( 
.A1(n_3494),
.A2(n_761),
.B(n_750),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_3466),
.B(n_3036),
.Y(n_3906)
);

NAND2x1p5_ASAP7_75t_L g3907 ( 
.A(n_3741),
.B(n_3362),
.Y(n_3907)
);

O2A1O1Ixp5_ASAP7_75t_L g3908 ( 
.A1(n_3672),
.A2(n_3167),
.B(n_3249),
.C(n_3245),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3626),
.A2(n_3377),
.B(n_3372),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3515),
.A2(n_2878),
.B(n_2789),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_3551),
.B(n_3047),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3633),
.A2(n_2878),
.B(n_3000),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3446),
.A2(n_2878),
.B(n_3000),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3392),
.B(n_3254),
.Y(n_3914)
);

OR2x2_ASAP7_75t_L g3915 ( 
.A(n_3556),
.B(n_3761),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3461),
.A2(n_3002),
.B(n_3100),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3628),
.A2(n_3380),
.B(n_3379),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3510),
.A2(n_3002),
.B(n_3100),
.Y(n_3918)
);

AOI21x1_ASAP7_75t_L g3919 ( 
.A1(n_3659),
.A2(n_3680),
.B(n_3637),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3587),
.A2(n_3601),
.B(n_3614),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3715),
.B(n_3337),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_3560),
.B(n_3047),
.Y(n_3922)
);

NAND2x1p5_ASAP7_75t_L g3923 ( 
.A(n_3741),
.B(n_3389),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3718),
.B(n_3302),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3654),
.A2(n_3644),
.B(n_3705),
.C(n_3699),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3476),
.A2(n_2659),
.B(n_2488),
.Y(n_3926)
);

NOR2xp33_ASAP7_75t_L g3927 ( 
.A(n_3724),
.B(n_3357),
.Y(n_3927)
);

AOI22xp5_ASAP7_75t_L g3928 ( 
.A1(n_3724),
.A2(n_3241),
.B1(n_3132),
.B2(n_3366),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3497),
.B(n_3337),
.Y(n_3929)
);

O2A1O1Ixp33_ASAP7_75t_L g3930 ( 
.A1(n_3572),
.A2(n_3259),
.B(n_3265),
.C(n_3264),
.Y(n_3930)
);

HB1xp67_ASAP7_75t_L g3931 ( 
.A(n_3398),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3459),
.B(n_3273),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3570),
.B(n_3630),
.Y(n_3933)
);

BUFx4f_ASAP7_75t_L g3934 ( 
.A(n_3496),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3720),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3630),
.B(n_3277),
.Y(n_3936)
);

AOI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3517),
.A2(n_3132),
.B1(n_3368),
.B2(n_3366),
.Y(n_3937)
);

A2O1A1Ixp33_ASAP7_75t_L g3938 ( 
.A1(n_3699),
.A2(n_3281),
.B(n_3282),
.C(n_3279),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3543),
.A2(n_2673),
.B(n_2659),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3543),
.A2(n_2673),
.B(n_2659),
.Y(n_3940)
);

AOI21xp5_ASAP7_75t_L g3941 ( 
.A1(n_3553),
.A2(n_3558),
.B(n_3557),
.Y(n_3941)
);

AOI21x1_ASAP7_75t_L g3942 ( 
.A1(n_3563),
.A2(n_2887),
.B(n_2770),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3441),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3418),
.B(n_3486),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3442),
.Y(n_3945)
);

BUFx3_ASAP7_75t_L g3946 ( 
.A(n_3421),
.Y(n_3946)
);

NAND2x1p5_ASAP7_75t_L g3947 ( 
.A(n_3663),
.B(n_3386),
.Y(n_3947)
);

NOR2x1_ASAP7_75t_R g3948 ( 
.A(n_3657),
.B(n_1780),
.Y(n_3948)
);

NAND2x1p5_ASAP7_75t_L g3949 ( 
.A(n_3663),
.B(n_3385),
.Y(n_3949)
);

NOR2xp67_ASAP7_75t_L g3950 ( 
.A(n_3752),
.B(n_3261),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3553),
.A2(n_2678),
.B(n_2673),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_3706),
.B(n_3132),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3420),
.B(n_3288),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3722),
.B(n_3046),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3443),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3406),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3754),
.A2(n_3291),
.B1(n_3292),
.B2(n_3289),
.Y(n_3957)
);

AOI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3735),
.A2(n_3366),
.B1(n_3368),
.B2(n_3337),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3557),
.A2(n_2780),
.B(n_2678),
.Y(n_3959)
);

OAI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3600),
.A2(n_3308),
.B1(n_3310),
.B2(n_3297),
.Y(n_3960)
);

O2A1O1Ixp33_ASAP7_75t_L g3961 ( 
.A1(n_3696),
.A2(n_3313),
.B(n_3317),
.C(n_3316),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3406),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3486),
.B(n_3323),
.Y(n_3963)
);

OAI21x1_ASAP7_75t_L g3964 ( 
.A1(n_3470),
.A2(n_2887),
.B(n_3371),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3739),
.B(n_1813),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3558),
.A2(n_2780),
.B(n_2678),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3452),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3646),
.B(n_3047),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3727),
.A2(n_2819),
.B(n_2780),
.Y(n_3969)
);

BUFx4f_ASAP7_75t_L g3970 ( 
.A(n_3496),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3431),
.A2(n_2843),
.B(n_2819),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3453),
.Y(n_3972)
);

HB1xp67_ASAP7_75t_L g3973 ( 
.A(n_3398),
.Y(n_3973)
);

A2O1A1Ixp33_ASAP7_75t_L g3974 ( 
.A1(n_3705),
.A2(n_3328),
.B(n_3332),
.C(n_3324),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3425),
.B(n_3334),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3465),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3431),
.A2(n_2843),
.B(n_2819),
.Y(n_3977)
);

O2A1O1Ixp33_ASAP7_75t_L g3978 ( 
.A1(n_3541),
.A2(n_2042),
.B(n_1809),
.C(n_1821),
.Y(n_3978)
);

AOI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3445),
.A2(n_3450),
.B(n_3574),
.Y(n_3979)
);

HB1xp67_ASAP7_75t_L g3980 ( 
.A(n_3454),
.Y(n_3980)
);

AOI21xp5_ASAP7_75t_L g3981 ( 
.A1(n_3445),
.A2(n_2843),
.B(n_3051),
.Y(n_3981)
);

INVx3_ASAP7_75t_L g3982 ( 
.A(n_3651),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3450),
.A2(n_2991),
.B(n_2959),
.Y(n_3983)
);

INVxp67_ASAP7_75t_SL g3984 ( 
.A(n_3607),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_L g3985 ( 
.A(n_3745),
.B(n_1822),
.Y(n_3985)
);

AOI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3574),
.A2(n_2991),
.B(n_2959),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3774),
.B(n_1831),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3479),
.B(n_3222),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3480),
.B(n_3222),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3463),
.B(n_3247),
.Y(n_3990)
);

AND2x4_ASAP7_75t_L g3991 ( 
.A(n_3685),
.B(n_3629),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3412),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3472),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3585),
.A2(n_2706),
.B(n_2670),
.Y(n_3994)
);

AO21x1_ASAP7_75t_L g3995 ( 
.A1(n_3678),
.A2(n_3329),
.B(n_3338),
.Y(n_3995)
);

OAI21x1_ASAP7_75t_L g3996 ( 
.A1(n_3468),
.A2(n_3388),
.B(n_3371),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_L g3997 ( 
.A(n_3589),
.B(n_1831),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3589),
.B(n_1839),
.Y(n_3998)
);

BUFx3_ASAP7_75t_L g3999 ( 
.A(n_3454),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3412),
.Y(n_4000)
);

AOI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3735),
.A2(n_3368),
.B1(n_3009),
.B2(n_3017),
.Y(n_4001)
);

AOI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3585),
.A2(n_2871),
.B(n_2670),
.Y(n_4002)
);

O2A1O1Ixp33_ASAP7_75t_L g4003 ( 
.A1(n_3529),
.A2(n_3494),
.B(n_3738),
.C(n_3564),
.Y(n_4003)
);

O2A1O1Ixp33_ASAP7_75t_L g4004 ( 
.A1(n_3737),
.A2(n_1827),
.B(n_1859),
.C(n_1806),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3547),
.B(n_3247),
.Y(n_4005)
);

AOI21x1_ASAP7_75t_L g4006 ( 
.A1(n_3592),
.A2(n_3343),
.B(n_3342),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3501),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3513),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3592),
.A2(n_2706),
.B(n_2670),
.Y(n_4009)
);

INVx3_ASAP7_75t_L g4010 ( 
.A(n_3685),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3595),
.A2(n_3647),
.B(n_3623),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3471),
.B(n_3520),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3527),
.B(n_3253),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3530),
.B(n_3253),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3427),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3595),
.A2(n_2706),
.B(n_2670),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3549),
.B(n_3255),
.Y(n_4017)
);

OAI21xp33_ASAP7_75t_L g4018 ( 
.A1(n_3429),
.A2(n_850),
.B(n_803),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3524),
.B(n_3142),
.Y(n_4019)
);

AOI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3623),
.A2(n_3653),
.B(n_3647),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3653),
.A2(n_2791),
.B(n_2706),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3546),
.Y(n_4022)
);

INVx3_ASAP7_75t_L g4023 ( 
.A(n_3458),
.Y(n_4023)
);

NOR2xp33_ASAP7_75t_L g4024 ( 
.A(n_3773),
.B(n_1944),
.Y(n_4024)
);

BUFx6f_ASAP7_75t_L g4025 ( 
.A(n_3427),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3666),
.A2(n_2871),
.B(n_2825),
.Y(n_4026)
);

NOR2xp33_ASAP7_75t_L g4027 ( 
.A(n_3464),
.B(n_2013),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3550),
.Y(n_4028)
);

BUFx6f_ASAP7_75t_L g4029 ( 
.A(n_3427),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3555),
.B(n_3255),
.Y(n_4030)
);

AOI21xp5_ASAP7_75t_L g4031 ( 
.A1(n_3666),
.A2(n_2871),
.B(n_2825),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_3667),
.A2(n_2871),
.B(n_2825),
.Y(n_4032)
);

NOR2x1_ASAP7_75t_L g4033 ( 
.A(n_3580),
.B(n_3017),
.Y(n_4033)
);

NOR2xp33_ASAP7_75t_L g4034 ( 
.A(n_3665),
.B(n_2013),
.Y(n_4034)
);

INVxp67_ASAP7_75t_L g4035 ( 
.A(n_3697),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3531),
.B(n_3256),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3578),
.B(n_3256),
.Y(n_4037)
);

OAI321xp33_ASAP7_75t_L g4038 ( 
.A1(n_3433),
.A2(n_882),
.A3(n_884),
.B1(n_891),
.B2(n_888),
.C(n_879),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3582),
.B(n_3263),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3414),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3679),
.B(n_3142),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_3635),
.B(n_3142),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3414),
.Y(n_4043)
);

A2O1A1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3602),
.A2(n_3145),
.B(n_3163),
.C(n_3147),
.Y(n_4044)
);

BUFx2_ASAP7_75t_L g4045 ( 
.A(n_3447),
.Y(n_4045)
);

OAI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_3600),
.A2(n_3695),
.B1(n_3782),
.B2(n_3410),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3586),
.B(n_3602),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3565),
.B(n_3263),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3430),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_3786),
.Y(n_4050)
);

OAI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3611),
.A2(n_3147),
.B(n_3145),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3566),
.B(n_3145),
.Y(n_4052)
);

NAND2xp33_ASAP7_75t_L g4053 ( 
.A(n_3755),
.B(n_3369),
.Y(n_4053)
);

O2A1O1Ixp33_ASAP7_75t_L g4054 ( 
.A1(n_3559),
.A2(n_1871),
.B(n_1878),
.C(n_1868),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3667),
.A2(n_3483),
.B(n_3468),
.Y(n_4055)
);

O2A1O1Ixp33_ASAP7_75t_L g4056 ( 
.A1(n_3561),
.A2(n_1887),
.B(n_1888),
.C(n_1880),
.Y(n_4056)
);

A2O1A1Ixp33_ASAP7_75t_L g4057 ( 
.A1(n_3627),
.A2(n_3147),
.B(n_3163),
.C(n_3345),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3483),
.A2(n_2825),
.B(n_2791),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3435),
.A2(n_3163),
.B1(n_2761),
.B2(n_3014),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3568),
.B(n_3388),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3492),
.A2(n_2791),
.B(n_2810),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3569),
.B(n_3573),
.Y(n_4062)
);

INVx11_ASAP7_75t_L g4063 ( 
.A(n_3448),
.Y(n_4063)
);

BUFx8_ASAP7_75t_L g4064 ( 
.A(n_3562),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3579),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3590),
.B(n_3358),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3430),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_3567),
.B(n_2989),
.Y(n_4068)
);

OAI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3449),
.A2(n_3643),
.B(n_3640),
.Y(n_4069)
);

OAI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3460),
.A2(n_3353),
.B(n_3350),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3635),
.B(n_2013),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3598),
.B(n_3605),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_3438),
.Y(n_4073)
);

AOI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3554),
.A2(n_3131),
.B1(n_3014),
.B2(n_2052),
.Y(n_4074)
);

AOI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_3492),
.A2(n_2791),
.B(n_3149),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3606),
.B(n_3267),
.Y(n_4076)
);

INVx3_ASAP7_75t_L g4077 ( 
.A(n_3458),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3622),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3645),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_3655),
.B(n_3267),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3658),
.B(n_3284),
.Y(n_4081)
);

OR2x2_ASAP7_75t_L g4082 ( 
.A(n_3660),
.B(n_3014),
.Y(n_4082)
);

HB1xp67_ASAP7_75t_L g4083 ( 
.A(n_3669),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3686),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3437),
.A2(n_2761),
.B1(n_3131),
.B2(n_3014),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3567),
.B(n_3131),
.Y(n_4086)
);

INVx4_ASAP7_75t_L g4087 ( 
.A(n_3467),
.Y(n_4087)
);

AOI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_3678),
.A2(n_3186),
.B(n_3180),
.Y(n_4088)
);

OAI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_3612),
.A2(n_3355),
.B(n_3315),
.Y(n_4089)
);

BUFx6f_ASAP7_75t_L g4090 ( 
.A(n_3467),
.Y(n_4090)
);

NAND3xp33_ASAP7_75t_L g4091 ( 
.A(n_3548),
.B(n_2052),
.C(n_858),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_3635),
.B(n_2052),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3688),
.A2(n_3186),
.B(n_3180),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3778),
.B(n_3779),
.Y(n_4094)
);

BUFx2_ASAP7_75t_L g4095 ( 
.A(n_3712),
.Y(n_4095)
);

INVx1_ASAP7_75t_SL g4096 ( 
.A(n_3712),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3390),
.B(n_3131),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3692),
.B(n_3327),
.Y(n_4098)
);

INVx2_ASAP7_75t_SL g4099 ( 
.A(n_3581),
.Y(n_4099)
);

AOI22xp33_ASAP7_75t_L g4100 ( 
.A1(n_3567),
.A2(n_2761),
.B1(n_3211),
.B2(n_3190),
.Y(n_4100)
);

OAI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_3618),
.A2(n_3331),
.B(n_3327),
.Y(n_4101)
);

NAND2x1p5_ASAP7_75t_L g4102 ( 
.A(n_3663),
.B(n_3190),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3778),
.B(n_3211),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3702),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3779),
.B(n_3225),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3704),
.B(n_3358),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3688),
.A2(n_3240),
.B(n_3225),
.Y(n_4107)
);

CKINVDCx8_ASAP7_75t_R g4108 ( 
.A(n_3652),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3732),
.B(n_3240),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3390),
.B(n_3246),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_3743),
.Y(n_4111)
);

A2O1A1Ixp33_ASAP7_75t_L g4112 ( 
.A1(n_3757),
.A2(n_3284),
.B(n_3285),
.C(n_3246),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_3757),
.A2(n_3315),
.B(n_3318),
.C(n_3285),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3438),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3746),
.B(n_3318),
.Y(n_4115)
);

OAI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_3695),
.A2(n_3759),
.B1(n_3763),
.B2(n_3758),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_3467),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3764),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3776),
.Y(n_4119)
);

OAI21xp33_ASAP7_75t_L g4120 ( 
.A1(n_3552),
.A2(n_1028),
.B(n_894),
.Y(n_4120)
);

AOI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_3693),
.A2(n_3710),
.B(n_3709),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_3783),
.A2(n_3349),
.B1(n_3326),
.B2(n_3331),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_3396),
.B(n_3319),
.Y(n_4123)
);

OR2x6_ASAP7_75t_L g4124 ( 
.A(n_3458),
.B(n_3319),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3783),
.B(n_3326),
.Y(n_4125)
);

CKINVDCx8_ASAP7_75t_R g4126 ( 
.A(n_3467),
.Y(n_4126)
);

BUFx6f_ASAP7_75t_L g4127 ( 
.A(n_3663),
.Y(n_4127)
);

INVx4_ASAP7_75t_L g4128 ( 
.A(n_3682),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_3693),
.A2(n_3349),
.B(n_2950),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3440),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3604),
.B(n_2761),
.Y(n_4131)
);

AO21x1_ASAP7_75t_L g4132 ( 
.A1(n_3709),
.A2(n_2409),
.B(n_2406),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3607),
.B(n_2483),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3608),
.B(n_2483),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_3571),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3613),
.B(n_2486),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_L g4137 ( 
.A(n_3396),
.B(n_2486),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3755),
.B(n_2495),
.Y(n_4138)
);

NOR2x1_ASAP7_75t_L g4139 ( 
.A(n_3424),
.B(n_2495),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_3571),
.B(n_824),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_3710),
.A2(n_2498),
.B(n_2495),
.Y(n_4141)
);

AO21x1_ASAP7_75t_L g4142 ( 
.A1(n_3711),
.A2(n_2409),
.B(n_2454),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3487),
.B(n_2761),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3490),
.B(n_2761),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_L g4145 ( 
.A(n_3554),
.B(n_2498),
.Y(n_4145)
);

CKINVDCx8_ASAP7_75t_R g4146 ( 
.A(n_3661),
.Y(n_4146)
);

OR2x2_ASAP7_75t_L g4147 ( 
.A(n_3491),
.B(n_3493),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_SL g4148 ( 
.A(n_3661),
.B(n_2885),
.Y(n_4148)
);

INVx3_ASAP7_75t_SL g4149 ( 
.A(n_3581),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3711),
.A2(n_2498),
.B(n_2620),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3499),
.B(n_3369),
.Y(n_4151)
);

NOR2x1p5_ASAP7_75t_L g4152 ( 
.A(n_3624),
.B(n_1506),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3440),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3505),
.B(n_3369),
.Y(n_4154)
);

BUFx6f_ASAP7_75t_L g4155 ( 
.A(n_3682),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_SL g4156 ( 
.A(n_3661),
.B(n_2885),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3571),
.B(n_2582),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3760),
.B(n_2582),
.Y(n_4158)
);

NAND2x1_ASAP7_75t_L g4159 ( 
.A(n_3682),
.B(n_2582),
.Y(n_4159)
);

O2A1O1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_3781),
.A2(n_1028),
.B(n_1091),
.C(n_894),
.Y(n_4160)
);

INVx3_ASAP7_75t_L g4161 ( 
.A(n_3691),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3750),
.A2(n_2620),
.B(n_2587),
.Y(n_4162)
);

AOI21xp33_ASAP7_75t_L g4163 ( 
.A1(n_3500),
.A2(n_2587),
.B(n_2584),
.Y(n_4163)
);

OAI321xp33_ASAP7_75t_L g4164 ( 
.A1(n_3748),
.A2(n_888),
.A3(n_891),
.B1(n_896),
.B2(n_895),
.C(n_884),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4062),
.Y(n_4165)
);

NAND2x1p5_ASAP7_75t_L g4166 ( 
.A(n_4023),
.B(n_3682),
.Y(n_4166)
);

AOI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_3791),
.A2(n_3610),
.B(n_3750),
.Y(n_4167)
);

OAI21xp33_ASAP7_75t_L g4168 ( 
.A1(n_3905),
.A2(n_3775),
.B(n_3617),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_3899),
.B(n_3624),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3793),
.B(n_3760),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_3847),
.A2(n_3634),
.B1(n_3577),
.B2(n_3662),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3790),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_SL g4173 ( 
.A(n_3859),
.B(n_3762),
.Y(n_4173)
);

AND2x4_ASAP7_75t_L g4174 ( 
.A(n_3899),
.B(n_3662),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_SL g4175 ( 
.A(n_3827),
.B(n_3762),
.Y(n_4175)
);

BUFx3_ASAP7_75t_L g4176 ( 
.A(n_3796),
.Y(n_4176)
);

AOI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_4053),
.A2(n_3691),
.B(n_3781),
.Y(n_4177)
);

INVxp67_ASAP7_75t_SL g4178 ( 
.A(n_4137),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_3820),
.A2(n_3691),
.B(n_3784),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_SL g4180 ( 
.A(n_3825),
.B(n_3725),
.Y(n_4180)
);

AOI21xp5_ASAP7_75t_L g4181 ( 
.A1(n_3834),
.A2(n_3784),
.B(n_3787),
.Y(n_4181)
);

BUFx2_ASAP7_75t_L g4182 ( 
.A(n_3821),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3792),
.B(n_3451),
.Y(n_4183)
);

AOI22xp33_ASAP7_75t_SL g4184 ( 
.A1(n_3924),
.A2(n_3525),
.B1(n_3755),
.B2(n_1097),
.Y(n_4184)
);

AO22x1_ASAP7_75t_L g4185 ( 
.A1(n_4027),
.A2(n_3525),
.B1(n_1194),
.B2(n_1097),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_3850),
.Y(n_4186)
);

BUFx8_ASAP7_75t_L g4187 ( 
.A(n_3824),
.Y(n_4187)
);

AOI33xp33_ASAP7_75t_L g4188 ( 
.A1(n_4160),
.A2(n_1248),
.A3(n_1112),
.B1(n_1154),
.B2(n_1091),
.B3(n_896),
.Y(n_4188)
);

INVxp67_ASAP7_75t_L g4189 ( 
.A(n_3853),
.Y(n_4189)
);

HB1xp67_ASAP7_75t_L g4190 ( 
.A(n_3800),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3933),
.B(n_3451),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_3867),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3838),
.B(n_3455),
.Y(n_4193)
);

AOI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3788),
.A2(n_3537),
.B1(n_3535),
.B2(n_3755),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3804),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_3835),
.B(n_3455),
.Y(n_4196)
);

OA22x2_ASAP7_75t_L g4197 ( 
.A1(n_4001),
.A2(n_1154),
.B1(n_1248),
.B2(n_1112),
.Y(n_4197)
);

NOR3xp33_ASAP7_75t_L g4198 ( 
.A(n_3877),
.B(n_1512),
.C(n_1508),
.Y(n_4198)
);

AOI21x1_ASAP7_75t_L g4199 ( 
.A1(n_3942),
.A2(n_3794),
.B(n_3919),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_3860),
.B(n_1582),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3863),
.B(n_3681),
.Y(n_4201)
);

OA22x2_ASAP7_75t_L g4202 ( 
.A1(n_3799),
.A2(n_3928),
.B1(n_3798),
.B2(n_3836),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3840),
.A2(n_3733),
.B(n_3780),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3944),
.B(n_3469),
.Y(n_4204)
);

NAND2x1p5_ASAP7_75t_L g4205 ( 
.A(n_4023),
.B(n_3733),
.Y(n_4205)
);

NOR2xp33_ASAP7_75t_L g4206 ( 
.A(n_3803),
.B(n_3687),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3914),
.B(n_3469),
.Y(n_4207)
);

NOR2x1_ASAP7_75t_L g4208 ( 
.A(n_3822),
.B(n_3411),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3823),
.B(n_3473),
.Y(n_4209)
);

NOR2xp33_ASAP7_75t_L g4210 ( 
.A(n_3861),
.B(n_3690),
.Y(n_4210)
);

OAI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4094),
.A2(n_3751),
.B1(n_3670),
.B2(n_3721),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4072),
.Y(n_4212)
);

OA22x2_ASAP7_75t_L g4213 ( 
.A1(n_3846),
.A2(n_3875),
.B1(n_3844),
.B2(n_4035),
.Y(n_4213)
);

INVxp33_ASAP7_75t_SL g4214 ( 
.A(n_4050),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_3828),
.A2(n_3733),
.B(n_3785),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3837),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3854),
.Y(n_4217)
);

A2O1A1Ixp33_ASAP7_75t_SL g4218 ( 
.A1(n_3998),
.A2(n_3599),
.B(n_3771),
.C(n_3769),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3823),
.B(n_3915),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_3869),
.B(n_3700),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3849),
.B(n_3473),
.Y(n_4221)
);

BUFx6f_ASAP7_75t_SL g4222 ( 
.A(n_3894),
.Y(n_4222)
);

AOI21x1_ASAP7_75t_L g4223 ( 
.A1(n_3808),
.A2(n_3717),
.B(n_3707),
.Y(n_4223)
);

NOR2xp67_ASAP7_75t_L g4224 ( 
.A(n_3952),
.B(n_3411),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_3843),
.B(n_3482),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3817),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3802),
.B(n_3482),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_3956),
.Y(n_4228)
);

OAI22xp5_ASAP7_75t_L g4229 ( 
.A1(n_4094),
.A2(n_3698),
.B1(n_3765),
.B2(n_3749),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_R g4230 ( 
.A(n_4146),
.B(n_3733),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3802),
.B(n_3485),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3932),
.B(n_3485),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_3829),
.A2(n_3768),
.B(n_3766),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_SL g4234 ( 
.A(n_3948),
.B(n_4108),
.Y(n_4234)
);

INVxp67_ASAP7_75t_L g4235 ( 
.A(n_3980),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_3813),
.A2(n_3814),
.B1(n_3819),
.B2(n_3815),
.Y(n_4236)
);

BUFx8_ASAP7_75t_L g4237 ( 
.A(n_4045),
.Y(n_4237)
);

HB1xp67_ASAP7_75t_L g4238 ( 
.A(n_3935),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3873),
.B(n_3488),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_3921),
.B(n_1583),
.Y(n_4240)
);

NOR2xp33_ASAP7_75t_SL g4241 ( 
.A(n_3934),
.B(n_3755),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3831),
.A2(n_3777),
.B(n_3770),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3870),
.A2(n_3708),
.B(n_3701),
.Y(n_4243)
);

INVx3_ASAP7_75t_L g4244 ( 
.A(n_4124),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_3927),
.B(n_3795),
.Y(n_4245)
);

OAI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_3813),
.A2(n_3719),
.B1(n_3723),
.B2(n_3716),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3887),
.B(n_3488),
.Y(n_4247)
);

NOR2xp67_ASAP7_75t_SL g4248 ( 
.A(n_3851),
.B(n_3477),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_3814),
.A2(n_3731),
.B1(n_3730),
.B2(n_3729),
.Y(n_4249)
);

AND2x4_ASAP7_75t_L g4250 ( 
.A(n_3991),
.B(n_3477),
.Y(n_4250)
);

AOI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3789),
.A2(n_3522),
.B(n_3504),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3997),
.B(n_3756),
.Y(n_4252)
);

NOR2xp33_ASAP7_75t_L g4253 ( 
.A(n_3874),
.B(n_856),
.Y(n_4253)
);

AOI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_3881),
.A2(n_3522),
.B(n_3504),
.Y(n_4254)
);

O2A1O1Ixp33_ASAP7_75t_L g4255 ( 
.A1(n_3807),
.A2(n_905),
.B(n_906),
.C(n_895),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_3962),
.Y(n_4256)
);

OR2x2_ASAP7_75t_L g4257 ( 
.A(n_4096),
.B(n_3523),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_SL g4258 ( 
.A(n_3815),
.B(n_3756),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_3865),
.A2(n_3534),
.B(n_3523),
.Y(n_4259)
);

O2A1O1Ixp33_ASAP7_75t_L g4260 ( 
.A1(n_4164),
.A2(n_906),
.B(n_914),
.C(n_905),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_3819),
.B(n_3534),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_SL g4262 ( 
.A1(n_3866),
.A2(n_4024),
.B1(n_3903),
.B2(n_4034),
.Y(n_4262)
);

CKINVDCx16_ASAP7_75t_R g4263 ( 
.A(n_3946),
.Y(n_4263)
);

AOI21xp5_ASAP7_75t_L g4264 ( 
.A1(n_3818),
.A2(n_3583),
.B(n_3545),
.Y(n_4264)
);

O2A1O1Ixp33_ASAP7_75t_L g4265 ( 
.A1(n_3801),
.A2(n_918),
.B(n_923),
.C(n_914),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_3812),
.B(n_3545),
.Y(n_4266)
);

INVx5_ASAP7_75t_L g4267 ( 
.A(n_4124),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3958),
.B(n_3756),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3812),
.B(n_3583),
.Y(n_4269)
);

OAI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4046),
.A2(n_3713),
.B1(n_3714),
.B2(n_3703),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3992),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_4046),
.A2(n_3833),
.B1(n_3822),
.B2(n_4047),
.Y(n_4272)
);

AOI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_3950),
.A2(n_862),
.B1(n_865),
.B2(n_859),
.Y(n_4273)
);

OAI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_3896),
.A2(n_3728),
.B1(n_3729),
.B2(n_3726),
.Y(n_4274)
);

NOR2x1_ASAP7_75t_L g4275 ( 
.A(n_3968),
.B(n_3597),
.Y(n_4275)
);

HB1xp67_ASAP7_75t_L g4276 ( 
.A(n_4135),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_3963),
.B(n_4018),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_3876),
.B(n_1585),
.Y(n_4278)
);

A2O1A1Ixp33_ASAP7_75t_L g4279 ( 
.A1(n_4003),
.A2(n_3603),
.B(n_3625),
.C(n_3597),
.Y(n_4279)
);

INVx3_ASAP7_75t_L g4280 ( 
.A(n_4124),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_3855),
.Y(n_4281)
);

CKINVDCx5p33_ASAP7_75t_R g4282 ( 
.A(n_4063),
.Y(n_4282)
);

OAI22xp5_ASAP7_75t_L g4283 ( 
.A1(n_3890),
.A2(n_3740),
.B1(n_3747),
.B2(n_3736),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3856),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3888),
.B(n_3603),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_3883),
.B(n_866),
.Y(n_4286)
);

AO21x1_ASAP7_75t_L g4287 ( 
.A1(n_3960),
.A2(n_3636),
.B(n_3625),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3936),
.B(n_3636),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_4126),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_SL g4290 ( 
.A(n_3839),
.B(n_3756),
.Y(n_4290)
);

NOR2xp33_ASAP7_75t_L g4291 ( 
.A(n_4095),
.B(n_869),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_3920),
.A2(n_3639),
.B(n_3638),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4012),
.B(n_3638),
.Y(n_4293)
);

AOI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_3886),
.A2(n_3671),
.B(n_3639),
.Y(n_4294)
);

OAI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_3925),
.A2(n_3675),
.B(n_3671),
.Y(n_4295)
);

OR2x6_ASAP7_75t_L g4296 ( 
.A(n_3941),
.B(n_3675),
.Y(n_4296)
);

A2O1A1Ixp33_ASAP7_75t_SL g4297 ( 
.A1(n_3965),
.A2(n_3677),
.B(n_3703),
.C(n_3694),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3871),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4012),
.B(n_3676),
.Y(n_4299)
);

AO22x1_ASAP7_75t_L g4300 ( 
.A1(n_4033),
.A2(n_872),
.B1(n_874),
.B2(n_871),
.Y(n_4300)
);

CKINVDCx16_ASAP7_75t_R g4301 ( 
.A(n_3999),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4120),
.B(n_3676),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4147),
.B(n_3677),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4000),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_3848),
.A2(n_3713),
.B(n_3694),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_3929),
.B(n_3714),
.Y(n_4306)
);

AOI21xp33_ASAP7_75t_L g4307 ( 
.A1(n_3845),
.A2(n_3728),
.B(n_3726),
.Y(n_4307)
);

INVx3_ASAP7_75t_L g4308 ( 
.A(n_3934),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_L g4309 ( 
.A(n_3954),
.B(n_3892),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_3953),
.B(n_3975),
.Y(n_4310)
);

AND2x4_ASAP7_75t_L g4311 ( 
.A(n_3991),
.B(n_3736),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_3953),
.B(n_3740),
.Y(n_4312)
);

NOR2xp33_ASAP7_75t_L g4313 ( 
.A(n_3906),
.B(n_876),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4040),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4083),
.B(n_4111),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_3884),
.A2(n_3753),
.B(n_3747),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4091),
.B(n_3756),
.Y(n_4317)
);

O2A1O1Ixp33_ASAP7_75t_L g4318 ( 
.A1(n_3878),
.A2(n_3868),
.B(n_3889),
.C(n_4071),
.Y(n_4318)
);

OAI22xp5_ASAP7_75t_L g4319 ( 
.A1(n_3937),
.A2(n_3767),
.B1(n_3769),
.B2(n_3753),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4140),
.B(n_3767),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4052),
.B(n_3771),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_3983),
.A2(n_3756),
.B(n_2587),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_3880),
.B(n_1586),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_3868),
.B(n_877),
.Y(n_4324)
);

NOR2xp33_ASAP7_75t_L g4325 ( 
.A(n_3911),
.B(n_3922),
.Y(n_4325)
);

AOI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_3994),
.A2(n_2588),
.B(n_2584),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4002),
.A2(n_2588),
.B(n_2584),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3806),
.B(n_878),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_4009),
.A2(n_2597),
.B(n_2588),
.Y(n_4329)
);

NOR2xp33_ASAP7_75t_L g4330 ( 
.A(n_3985),
.B(n_880),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_3806),
.B(n_881),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_4044),
.A2(n_886),
.B1(n_890),
.B2(n_885),
.Y(n_4332)
);

OR2x6_ASAP7_75t_L g4333 ( 
.A(n_4077),
.B(n_2597),
.Y(n_4333)
);

AND2x4_ASAP7_75t_L g4334 ( 
.A(n_4068),
.B(n_2603),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4043),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_SL g4336 ( 
.A(n_3811),
.B(n_2885),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3885),
.B(n_892),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_3943),
.B(n_899),
.Y(n_4338)
);

INVx6_ASAP7_75t_L g4339 ( 
.A(n_4064),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3945),
.B(n_901),
.Y(n_4340)
);

AO21x1_ASAP7_75t_L g4341 ( 
.A1(n_3960),
.A2(n_923),
.B(n_918),
.Y(n_4341)
);

NOR2xp67_ASAP7_75t_SL g4342 ( 
.A(n_4038),
.B(n_926),
.Y(n_4342)
);

INVx5_ASAP7_75t_L g4343 ( 
.A(n_3895),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_3955),
.B(n_902),
.Y(n_4344)
);

A2O1A1Ixp33_ASAP7_75t_L g4345 ( 
.A1(n_3882),
.A2(n_929),
.B(n_930),
.C(n_926),
.Y(n_4345)
);

NAND3xp33_ASAP7_75t_SL g4346 ( 
.A(n_4074),
.B(n_908),
.C(n_904),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_3987),
.B(n_907),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3967),
.B(n_915),
.Y(n_4348)
);

BUFx4f_ASAP7_75t_L g4349 ( 
.A(n_4149),
.Y(n_4349)
);

O2A1O1Ixp33_ASAP7_75t_L g4350 ( 
.A1(n_4092),
.A2(n_930),
.B(n_932),
.C(n_929),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4019),
.B(n_1587),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_4059),
.A2(n_922),
.B1(n_927),
.B2(n_921),
.Y(n_4352)
);

BUFx3_ASAP7_75t_L g4353 ( 
.A(n_4064),
.Y(n_4353)
);

AOI21xp5_ASAP7_75t_L g4354 ( 
.A1(n_4016),
.A2(n_2603),
.B(n_2597),
.Y(n_4354)
);

OAI21xp33_ASAP7_75t_L g4355 ( 
.A1(n_4139),
.A2(n_935),
.B(n_934),
.Y(n_4355)
);

AOI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4021),
.A2(n_2607),
.B(n_2603),
.Y(n_4356)
);

NOR2xp33_ASAP7_75t_L g4357 ( 
.A(n_4082),
.B(n_937),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3862),
.A2(n_2610),
.B(n_2607),
.Y(n_4358)
);

BUFx3_ASAP7_75t_L g4359 ( 
.A(n_4099),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_3972),
.B(n_3993),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4049),
.Y(n_4361)
);

OAI21xp33_ASAP7_75t_SL g4362 ( 
.A1(n_4060),
.A2(n_938),
.B(n_932),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_3976),
.Y(n_4363)
);

AOI22xp33_ASAP7_75t_L g4364 ( 
.A1(n_3830),
.A2(n_837),
.B1(n_920),
.B2(n_824),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4007),
.B(n_939),
.Y(n_4365)
);

AOI22xp5_ASAP7_75t_L g4366 ( 
.A1(n_4152),
.A2(n_942),
.B1(n_944),
.B2(n_941),
.Y(n_4366)
);

O2A1O1Ixp33_ASAP7_75t_L g4367 ( 
.A1(n_3897),
.A2(n_943),
.B(n_949),
.C(n_938),
.Y(n_4367)
);

OR2x6_ASAP7_75t_L g4368 ( 
.A(n_4077),
.B(n_2607),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_4008),
.B(n_945),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4022),
.B(n_947),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_4086),
.B(n_4028),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_3797),
.B(n_2885),
.Y(n_4372)
);

NOR2xp33_ASAP7_75t_L g4373 ( 
.A(n_4042),
.B(n_948),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4065),
.B(n_953),
.Y(n_4374)
);

OAI22xp5_ASAP7_75t_L g4375 ( 
.A1(n_3970),
.A2(n_960),
.B1(n_965),
.B2(n_954),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4078),
.B(n_967),
.Y(n_4376)
);

A2O1A1Ixp33_ASAP7_75t_L g4377 ( 
.A1(n_3930),
.A2(n_949),
.B(n_952),
.C(n_943),
.Y(n_4377)
);

AOI22xp5_ASAP7_75t_L g4378 ( 
.A1(n_4041),
.A2(n_978),
.B1(n_980),
.B2(n_971),
.Y(n_4378)
);

AOI21xp5_ASAP7_75t_L g4379 ( 
.A1(n_4026),
.A2(n_2617),
.B(n_2610),
.Y(n_4379)
);

OAI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_3908),
.A2(n_2617),
.B(n_2610),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4067),
.Y(n_4381)
);

OR2x2_ASAP7_75t_L g4382 ( 
.A(n_4079),
.B(n_1625),
.Y(n_4382)
);

OAI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_3926),
.A2(n_2642),
.B(n_2617),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_3931),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4084),
.Y(n_4385)
);

OA22x2_ASAP7_75t_L g4386 ( 
.A1(n_4104),
.A2(n_956),
.B1(n_957),
.B2(n_952),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4118),
.Y(n_4387)
);

AND2x2_ASAP7_75t_SL g4388 ( 
.A(n_3970),
.B(n_956),
.Y(n_4388)
);

NOR2xp33_ASAP7_75t_L g4389 ( 
.A(n_3973),
.B(n_985),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_4031),
.A2(n_2645),
.B(n_2642),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_4032),
.A2(n_4058),
.B(n_3842),
.Y(n_4391)
);

O2A1O1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_3938),
.A2(n_958),
.B(n_959),
.C(n_957),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_SL g4393 ( 
.A(n_3797),
.B(n_2907),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_SL g4394 ( 
.A(n_3816),
.B(n_2907),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_3816),
.B(n_2907),
.Y(n_4395)
);

A2O1A1Ixp33_ASAP7_75t_L g4396 ( 
.A1(n_3978),
.A2(n_959),
.B(n_961),
.C(n_958),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4119),
.B(n_986),
.Y(n_4397)
);

OAI21x1_ASAP7_75t_L g4398 ( 
.A1(n_4129),
.A2(n_2677),
.B(n_2666),
.Y(n_4398)
);

A2O1A1Ixp33_ASAP7_75t_SL g4399 ( 
.A1(n_4097),
.A2(n_2645),
.B(n_2650),
.C(n_2642),
.Y(n_4399)
);

BUFx6f_ASAP7_75t_L g4400 ( 
.A(n_3895),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_3986),
.A2(n_2650),
.B(n_2645),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4085),
.A2(n_991),
.B1(n_993),
.B2(n_987),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_3805),
.B(n_995),
.Y(n_4403)
);

INVx4_ASAP7_75t_L g4404 ( 
.A(n_3895),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4073),
.Y(n_4405)
);

NOR2xp33_ASAP7_75t_L g4406 ( 
.A(n_4004),
.B(n_996),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_3805),
.A2(n_998),
.B1(n_999),
.B2(n_997),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4145),
.B(n_1000),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4161),
.B(n_1515),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_3809),
.B(n_1001),
.Y(n_4410)
);

OAI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_3969),
.A2(n_2652),
.B(n_2650),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4069),
.A2(n_2657),
.B(n_2652),
.Y(n_4412)
);

OAI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_3872),
.A2(n_3957),
.B1(n_4116),
.B2(n_4105),
.Y(n_4413)
);

AND2x4_ASAP7_75t_L g4414 ( 
.A(n_3832),
.B(n_2660),
.Y(n_4414)
);

BUFx2_ASAP7_75t_L g4415 ( 
.A(n_4015),
.Y(n_4415)
);

INVx5_ASAP7_75t_L g4416 ( 
.A(n_4015),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_3904),
.A2(n_3910),
.B(n_3857),
.Y(n_4417)
);

AOI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_3852),
.A2(n_2657),
.B(n_2652),
.Y(n_4418)
);

AOI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_3893),
.A2(n_2660),
.B(n_2657),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_SL g4420 ( 
.A(n_3872),
.B(n_2907),
.Y(n_4420)
);

INVx2_ASAP7_75t_SL g4421 ( 
.A(n_4015),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_3809),
.B(n_1005),
.Y(n_4422)
);

AOI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_3832),
.A2(n_3864),
.B1(n_4161),
.B2(n_3826),
.Y(n_4423)
);

INVx8_ASAP7_75t_L g4424 ( 
.A(n_4025),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4066),
.B(n_1006),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4025),
.Y(n_4426)
);

O2A1O1Ixp33_ASAP7_75t_L g4427 ( 
.A1(n_3974),
.A2(n_964),
.B(n_970),
.C(n_961),
.Y(n_4427)
);

OAI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_3957),
.A2(n_970),
.B1(n_972),
.B2(n_964),
.Y(n_4428)
);

O2A1O1Ixp33_ASAP7_75t_L g4429 ( 
.A1(n_3826),
.A2(n_977),
.B(n_981),
.C(n_972),
.Y(n_4429)
);

O2A1O1Ixp5_ASAP7_75t_L g4430 ( 
.A1(n_3995),
.A2(n_2662),
.B(n_2666),
.C(n_2660),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_SL g4431 ( 
.A(n_4051),
.B(n_4116),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4076),
.B(n_1009),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4080),
.B(n_4081),
.Y(n_4433)
);

AOI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_3864),
.A2(n_1012),
.B1(n_1014),
.B2(n_1011),
.Y(n_4434)
);

AOI33xp33_ASAP7_75t_L g4435 ( 
.A1(n_4054),
.A2(n_989),
.A3(n_981),
.B1(n_992),
.B2(n_988),
.B3(n_977),
.Y(n_4435)
);

AOI21xp5_ASAP7_75t_L g4436 ( 
.A1(n_3841),
.A2(n_2666),
.B(n_2662),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4114),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_3858),
.A2(n_2677),
.B(n_2662),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4098),
.B(n_1015),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_SL g4440 ( 
.A(n_3909),
.B(n_2697),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4106),
.B(n_1019),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_3917),
.B(n_3982),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_SL g4443 ( 
.A(n_3982),
.B(n_2677),
.Y(n_4443)
);

AND2x4_ASAP7_75t_L g4444 ( 
.A(n_3891),
.B(n_2679),
.Y(n_4444)
);

INVx4_ASAP7_75t_L g4445 ( 
.A(n_4025),
.Y(n_4445)
);

AOI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_3879),
.A2(n_2681),
.B(n_2679),
.Y(n_4446)
);

AOI21x1_ASAP7_75t_L g4447 ( 
.A1(n_4006),
.A2(n_2681),
.B(n_2679),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4130),
.Y(n_4448)
);

OAI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_3913),
.A2(n_2685),
.B(n_2681),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4157),
.B(n_1519),
.Y(n_4450)
);

AOI22xp33_ASAP7_75t_L g4451 ( 
.A1(n_3891),
.A2(n_837),
.B1(n_920),
.B2(n_824),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4109),
.B(n_1020),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4153),
.Y(n_4453)
);

BUFx6f_ASAP7_75t_L g4454 ( 
.A(n_4029),
.Y(n_4454)
);

AND2x4_ASAP7_75t_L g4455 ( 
.A(n_4010),
.B(n_2695),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4115),
.B(n_1024),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_SL g4457 ( 
.A(n_4128),
.B(n_946),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_3984),
.B(n_4110),
.Y(n_4458)
);

AND2x4_ASAP7_75t_L g4459 ( 
.A(n_4010),
.B(n_2697),
.Y(n_4459)
);

BUFx2_ASAP7_75t_L g4460 ( 
.A(n_4029),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4133),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4133),
.Y(n_4462)
);

AOI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_4148),
.A2(n_4156),
.B1(n_4123),
.B2(n_4057),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_3988),
.B(n_1027),
.Y(n_4464)
);

AND2x4_ASAP7_75t_L g4465 ( 
.A(n_4128),
.B(n_2698),
.Y(n_4465)
);

CKINVDCx20_ASAP7_75t_R g4466 ( 
.A(n_4029),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3988),
.B(n_1030),
.Y(n_4467)
);

BUFx6f_ASAP7_75t_L g4468 ( 
.A(n_4090),
.Y(n_4468)
);

NOR2xp33_ASAP7_75t_L g4469 ( 
.A(n_4056),
.B(n_1033),
.Y(n_4469)
);

INVx2_ASAP7_75t_SL g4470 ( 
.A(n_4090),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_3979),
.B(n_2685),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4090),
.B(n_1520),
.Y(n_4472)
);

NAND2x1p5_ASAP7_75t_L g4473 ( 
.A(n_4087),
.B(n_2685),
.Y(n_4473)
);

INVx1_ASAP7_75t_SL g4474 ( 
.A(n_4138),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_3961),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_3989),
.B(n_1036),
.Y(n_4476)
);

NOR2xp33_ASAP7_75t_L g4477 ( 
.A(n_4087),
.B(n_1039),
.Y(n_4477)
);

O2A1O1Ixp33_ASAP7_75t_L g4478 ( 
.A1(n_4131),
.A2(n_989),
.B(n_992),
.C(n_988),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_3996),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4117),
.B(n_1522),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_4100),
.A2(n_1045),
.B1(n_1048),
.B2(n_1043),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_SL g4482 ( 
.A(n_4070),
.B(n_2686),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_3989),
.B(n_1051),
.Y(n_4483)
);

O2A1O1Ixp33_ASAP7_75t_L g4484 ( 
.A1(n_4143),
.A2(n_1007),
.B(n_1016),
.C(n_994),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_3990),
.B(n_1053),
.Y(n_4485)
);

AOI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_3810),
.A2(n_2690),
.B(n_2686),
.Y(n_4486)
);

AOI21xp5_ASAP7_75t_L g4487 ( 
.A1(n_4061),
.A2(n_2690),
.B(n_2686),
.Y(n_4487)
);

OAI22xp5_ASAP7_75t_L g4488 ( 
.A1(n_4103),
.A2(n_1070),
.B1(n_1071),
.B2(n_1055),
.Y(n_4488)
);

NOR2xp33_ASAP7_75t_R g4489 ( 
.A(n_4117),
.B(n_1074),
.Y(n_4489)
);

AOI21xp5_ASAP7_75t_L g4490 ( 
.A1(n_4011),
.A2(n_2695),
.B(n_2690),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_4020),
.A2(n_2697),
.B(n_2695),
.Y(n_4491)
);

O2A1O1Ixp5_ASAP7_75t_L g4492 ( 
.A1(n_3981),
.A2(n_2703),
.B(n_2698),
.C(n_2507),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_4055),
.A2(n_2703),
.B(n_2698),
.Y(n_4493)
);

AO22x1_ASAP7_75t_L g4494 ( 
.A1(n_4089),
.A2(n_1077),
.B1(n_1078),
.B2(n_1076),
.Y(n_4494)
);

OAI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_4121),
.A2(n_2703),
.B(n_2507),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_3990),
.B(n_1080),
.Y(n_4496)
);

BUFx8_ASAP7_75t_L g4497 ( 
.A(n_4117),
.Y(n_4497)
);

BUFx8_ASAP7_75t_SL g4498 ( 
.A(n_4127),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4048),
.B(n_1081),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_3916),
.A2(n_2507),
.B(n_2500),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4122),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_3947),
.Y(n_4502)
);

A2O1A1Ixp33_ASAP7_75t_L g4503 ( 
.A1(n_3959),
.A2(n_1007),
.B(n_1016),
.C(n_994),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_SL g4504 ( 
.A(n_3939),
.B(n_837),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4005),
.B(n_1083),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_SL g4506 ( 
.A(n_3940),
.B(n_837),
.Y(n_4506)
);

AOI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_3918),
.A2(n_2511),
.B(n_2500),
.Y(n_4507)
);

OAI22xp5_ASAP7_75t_L g4508 ( 
.A1(n_4103),
.A2(n_1035),
.B1(n_1037),
.B2(n_1025),
.Y(n_4508)
);

INVx3_ASAP7_75t_L g4509 ( 
.A(n_4127),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4017),
.B(n_1086),
.Y(n_4510)
);

AOI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_4105),
.A2(n_2511),
.B(n_2500),
.Y(n_4511)
);

AOI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_4125),
.A2(n_2513),
.B(n_2511),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_3947),
.Y(n_4513)
);

BUFx2_ASAP7_75t_L g4514 ( 
.A(n_4127),
.Y(n_4514)
);

O2A1O1Ixp5_ASAP7_75t_L g4515 ( 
.A1(n_3900),
.A2(n_2518),
.B(n_2520),
.C(n_2513),
.Y(n_4515)
);

NOR3xp33_ASAP7_75t_L g4516 ( 
.A(n_4144),
.B(n_1528),
.C(n_1523),
.Y(n_4516)
);

O2A1O1Ixp33_ASAP7_75t_L g4517 ( 
.A1(n_4151),
.A2(n_1035),
.B(n_1037),
.C(n_1025),
.Y(n_4517)
);

A2O1A1Ixp33_ASAP7_75t_L g4518 ( 
.A1(n_3966),
.A2(n_1052),
.B(n_1054),
.C(n_1038),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4030),
.B(n_4037),
.Y(n_4519)
);

AOI22x1_ASAP7_75t_L g4520 ( 
.A1(n_3907),
.A2(n_2518),
.B1(n_2520),
.B2(n_2513),
.Y(n_4520)
);

CKINVDCx5p33_ASAP7_75t_R g4521 ( 
.A(n_4155),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4039),
.B(n_1089),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_4125),
.A2(n_2520),
.B(n_2518),
.Y(n_4523)
);

BUFx2_ASAP7_75t_L g4524 ( 
.A(n_4155),
.Y(n_4524)
);

NOR2xp33_ASAP7_75t_SL g4525 ( 
.A(n_3898),
.B(n_946),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_3901),
.A2(n_2568),
.B(n_2522),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4013),
.B(n_1092),
.Y(n_4527)
);

NAND2xp33_ASAP7_75t_L g4528 ( 
.A(n_4155),
.B(n_1094),
.Y(n_4528)
);

NOR2xp33_ASAP7_75t_L g4529 ( 
.A(n_4138),
.B(n_1095),
.Y(n_4529)
);

NOR2x1_ASAP7_75t_R g4530 ( 
.A(n_4154),
.B(n_1096),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_3949),
.Y(n_4531)
);

BUFx8_ASAP7_75t_L g4532 ( 
.A(n_3949),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4013),
.B(n_1098),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_3951),
.B(n_837),
.Y(n_4534)
);

NOR2xp67_ASAP7_75t_SL g4535 ( 
.A(n_3971),
.B(n_1038),
.Y(n_4535)
);

BUFx2_ASAP7_75t_L g4536 ( 
.A(n_4102),
.Y(n_4536)
);

AOI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_3902),
.A2(n_2568),
.B(n_2522),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_3912),
.A2(n_2568),
.B(n_2522),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4014),
.B(n_4036),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_SL g4540 ( 
.A(n_3977),
.B(n_920),
.Y(n_4540)
);

OAI22x1_ASAP7_75t_L g4541 ( 
.A1(n_3907),
.A2(n_1054),
.B1(n_1060),
.B2(n_1052),
.Y(n_4541)
);

AOI22xp5_ASAP7_75t_L g4542 ( 
.A1(n_3923),
.A2(n_4122),
.B1(n_4014),
.B2(n_1104),
.Y(n_4542)
);

BUFx4f_ASAP7_75t_L g4543 ( 
.A(n_4102),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4134),
.B(n_1101),
.Y(n_4544)
);

INVx6_ASAP7_75t_L g4545 ( 
.A(n_3898),
.Y(n_4545)
);

OAI22xp5_ASAP7_75t_L g4546 ( 
.A1(n_4158),
.A2(n_1065),
.B1(n_1066),
.B2(n_1060),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_4134),
.B(n_4136),
.Y(n_4547)
);

AOI21xp5_ASAP7_75t_L g4548 ( 
.A1(n_4075),
.A2(n_4101),
.B(n_4150),
.Y(n_4548)
);

OAI321xp33_ASAP7_75t_L g4549 ( 
.A1(n_3923),
.A2(n_1072),
.A3(n_1066),
.B1(n_1073),
.B2(n_1067),
.C(n_1065),
.Y(n_4549)
);

AOI33xp33_ASAP7_75t_L g4550 ( 
.A1(n_4142),
.A2(n_1079),
.A3(n_1072),
.B1(n_1084),
.B2(n_1073),
.B3(n_1067),
.Y(n_4550)
);

OAI21x1_ASAP7_75t_L g4551 ( 
.A1(n_3964),
.A2(n_2570),
.B(n_2569),
.Y(n_4551)
);

AOI21xp5_ASAP7_75t_L g4552 ( 
.A1(n_4112),
.A2(n_2570),
.B(n_2569),
.Y(n_4552)
);

BUFx6f_ASAP7_75t_L g4553 ( 
.A(n_4159),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4136),
.B(n_4141),
.Y(n_4554)
);

OAI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4113),
.A2(n_1084),
.B1(n_1085),
.B2(n_1079),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4088),
.B(n_1107),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_L g4557 ( 
.A(n_4093),
.B(n_1108),
.Y(n_4557)
);

AOI21x1_ASAP7_75t_L g4558 ( 
.A1(n_4132),
.A2(n_2461),
.B(n_2454),
.Y(n_4558)
);

AOI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_4162),
.A2(n_2570),
.B(n_2569),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4107),
.Y(n_4560)
);

AO22x1_ASAP7_75t_L g4561 ( 
.A1(n_4163),
.A2(n_1113),
.B1(n_1114),
.B2(n_1110),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_4163),
.A2(n_2577),
.B(n_2571),
.Y(n_4562)
);

AOI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_3788),
.A2(n_1129),
.B1(n_1130),
.B2(n_1121),
.Y(n_4563)
);

AOI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_3791),
.A2(n_2577),
.B(n_2571),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_3791),
.A2(n_2577),
.B(n_2571),
.Y(n_4565)
);

NOR2xp33_ASAP7_75t_L g4566 ( 
.A(n_3863),
.B(n_1136),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4236),
.B(n_1085),
.Y(n_4567)
);

BUFx2_ASAP7_75t_L g4568 ( 
.A(n_4466),
.Y(n_4568)
);

OAI21x1_ASAP7_75t_SL g4569 ( 
.A1(n_4341),
.A2(n_1103),
.B(n_1087),
.Y(n_4569)
);

NOR2xp67_ASAP7_75t_L g4570 ( 
.A(n_4189),
.B(n_1530),
.Y(n_4570)
);

AND2x4_ASAP7_75t_L g4571 ( 
.A(n_4244),
.B(n_2449),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4172),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_SL g4573 ( 
.A(n_4184),
.B(n_1625),
.Y(n_4573)
);

OAI21x1_ASAP7_75t_L g4574 ( 
.A1(n_4417),
.A2(n_2062),
.B(n_2057),
.Y(n_4574)
);

AOI221xp5_ASAP7_75t_SL g4575 ( 
.A1(n_4318),
.A2(n_4410),
.B1(n_4422),
.B2(n_4403),
.C(n_4428),
.Y(n_4575)
);

AOI21x1_ASAP7_75t_L g4576 ( 
.A1(n_4494),
.A2(n_1637),
.B(n_1629),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4226),
.Y(n_4577)
);

AOI21x1_ASAP7_75t_SL g4578 ( 
.A1(n_4328),
.A2(n_931),
.B(n_920),
.Y(n_4578)
);

AOI21xp5_ASAP7_75t_SL g4579 ( 
.A1(n_4168),
.A2(n_4310),
.B(n_4530),
.Y(n_4579)
);

OAI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4243),
.A2(n_2463),
.B(n_2461),
.Y(n_4580)
);

OAI21x1_ASAP7_75t_L g4581 ( 
.A1(n_4391),
.A2(n_2062),
.B(n_2057),
.Y(n_4581)
);

NOR2x1_ASAP7_75t_L g4582 ( 
.A(n_4208),
.B(n_1087),
.Y(n_4582)
);

INVxp67_ASAP7_75t_L g4583 ( 
.A(n_4238),
.Y(n_4583)
);

OAI22xp5_ASAP7_75t_L g4584 ( 
.A1(n_4197),
.A2(n_1105),
.B1(n_1118),
.B2(n_1103),
.Y(n_4584)
);

INVx1_ASAP7_75t_SL g4585 ( 
.A(n_4315),
.Y(n_4585)
);

AOI21xp5_ASAP7_75t_L g4586 ( 
.A1(n_4167),
.A2(n_2070),
.B(n_2069),
.Y(n_4586)
);

AOI21xp5_ASAP7_75t_L g4587 ( 
.A1(n_4548),
.A2(n_2070),
.B(n_2069),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4371),
.B(n_1629),
.Y(n_4588)
);

OAI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4175),
.A2(n_2464),
.B(n_2463),
.Y(n_4589)
);

BUFx3_ASAP7_75t_L g4590 ( 
.A(n_4349),
.Y(n_4590)
);

AOI21x1_ASAP7_75t_SL g4591 ( 
.A1(n_4331),
.A2(n_931),
.B(n_920),
.Y(n_4591)
);

OAI21x1_ASAP7_75t_L g4592 ( 
.A1(n_4199),
.A2(n_2075),
.B(n_2071),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4219),
.B(n_1137),
.Y(n_4593)
);

INVx2_ASAP7_75t_SL g4594 ( 
.A(n_4349),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4206),
.B(n_1637),
.Y(n_4595)
);

AOI221x1_ASAP7_75t_L g4596 ( 
.A1(n_4406),
.A2(n_1119),
.B1(n_1124),
.B2(n_1118),
.C(n_1105),
.Y(n_4596)
);

OAI21x1_ASAP7_75t_L g4597 ( 
.A1(n_4447),
.A2(n_2075),
.B(n_2071),
.Y(n_4597)
);

CKINVDCx5p33_ASAP7_75t_R g4598 ( 
.A(n_4214),
.Y(n_4598)
);

OA22x2_ASAP7_75t_L g4599 ( 
.A1(n_4423),
.A2(n_1124),
.B1(n_1128),
.B2(n_1119),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4281),
.Y(n_4600)
);

NOR2x1_ASAP7_75t_SL g4601 ( 
.A(n_4267),
.B(n_2464),
.Y(n_4601)
);

BUFx6f_ASAP7_75t_L g4602 ( 
.A(n_4186),
.Y(n_4602)
);

A2O1A1Ixp33_ASAP7_75t_L g4603 ( 
.A1(n_4469),
.A2(n_1132),
.B(n_1133),
.C(n_1128),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4220),
.B(n_1640),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4284),
.Y(n_4605)
);

BUFx4f_ASAP7_75t_L g4606 ( 
.A(n_4289),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4165),
.B(n_1139),
.Y(n_4607)
);

AO31x2_ASAP7_75t_L g4608 ( 
.A1(n_4287),
.A2(n_2088),
.A3(n_2090),
.B(n_2077),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_SL g4609 ( 
.A(n_4213),
.B(n_1640),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4212),
.B(n_1142),
.Y(n_4610)
);

NAND2x1p5_ASAP7_75t_L g4611 ( 
.A(n_4267),
.B(n_2077),
.Y(n_4611)
);

OR2x2_ASAP7_75t_L g4612 ( 
.A(n_4474),
.B(n_1647),
.Y(n_4612)
);

NOR2xp33_ASAP7_75t_L g4613 ( 
.A(n_4245),
.B(n_1151),
.Y(n_4613)
);

NOR3xp33_ASAP7_75t_L g4614 ( 
.A(n_4346),
.B(n_1535),
.C(n_1532),
.Y(n_4614)
);

AO31x2_ASAP7_75t_L g4615 ( 
.A1(n_4479),
.A2(n_2090),
.A3(n_2102),
.B(n_2088),
.Y(n_4615)
);

INVx3_ASAP7_75t_L g4616 ( 
.A(n_4308),
.Y(n_4616)
);

OA22x2_ASAP7_75t_L g4617 ( 
.A1(n_4194),
.A2(n_1133),
.B1(n_1134),
.B2(n_1132),
.Y(n_4617)
);

OAI21x1_ASAP7_75t_L g4618 ( 
.A1(n_4322),
.A2(n_2108),
.B(n_2102),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4409),
.B(n_1647),
.Y(n_4619)
);

NOR2x1_ASAP7_75t_L g4620 ( 
.A(n_4224),
.B(n_1134),
.Y(n_4620)
);

OAI21x1_ASAP7_75t_L g4621 ( 
.A1(n_4215),
.A2(n_2110),
.B(n_2108),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_SL g4622 ( 
.A(n_4213),
.B(n_1649),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_SL g4623 ( 
.A(n_4210),
.B(n_1649),
.Y(n_4623)
);

OAI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4556),
.A2(n_4557),
.B(n_4255),
.Y(n_4624)
);

OAI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4431),
.A2(n_2473),
.B(n_2465),
.Y(n_4625)
);

NOR2xp33_ASAP7_75t_L g4626 ( 
.A(n_4309),
.B(n_1155),
.Y(n_4626)
);

O2A1O1Ixp5_ASAP7_75t_SL g4627 ( 
.A1(n_4504),
.A2(n_1141),
.B(n_1146),
.C(n_1138),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4195),
.Y(n_4628)
);

AND2x4_ASAP7_75t_L g4629 ( 
.A(n_4244),
.B(n_4280),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_SL g4630 ( 
.A(n_4202),
.B(n_1650),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4272),
.B(n_1138),
.Y(n_4631)
);

OR2x6_ASAP7_75t_L g4632 ( 
.A(n_4179),
.B(n_2110),
.Y(n_4632)
);

NOR2xp33_ASAP7_75t_L g4633 ( 
.A(n_4253),
.B(n_1159),
.Y(n_4633)
);

OA21x2_ASAP7_75t_L g4634 ( 
.A1(n_4430),
.A2(n_1597),
.B(n_1596),
.Y(n_4634)
);

OR2x6_ASAP7_75t_L g4635 ( 
.A(n_4177),
.B(n_2116),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4529),
.B(n_1650),
.Y(n_4636)
);

OAI21xp5_ASAP7_75t_L g4637 ( 
.A1(n_4181),
.A2(n_2473),
.B(n_2465),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4272),
.B(n_1141),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4216),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4539),
.B(n_1146),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4474),
.B(n_1147),
.Y(n_4641)
);

OAI21x1_ASAP7_75t_L g4642 ( 
.A1(n_4398),
.A2(n_2128),
.B(n_2116),
.Y(n_4642)
);

AO31x2_ASAP7_75t_L g4643 ( 
.A1(n_4413),
.A2(n_2130),
.A3(n_2141),
.B(n_2128),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4186),
.Y(n_4644)
);

AO31x2_ASAP7_75t_L g4645 ( 
.A1(n_4413),
.A2(n_4270),
.A3(n_4555),
.B(n_4560),
.Y(n_4645)
);

OAI21x1_ASAP7_75t_L g4646 ( 
.A1(n_4500),
.A2(n_2141),
.B(n_2130),
.Y(n_4646)
);

INVx5_ASAP7_75t_L g4647 ( 
.A(n_4296),
.Y(n_4647)
);

AO31x2_ASAP7_75t_L g4648 ( 
.A1(n_4270),
.A2(n_2143),
.A3(n_2148),
.B(n_2142),
.Y(n_4648)
);

AOI221x1_ASAP7_75t_L g4649 ( 
.A1(n_4428),
.A2(n_1152),
.B1(n_1158),
.B2(n_1150),
.C(n_1147),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4298),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4217),
.Y(n_4651)
);

OAI21x1_ASAP7_75t_L g4652 ( 
.A1(n_4507),
.A2(n_2143),
.B(n_2142),
.Y(n_4652)
);

OAI21x1_ASAP7_75t_SL g4653 ( 
.A1(n_4265),
.A2(n_1152),
.B(n_1150),
.Y(n_4653)
);

OAI21xp5_ASAP7_75t_L g4654 ( 
.A1(n_4475),
.A2(n_4203),
.B(n_4233),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4394),
.A2(n_2168),
.B(n_2148),
.Y(n_4655)
);

OAI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4242),
.A2(n_2478),
.B(n_2186),
.Y(n_4656)
);

INVx4_ASAP7_75t_L g4657 ( 
.A(n_4289),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4201),
.B(n_1161),
.Y(n_4658)
);

OAI21x1_ASAP7_75t_L g4659 ( 
.A1(n_4486),
.A2(n_2186),
.B(n_2168),
.Y(n_4659)
);

AND2x4_ASAP7_75t_L g4660 ( 
.A(n_4280),
.B(n_2449),
.Y(n_4660)
);

BUFx12f_ASAP7_75t_L g4661 ( 
.A(n_4187),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4519),
.B(n_1168),
.Y(n_4662)
);

BUFx6f_ASAP7_75t_L g4663 ( 
.A(n_4186),
.Y(n_4663)
);

OAI21x1_ASAP7_75t_L g4664 ( 
.A1(n_4401),
.A2(n_2194),
.B(n_2192),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4363),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_4289),
.Y(n_4666)
);

AOI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_4395),
.A2(n_2194),
.B(n_2192),
.Y(n_4667)
);

AOI21x1_ASAP7_75t_L g4668 ( 
.A1(n_4535),
.A2(n_4555),
.B(n_4534),
.Y(n_4668)
);

OAI21x1_ASAP7_75t_L g4669 ( 
.A1(n_4305),
.A2(n_2198),
.B(n_2196),
.Y(n_4669)
);

INVx2_ASAP7_75t_SL g4670 ( 
.A(n_4176),
.Y(n_4670)
);

OAI21x1_ASAP7_75t_SL g4671 ( 
.A1(n_4429),
.A2(n_1160),
.B(n_1158),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4372),
.A2(n_2198),
.B(n_2196),
.Y(n_4672)
);

INVx1_ASAP7_75t_SL g4673 ( 
.A(n_4458),
.Y(n_4673)
);

OAI21x1_ASAP7_75t_L g4674 ( 
.A1(n_4538),
.A2(n_2209),
.B(n_2204),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_L g4675 ( 
.A(n_4277),
.B(n_1169),
.Y(n_4675)
);

AOI221x1_ASAP7_75t_L g4676 ( 
.A1(n_4541),
.A2(n_1166),
.B1(n_1167),
.B2(n_1165),
.C(n_1160),
.Y(n_4676)
);

OAI21x1_ASAP7_75t_L g4677 ( 
.A1(n_4449),
.A2(n_2209),
.B(n_2204),
.Y(n_4677)
);

AOI31xp67_ASAP7_75t_L g4678 ( 
.A1(n_4202),
.A2(n_2220),
.A3(n_2222),
.B(n_2214),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4170),
.B(n_1170),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4385),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_4282),
.Y(n_4681)
);

AOI21xp5_ASAP7_75t_L g4682 ( 
.A1(n_4393),
.A2(n_2220),
.B(n_2214),
.Y(n_4682)
);

OAI21x1_ASAP7_75t_L g4683 ( 
.A1(n_4449),
.A2(n_2230),
.B(n_2222),
.Y(n_4683)
);

INVxp67_ASAP7_75t_SL g4684 ( 
.A(n_4178),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4408),
.B(n_1173),
.Y(n_4685)
);

CKINVDCx11_ASAP7_75t_R g4686 ( 
.A(n_4263),
.Y(n_4686)
);

INVx3_ASAP7_75t_SL g4687 ( 
.A(n_4339),
.Y(n_4687)
);

OAI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4478),
.A2(n_2478),
.B(n_2245),
.Y(n_4688)
);

AOI21xp5_ASAP7_75t_L g4689 ( 
.A1(n_4420),
.A2(n_2245),
.B(n_2230),
.Y(n_4689)
);

AO31x2_ASAP7_75t_L g4690 ( 
.A1(n_4501),
.A2(n_4274),
.A3(n_4283),
.B(n_4249),
.Y(n_4690)
);

OAI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4484),
.A2(n_2249),
.B(n_2248),
.Y(n_4691)
);

OAI21xp5_ASAP7_75t_L g4692 ( 
.A1(n_4517),
.A2(n_2249),
.B(n_2248),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4180),
.B(n_1175),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4228),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4387),
.Y(n_4695)
);

OAI22xp5_ASAP7_75t_L g4696 ( 
.A1(n_4197),
.A2(n_1166),
.B1(n_1167),
.B2(n_1165),
.Y(n_4696)
);

O2A1O1Ixp5_ASAP7_75t_L g4697 ( 
.A1(n_4561),
.A2(n_1178),
.B(n_1179),
.C(n_1174),
.Y(n_4697)
);

OAI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4516),
.A2(n_2261),
.B(n_2250),
.Y(n_4698)
);

OAI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4362),
.A2(n_2261),
.B(n_2250),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4544),
.B(n_1177),
.Y(n_4700)
);

OAI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4324),
.A2(n_2275),
.B(n_2262),
.Y(n_4701)
);

INVx2_ASAP7_75t_SL g4702 ( 
.A(n_4237),
.Y(n_4702)
);

AOI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4241),
.A2(n_2275),
.B(n_2262),
.Y(n_4703)
);

AOI21xp5_ASAP7_75t_L g4704 ( 
.A1(n_4241),
.A2(n_2302),
.B(n_2299),
.Y(n_4704)
);

AO21x2_ASAP7_75t_L g4705 ( 
.A1(n_4558),
.A2(n_4380),
.B(n_4218),
.Y(n_4705)
);

AOI221xp5_ASAP7_75t_SL g4706 ( 
.A1(n_4260),
.A2(n_1179),
.B1(n_1191),
.B2(n_1178),
.C(n_1174),
.Y(n_4706)
);

AO31x2_ASAP7_75t_L g4707 ( 
.A1(n_4274),
.A2(n_2302),
.A3(n_2311),
.B(n_2299),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4360),
.Y(n_4708)
);

OAI21x1_ASAP7_75t_L g4709 ( 
.A1(n_4326),
.A2(n_2314),
.B(n_2311),
.Y(n_4709)
);

OAI21x1_ASAP7_75t_L g4710 ( 
.A1(n_4327),
.A2(n_2315),
.B(n_2314),
.Y(n_4710)
);

NOR2x1_ASAP7_75t_SL g4711 ( 
.A(n_4267),
.B(n_2315),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4336),
.A2(n_2333),
.B(n_2319),
.Y(n_4712)
);

AOI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4442),
.A2(n_2333),
.B(n_2319),
.Y(n_4713)
);

INVx2_ASAP7_75t_SL g4714 ( 
.A(n_4237),
.Y(n_4714)
);

OAI22xp5_ASAP7_75t_L g4715 ( 
.A1(n_4407),
.A2(n_1198),
.B1(n_1210),
.B2(n_1191),
.Y(n_4715)
);

OAI22x1_ASAP7_75t_L g4716 ( 
.A1(n_4463),
.A2(n_1210),
.B1(n_1216),
.B2(n_1198),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4173),
.B(n_1180),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4240),
.B(n_1653),
.Y(n_4718)
);

OR2x6_ASAP7_75t_L g4719 ( 
.A(n_4296),
.B(n_2349),
.Y(n_4719)
);

INVx5_ASAP7_75t_L g4720 ( 
.A(n_4296),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4461),
.B(n_1216),
.Y(n_4721)
);

OAI21x1_ASAP7_75t_L g4722 ( 
.A1(n_4329),
.A2(n_2353),
.B(n_2349),
.Y(n_4722)
);

BUFx6f_ASAP7_75t_L g4723 ( 
.A(n_4400),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4543),
.A2(n_2355),
.B(n_2353),
.Y(n_4724)
);

A2O1A1Ixp33_ASAP7_75t_L g4725 ( 
.A1(n_4188),
.A2(n_1220),
.B(n_1222),
.C(n_1217),
.Y(n_4725)
);

A2O1A1Ixp33_ASAP7_75t_L g4726 ( 
.A1(n_4330),
.A2(n_1220),
.B(n_1222),
.C(n_1217),
.Y(n_4726)
);

AOI21x1_ASAP7_75t_L g4727 ( 
.A1(n_4506),
.A2(n_1655),
.B(n_1653),
.Y(n_4727)
);

OAI21xp5_ASAP7_75t_L g4728 ( 
.A1(n_4542),
.A2(n_2356),
.B(n_2355),
.Y(n_4728)
);

INVx1_ASAP7_75t_SL g4729 ( 
.A(n_4276),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_SL g4730 ( 
.A(n_4388),
.B(n_1655),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_SL g4731 ( 
.A1(n_4317),
.A2(n_2366),
.B(n_2356),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4462),
.B(n_1228),
.Y(n_4732)
);

HB1xp67_ASAP7_75t_L g4733 ( 
.A(n_4235),
.Y(n_4733)
);

INVx5_ASAP7_75t_L g4734 ( 
.A(n_4333),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4521),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_SL g4736 ( 
.A(n_4325),
.B(n_4262),
.Y(n_4736)
);

OAI22xp5_ASAP7_75t_L g4737 ( 
.A1(n_4171),
.A2(n_1230),
.B1(n_1232),
.B2(n_1228),
.Y(n_4737)
);

AOI21x1_ASAP7_75t_L g4738 ( 
.A1(n_4540),
.A2(n_1660),
.B(n_1658),
.Y(n_4738)
);

OAI21x1_ASAP7_75t_SL g4739 ( 
.A1(n_4367),
.A2(n_1232),
.B(n_1230),
.Y(n_4739)
);

INVx2_ASAP7_75t_SL g4740 ( 
.A(n_4301),
.Y(n_4740)
);

AO31x2_ASAP7_75t_L g4741 ( 
.A1(n_4283),
.A2(n_2371),
.A3(n_2377),
.B(n_2366),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4257),
.B(n_1658),
.Y(n_4742)
);

NOR2x1_ASAP7_75t_SL g4743 ( 
.A(n_4267),
.B(n_2371),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4547),
.B(n_1237),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4261),
.B(n_1237),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4227),
.B(n_1238),
.Y(n_4746)
);

AND2x2_ASAP7_75t_L g4747 ( 
.A(n_4278),
.B(n_1660),
.Y(n_4747)
);

AOI21xp33_ASAP7_75t_L g4748 ( 
.A1(n_4392),
.A2(n_4427),
.B(n_4566),
.Y(n_4748)
);

AOI21xp5_ASAP7_75t_L g4749 ( 
.A1(n_4543),
.A2(n_2379),
.B(n_2377),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4231),
.B(n_1238),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4293),
.B(n_1239),
.Y(n_4751)
);

BUFx2_ASAP7_75t_L g4752 ( 
.A(n_4182),
.Y(n_4752)
);

AOI21xp5_ASAP7_75t_L g4753 ( 
.A1(n_4292),
.A2(n_2385),
.B(n_2379),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4303),
.B(n_1182),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4299),
.B(n_1239),
.Y(n_4755)
);

OR2x6_ASAP7_75t_L g4756 ( 
.A(n_4268),
.B(n_4264),
.Y(n_4756)
);

NOR2xp33_ASAP7_75t_L g4757 ( 
.A(n_4347),
.B(n_1183),
.Y(n_4757)
);

NAND3xp33_ASAP7_75t_L g4758 ( 
.A(n_4273),
.B(n_1185),
.C(n_1184),
.Y(n_4758)
);

NOR2xp67_ASAP7_75t_SL g4759 ( 
.A(n_4339),
.B(n_1537),
.Y(n_4759)
);

OAI21x1_ASAP7_75t_L g4760 ( 
.A1(n_4354),
.A2(n_4379),
.B(n_4356),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4256),
.Y(n_4761)
);

BUFx4_ASAP7_75t_SL g4762 ( 
.A(n_4353),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4448),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_L g4764 ( 
.A(n_4191),
.B(n_1242),
.Y(n_4764)
);

OAI21x1_ASAP7_75t_L g4765 ( 
.A1(n_4390),
.A2(n_2390),
.B(n_2385),
.Y(n_4765)
);

AOI21xp5_ASAP7_75t_L g4766 ( 
.A1(n_4554),
.A2(n_2392),
.B(n_2390),
.Y(n_4766)
);

OAI21x1_ASAP7_75t_L g4767 ( 
.A1(n_4223),
.A2(n_2400),
.B(n_2392),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4351),
.B(n_1662),
.Y(n_4768)
);

OAI21x1_ASAP7_75t_L g4769 ( 
.A1(n_4436),
.A2(n_2401),
.B(n_2400),
.Y(n_4769)
);

BUFx6f_ASAP7_75t_L g4770 ( 
.A(n_4400),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4472),
.B(n_1662),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4453),
.Y(n_4772)
);

OAI21x1_ASAP7_75t_L g4773 ( 
.A1(n_4564),
.A2(n_2418),
.B(n_2401),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4450),
.B(n_1190),
.Y(n_4774)
);

OAI21x1_ASAP7_75t_L g4775 ( 
.A1(n_4565),
.A2(n_2433),
.B(n_2418),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4271),
.Y(n_4776)
);

NOR2xp33_ASAP7_75t_SL g4777 ( 
.A(n_4457),
.B(n_931),
.Y(n_4777)
);

NOR2xp33_ASAP7_75t_SL g4778 ( 
.A(n_4457),
.B(n_931),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4396),
.A2(n_2447),
.B(n_2433),
.Y(n_4779)
);

BUFx3_ASAP7_75t_L g4780 ( 
.A(n_4498),
.Y(n_4780)
);

CKINVDCx16_ASAP7_75t_R g4781 ( 
.A(n_4234),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4464),
.B(n_1195),
.Y(n_4782)
);

NAND2x1p5_ASAP7_75t_L g4783 ( 
.A(n_4252),
.B(n_4531),
.Y(n_4783)
);

OAI21xp33_ASAP7_75t_L g4784 ( 
.A1(n_4435),
.A2(n_1199),
.B(n_1196),
.Y(n_4784)
);

INVx2_ASAP7_75t_SL g4785 ( 
.A(n_4359),
.Y(n_4785)
);

AND2x2_ASAP7_75t_SL g4786 ( 
.A(n_4525),
.B(n_1242),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4482),
.A2(n_2452),
.B(n_2447),
.Y(n_4787)
);

BUFx3_ASAP7_75t_L g4788 ( 
.A(n_4384),
.Y(n_4788)
);

OAI21x1_ASAP7_75t_L g4789 ( 
.A1(n_4316),
.A2(n_2453),
.B(n_2452),
.Y(n_4789)
);

A2O1A1Ixp33_ASAP7_75t_L g4790 ( 
.A1(n_4373),
.A2(n_1250),
.B(n_1665),
.C(n_1663),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4209),
.B(n_1663),
.Y(n_4791)
);

OAI21x1_ASAP7_75t_L g4792 ( 
.A1(n_4493),
.A2(n_2453),
.B(n_2294),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4304),
.Y(n_4793)
);

OAI21x1_ASAP7_75t_L g4794 ( 
.A1(n_4490),
.A2(n_2294),
.B(n_2277),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4288),
.B(n_1665),
.Y(n_4795)
);

AOI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4246),
.A2(n_2294),
.B(n_2277),
.Y(n_4796)
);

OA21x2_ASAP7_75t_L g4797 ( 
.A1(n_4380),
.A2(n_1598),
.B(n_1597),
.Y(n_4797)
);

OA21x2_ASAP7_75t_L g4798 ( 
.A1(n_4411),
.A2(n_1599),
.B(n_1598),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4266),
.B(n_1666),
.Y(n_4799)
);

INVx5_ASAP7_75t_L g4800 ( 
.A(n_4333),
.Y(n_4800)
);

AND3x2_ASAP7_75t_L g4801 ( 
.A(n_4234),
.B(n_1540),
.C(n_1539),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4246),
.A2(n_2294),
.B(n_2277),
.Y(n_4802)
);

OAI21x1_ASAP7_75t_L g4803 ( 
.A1(n_4491),
.A2(n_2312),
.B(n_2308),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4314),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_4480),
.B(n_1666),
.Y(n_4805)
);

OAI21xp33_ASAP7_75t_L g4806 ( 
.A1(n_4364),
.A2(n_1207),
.B(n_1202),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_4286),
.B(n_1208),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4467),
.B(n_1211),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4487),
.A2(n_4383),
.B(n_4254),
.Y(n_4809)
);

INVx4_ASAP7_75t_L g4810 ( 
.A(n_4343),
.Y(n_4810)
);

OAI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4377),
.A2(n_1669),
.B(n_1668),
.Y(n_4811)
);

AOI21xp5_ASAP7_75t_SL g4812 ( 
.A1(n_4229),
.A2(n_4222),
.B(n_4476),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4335),
.Y(n_4813)
);

INVxp67_ASAP7_75t_SL g4814 ( 
.A(n_4196),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4313),
.A2(n_1213),
.B1(n_1214),
.B2(n_1212),
.Y(n_4815)
);

INVx1_ASAP7_75t_SL g4816 ( 
.A(n_4190),
.Y(n_4816)
);

AOI221x1_ASAP7_75t_L g4817 ( 
.A1(n_4355),
.A2(n_1670),
.B1(n_1672),
.B2(n_1669),
.C(n_1668),
.Y(n_4817)
);

NOR2xp33_ASAP7_75t_SL g4818 ( 
.A(n_4525),
.B(n_931),
.Y(n_4818)
);

OAI21x1_ASAP7_75t_L g4819 ( 
.A1(n_4383),
.A2(n_4559),
.B(n_4551),
.Y(n_4819)
);

AO31x2_ASAP7_75t_L g4820 ( 
.A1(n_4249),
.A2(n_1600),
.A3(n_1602),
.B(n_1599),
.Y(n_4820)
);

BUFx6f_ASAP7_75t_L g4821 ( 
.A(n_4400),
.Y(n_4821)
);

OAI21x1_ASAP7_75t_L g4822 ( 
.A1(n_4418),
.A2(n_2312),
.B(n_2308),
.Y(n_4822)
);

AND2x4_ASAP7_75t_L g4823 ( 
.A(n_4250),
.B(n_1542),
.Y(n_4823)
);

NAND2x1_ASAP7_75t_L g4824 ( 
.A(n_4545),
.B(n_2308),
.Y(n_4824)
);

AOI21xp5_ASAP7_75t_L g4825 ( 
.A1(n_4251),
.A2(n_2312),
.B(n_2308),
.Y(n_4825)
);

OAI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4259),
.A2(n_1672),
.B(n_1670),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4361),
.Y(n_4827)
);

AO31x2_ASAP7_75t_L g4828 ( 
.A1(n_4279),
.A2(n_1602),
.A3(n_1605),
.B(n_1600),
.Y(n_4828)
);

OAI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4295),
.A2(n_1677),
.B(n_1676),
.Y(n_4829)
);

INVxp67_ASAP7_75t_SL g4830 ( 
.A(n_4269),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4483),
.B(n_1215),
.Y(n_4831)
);

OAI21x1_ASAP7_75t_L g4832 ( 
.A1(n_4411),
.A2(n_2322),
.B(n_2312),
.Y(n_4832)
);

AO31x2_ASAP7_75t_L g4833 ( 
.A1(n_4503),
.A2(n_1611),
.A3(n_1612),
.B(n_1605),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4440),
.A2(n_4433),
.B(n_4471),
.Y(n_4834)
);

OAI21xp5_ASAP7_75t_L g4835 ( 
.A1(n_4295),
.A2(n_1677),
.B(n_1676),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4204),
.B(n_1683),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4239),
.B(n_1683),
.Y(n_4837)
);

BUFx3_ASAP7_75t_L g4838 ( 
.A(n_4497),
.Y(n_4838)
);

OAI21xp5_ASAP7_75t_L g4839 ( 
.A1(n_4211),
.A2(n_1691),
.B(n_1688),
.Y(n_4839)
);

OAI21x1_ASAP7_75t_L g4840 ( 
.A1(n_4495),
.A2(n_2327),
.B(n_2322),
.Y(n_4840)
);

INVx2_ASAP7_75t_L g4841 ( 
.A(n_4381),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_L g4842 ( 
.A(n_4247),
.B(n_1688),
.Y(n_4842)
);

OAI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4518),
.A2(n_1694),
.B(n_1691),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4334),
.B(n_1694),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4312),
.B(n_1543),
.Y(n_4845)
);

BUFx6f_ASAP7_75t_L g4846 ( 
.A(n_4454),
.Y(n_4846)
);

OAI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4485),
.A2(n_1612),
.B(n_1611),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_L g4848 ( 
.A(n_4183),
.B(n_1545),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4405),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4437),
.Y(n_4850)
);

OAI21x1_ASAP7_75t_L g4851 ( 
.A1(n_4495),
.A2(n_2327),
.B(n_2322),
.Y(n_4851)
);

OAI22xp5_ASAP7_75t_L g4852 ( 
.A1(n_4386),
.A2(n_1225),
.B1(n_1233),
.B2(n_1224),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4496),
.B(n_1234),
.Y(n_4853)
);

BUFx4f_ASAP7_75t_L g4854 ( 
.A(n_4308),
.Y(n_4854)
);

OAI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4527),
.A2(n_1619),
.B(n_1617),
.Y(n_4855)
);

AOI21xp5_ASAP7_75t_L g4856 ( 
.A1(n_4412),
.A2(n_2327),
.B(n_2322),
.Y(n_4856)
);

NOR2xp67_ASAP7_75t_SL g4857 ( 
.A(n_4549),
.B(n_1546),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4382),
.Y(n_4858)
);

OAI21x1_ASAP7_75t_L g4859 ( 
.A1(n_4438),
.A2(n_2334),
.B(n_2327),
.Y(n_4859)
);

AO21x2_ASAP7_75t_L g4860 ( 
.A1(n_4297),
.A2(n_1619),
.B(n_1617),
.Y(n_4860)
);

BUFx3_ASAP7_75t_L g4861 ( 
.A(n_4497),
.Y(n_4861)
);

AND2x2_ASAP7_75t_L g4862 ( 
.A(n_4334),
.B(n_1547),
.Y(n_4862)
);

INVx3_ASAP7_75t_SL g4863 ( 
.A(n_4169),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4323),
.Y(n_4864)
);

A2O1A1Ixp33_ASAP7_75t_L g4865 ( 
.A1(n_4550),
.A2(n_1245),
.B(n_1246),
.C(n_1243),
.Y(n_4865)
);

OAI22xp5_ASAP7_75t_L g4866 ( 
.A1(n_4386),
.A2(n_1249),
.B1(n_1550),
.B2(n_1549),
.Y(n_4866)
);

AOI21xp5_ASAP7_75t_L g4867 ( 
.A1(n_4412),
.A2(n_2337),
.B(n_2334),
.Y(n_4867)
);

BUFx6f_ASAP7_75t_L g4868 ( 
.A(n_4454),
.Y(n_4868)
);

OAI21x1_ASAP7_75t_L g4869 ( 
.A1(n_4446),
.A2(n_2337),
.B(n_2334),
.Y(n_4869)
);

AOI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4258),
.A2(n_2337),
.B(n_2334),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4533),
.B(n_4285),
.Y(n_4871)
);

OAI22x1_ASAP7_75t_L g4872 ( 
.A1(n_4434),
.A2(n_1557),
.B1(n_1559),
.B2(n_1551),
.Y(n_4872)
);

OAI21x1_ASAP7_75t_L g4873 ( 
.A1(n_4526),
.A2(n_2339),
.B(n_2337),
.Y(n_4873)
);

CKINVDCx12_ASAP7_75t_R g4874 ( 
.A(n_4200),
.Y(n_4874)
);

AOI21xp5_ASAP7_75t_L g4875 ( 
.A1(n_4232),
.A2(n_2360),
.B(n_2339),
.Y(n_4875)
);

INVx2_ASAP7_75t_L g4876 ( 
.A(n_4311),
.Y(n_4876)
);

BUFx2_ASAP7_75t_L g4877 ( 
.A(n_4426),
.Y(n_4877)
);

INVx3_ASAP7_75t_L g4878 ( 
.A(n_4509),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4358),
.A2(n_4294),
.B(n_4321),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4311),
.Y(n_4880)
);

AOI21xp5_ASAP7_75t_L g4881 ( 
.A1(n_4358),
.A2(n_2360),
.B(n_2339),
.Y(n_4881)
);

OAI21x1_ASAP7_75t_L g4882 ( 
.A1(n_4537),
.A2(n_2360),
.B(n_2339),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4306),
.Y(n_4883)
);

OAI21x1_ASAP7_75t_L g4884 ( 
.A1(n_4562),
.A2(n_2361),
.B(n_2360),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4207),
.B(n_1560),
.Y(n_4885)
);

AND2x2_ASAP7_75t_L g4886 ( 
.A(n_4357),
.B(n_1565),
.Y(n_4886)
);

BUFx3_ASAP7_75t_L g4887 ( 
.A(n_4169),
.Y(n_4887)
);

AOI21xp5_ASAP7_75t_L g4888 ( 
.A1(n_4290),
.A2(n_2374),
.B(n_2361),
.Y(n_4888)
);

OAI21x1_ASAP7_75t_L g4889 ( 
.A1(n_4552),
.A2(n_2374),
.B(n_2361),
.Y(n_4889)
);

OR2x6_ASAP7_75t_L g4890 ( 
.A(n_4333),
.B(n_4368),
.Y(n_4890)
);

BUFx10_ASAP7_75t_L g4891 ( 
.A(n_4222),
.Y(n_4891)
);

A2O1A1Ixp33_ASAP7_75t_L g4892 ( 
.A1(n_4350),
.A2(n_1567),
.B(n_1568),
.C(n_1566),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4307),
.A2(n_2374),
.B(n_2361),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4193),
.B(n_1569),
.Y(n_4894)
);

BUFx2_ASAP7_75t_L g4895 ( 
.A(n_4415),
.Y(n_4895)
);

NAND2x1p5_ASAP7_75t_L g4896 ( 
.A(n_4531),
.B(n_2374),
.Y(n_4896)
);

BUFx6f_ASAP7_75t_L g4897 ( 
.A(n_4454),
.Y(n_4897)
);

OAI21x1_ASAP7_75t_L g4898 ( 
.A1(n_4492),
.A2(n_2407),
.B(n_2396),
.Y(n_4898)
);

A2O1A1Ixp33_ASAP7_75t_L g4899 ( 
.A1(n_4345),
.A2(n_1572),
.B(n_1573),
.C(n_1570),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4221),
.Y(n_4900)
);

NAND2x1p5_ASAP7_75t_L g4901 ( 
.A(n_4275),
.B(n_2396),
.Y(n_4901)
);

CKINVDCx5p33_ASAP7_75t_R g4902 ( 
.A(n_4187),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4509),
.Y(n_4903)
);

INVx5_ASAP7_75t_L g4904 ( 
.A(n_4368),
.Y(n_4904)
);

BUFx6f_ASAP7_75t_L g4905 ( 
.A(n_4468),
.Y(n_4905)
);

AOI21xp5_ASAP7_75t_L g4906 ( 
.A1(n_4399),
.A2(n_4225),
.B(n_4419),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4460),
.B(n_1578),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4549),
.A2(n_2407),
.B(n_2396),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4499),
.B(n_1580),
.Y(n_4909)
);

AOI21x1_ASAP7_75t_L g4910 ( 
.A1(n_4511),
.A2(n_1622),
.B(n_1581),
.Y(n_4910)
);

OAI21x1_ASAP7_75t_L g4911 ( 
.A1(n_4520),
.A2(n_2407),
.B(n_2396),
.Y(n_4911)
);

AOI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4302),
.A2(n_4523),
.B(n_4512),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_4505),
.B(n_1622),
.Y(n_4913)
);

AOI221x1_ASAP7_75t_L g4914 ( 
.A1(n_4508),
.A2(n_1812),
.B1(n_1848),
.B2(n_1824),
.C(n_2040),
.Y(n_4914)
);

OAI22x1_ASAP7_75t_L g4915 ( 
.A1(n_4563),
.A2(n_984),
.B1(n_1050),
.B2(n_946),
.Y(n_4915)
);

BUFx6f_ASAP7_75t_SL g4916 ( 
.A(n_4174),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4510),
.B(n_946),
.Y(n_4917)
);

OAI21x1_ASAP7_75t_L g4918 ( 
.A1(n_4515),
.A2(n_2415),
.B(n_2407),
.Y(n_4918)
);

AOI22xp5_ASAP7_75t_L g4919 ( 
.A1(n_4389),
.A2(n_984),
.B1(n_1050),
.B2(n_946),
.Y(n_4919)
);

NOR2xp33_ASAP7_75t_L g4920 ( 
.A(n_4192),
.B(n_984),
.Y(n_4920)
);

BUFx6f_ASAP7_75t_L g4921 ( 
.A(n_4468),
.Y(n_4921)
);

OA21x2_ASAP7_75t_L g4922 ( 
.A1(n_4508),
.A2(n_1824),
.B(n_1812),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_SL g4923 ( 
.A(n_4320),
.B(n_984),
.Y(n_4923)
);

OAI21x1_ASAP7_75t_L g4924 ( 
.A1(n_4319),
.A2(n_2417),
.B(n_2415),
.Y(n_4924)
);

AO32x2_ASAP7_75t_L g4925 ( 
.A1(n_4546),
.A2(n_1082),
.A3(n_1192),
.B1(n_1050),
.B2(n_984),
.Y(n_4925)
);

OAI21x1_ASAP7_75t_L g4926 ( 
.A1(n_4502),
.A2(n_2417),
.B(n_2415),
.Y(n_4926)
);

AOI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4300),
.A2(n_1082),
.B1(n_1192),
.B2(n_1050),
.Y(n_4927)
);

OAI22xp5_ASAP7_75t_L g4928 ( 
.A1(n_4451),
.A2(n_4522),
.B1(n_4452),
.B2(n_4432),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4425),
.B(n_1050),
.Y(n_4929)
);

O2A1O1Ixp5_ASAP7_75t_L g4930 ( 
.A1(n_4248),
.A2(n_2415),
.B(n_2419),
.C(n_2417),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4546),
.B(n_3),
.Y(n_4931)
);

HB1xp67_ASAP7_75t_L g4932 ( 
.A(n_4368),
.Y(n_4932)
);

AOI21x1_ASAP7_75t_L g4933 ( 
.A1(n_4342),
.A2(n_1848),
.B(n_1945),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4439),
.B(n_1082),
.Y(n_4934)
);

AOI21x1_ASAP7_75t_L g4935 ( 
.A1(n_4443),
.A2(n_1970),
.B(n_1965),
.Y(n_4935)
);

CKINVDCx20_ASAP7_75t_R g4936 ( 
.A(n_4489),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_4513),
.A2(n_2419),
.B(n_2417),
.Y(n_4937)
);

INVx3_ASAP7_75t_L g4938 ( 
.A(n_4404),
.Y(n_4938)
);

AOI22xp5_ASAP7_75t_L g4939 ( 
.A1(n_4477),
.A2(n_1192),
.B1(n_1231),
.B2(n_1082),
.Y(n_4939)
);

OR2x2_ASAP7_75t_L g4940 ( 
.A(n_4337),
.B(n_4338),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4536),
.B(n_4),
.Y(n_4941)
);

AOI21xp33_ASAP7_75t_L g4942 ( 
.A1(n_4332),
.A2(n_4),
.B(n_5),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4414),
.B(n_5),
.Y(n_4943)
);

AOI211x1_ASAP7_75t_L g4944 ( 
.A1(n_4185),
.A2(n_1192),
.B(n_1231),
.C(n_1082),
.Y(n_4944)
);

AND3x4_ASAP7_75t_L g4945 ( 
.A(n_4174),
.B(n_4250),
.C(n_4198),
.Y(n_4945)
);

AO31x2_ASAP7_75t_L g4946 ( 
.A1(n_4514),
.A2(n_1970),
.A3(n_1971),
.B(n_1965),
.Y(n_4946)
);

INVx2_ASAP7_75t_SL g4947 ( 
.A(n_4424),
.Y(n_4947)
);

NOR2xp67_ASAP7_75t_L g4948 ( 
.A(n_4291),
.B(n_5),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_SL g4949 ( 
.A(n_4414),
.B(n_1192),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4441),
.B(n_1231),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4444),
.B(n_6),
.Y(n_4951)
);

AOI221x1_ASAP7_75t_L g4952 ( 
.A1(n_4402),
.A2(n_2040),
.B1(n_2053),
.B2(n_2050),
.C(n_2048),
.Y(n_4952)
);

OAI21x1_ASAP7_75t_L g4953 ( 
.A1(n_4166),
.A2(n_2448),
.B(n_2419),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4444),
.A2(n_2448),
.B(n_2419),
.Y(n_4954)
);

OAI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4456),
.A2(n_2450),
.B(n_2448),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4524),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4166),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_SL g4958 ( 
.A(n_4230),
.B(n_4532),
.Y(n_4958)
);

AO21x1_ASAP7_75t_L g4959 ( 
.A1(n_4352),
.A2(n_1231),
.B(n_6),
.Y(n_4959)
);

OAI21x1_ASAP7_75t_L g4960 ( 
.A1(n_4205),
.A2(n_4473),
.B(n_2450),
.Y(n_4960)
);

BUFx6f_ASAP7_75t_L g4961 ( 
.A(n_4468),
.Y(n_4961)
);

OAI21x1_ASAP7_75t_L g4962 ( 
.A1(n_4205),
.A2(n_2450),
.B(n_2448),
.Y(n_4962)
);

OAI22xp5_ASAP7_75t_L g4963 ( 
.A1(n_4340),
.A2(n_1231),
.B1(n_10),
.B2(n_7),
.Y(n_4963)
);

NOR2xp33_ASAP7_75t_L g4964 ( 
.A(n_4375),
.B(n_90),
.Y(n_4964)
);

NAND2xp5_ASAP7_75t_L g4965 ( 
.A(n_4488),
.B(n_4344),
.Y(n_4965)
);

OAI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4348),
.A2(n_2455),
.B(n_2450),
.Y(n_4966)
);

OAI21x1_ASAP7_75t_L g4967 ( 
.A1(n_4473),
.A2(n_2455),
.B(n_2066),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4365),
.Y(n_4968)
);

AO31x2_ASAP7_75t_L g4969 ( 
.A1(n_4404),
.A2(n_1980),
.A3(n_2006),
.B(n_1971),
.Y(n_4969)
);

OAI22xp5_ASAP7_75t_L g4970 ( 
.A1(n_4369),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_SL g4971 ( 
.A(n_4532),
.B(n_2040),
.Y(n_4971)
);

A2O1A1Ixp33_ASAP7_75t_L g4972 ( 
.A1(n_4378),
.A2(n_2455),
.B(n_1297),
.C(n_1300),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_SL g4973 ( 
.A(n_4553),
.B(n_4455),
.Y(n_4973)
);

OR2x6_ASAP7_75t_L g4974 ( 
.A(n_4545),
.B(n_1797),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_SL g4975 ( 
.A(n_4553),
.B(n_2040),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4455),
.B(n_7),
.Y(n_4976)
);

AOI21xp5_ASAP7_75t_L g4977 ( 
.A1(n_4459),
.A2(n_2455),
.B(n_2244),
.Y(n_4977)
);

OAI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4370),
.A2(n_2006),
.B(n_1980),
.Y(n_4978)
);

OAI22xp5_ASAP7_75t_L g4979 ( 
.A1(n_4374),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_4979)
);

CKINVDCx5p33_ASAP7_75t_R g4980 ( 
.A(n_4424),
.Y(n_4980)
);

OAI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4376),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_4981)
);

OAI21x1_ASAP7_75t_L g4982 ( 
.A1(n_4397),
.A2(n_2066),
.B(n_2060),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4459),
.B(n_11),
.Y(n_4983)
);

HB1xp67_ASAP7_75t_L g4984 ( 
.A(n_4343),
.Y(n_4984)
);

NAND2x1_ASAP7_75t_L g4985 ( 
.A(n_4553),
.B(n_2060),
.Y(n_4985)
);

BUFx6f_ASAP7_75t_L g4986 ( 
.A(n_4602),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4830),
.B(n_4814),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4577),
.Y(n_4988)
);

OAI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4818),
.A2(n_4777),
.B1(n_4778),
.B2(n_4939),
.Y(n_4989)
);

BUFx2_ASAP7_75t_L g4990 ( 
.A(n_4788),
.Y(n_4990)
);

NAND3xp33_ASAP7_75t_L g4991 ( 
.A(n_4624),
.B(n_4481),
.C(n_4366),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4624),
.A2(n_4416),
.B(n_4343),
.Y(n_4992)
);

OAI22xp5_ASAP7_75t_L g4993 ( 
.A1(n_4786),
.A2(n_4416),
.B1(n_4343),
.B2(n_4445),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4654),
.A2(n_4416),
.B(n_4528),
.Y(n_4994)
);

BUFx6f_ASAP7_75t_L g4995 ( 
.A(n_4602),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4684),
.B(n_4421),
.Y(n_4996)
);

OAI21x1_ASAP7_75t_L g4997 ( 
.A1(n_4809),
.A2(n_2025),
.B(n_2023),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4600),
.Y(n_4998)
);

CKINVDCx8_ASAP7_75t_R g4999 ( 
.A(n_4598),
.Y(n_4999)
);

INVx2_ASAP7_75t_SL g5000 ( 
.A(n_4602),
.Y(n_5000)
);

AOI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_4654),
.A2(n_4416),
.B(n_4465),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4605),
.Y(n_5002)
);

O2A1O1Ixp33_ASAP7_75t_L g5003 ( 
.A1(n_4736),
.A2(n_4470),
.B(n_4465),
.C(n_1297),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4650),
.Y(n_5004)
);

INVx2_ASAP7_75t_L g5005 ( 
.A(n_4665),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4680),
.Y(n_5006)
);

INVx3_ASAP7_75t_SL g5007 ( 
.A(n_4681),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4695),
.Y(n_5008)
);

AOI21xp33_ASAP7_75t_L g5009 ( 
.A1(n_4575),
.A2(n_4638),
.B(n_4631),
.Y(n_5009)
);

BUFx10_ASAP7_75t_L g5010 ( 
.A(n_4801),
.Y(n_5010)
);

INVxp67_ASAP7_75t_L g5011 ( 
.A(n_4733),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_4613),
.B(n_4445),
.Y(n_5012)
);

BUFx2_ASAP7_75t_L g5013 ( 
.A(n_4752),
.Y(n_5013)
);

AND2x2_ASAP7_75t_SL g5014 ( 
.A(n_4818),
.B(n_4424),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4673),
.B(n_90),
.Y(n_5015)
);

HB1xp67_ASAP7_75t_L g5016 ( 
.A(n_4729),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4763),
.Y(n_5017)
);

INVx1_ASAP7_75t_SL g5018 ( 
.A(n_4816),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4673),
.B(n_92),
.Y(n_5019)
);

CKINVDCx11_ASAP7_75t_R g5020 ( 
.A(n_4661),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4585),
.B(n_12),
.Y(n_5021)
);

OAI21xp5_ASAP7_75t_L g5022 ( 
.A1(n_4748),
.A2(n_2025),
.B(n_2023),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4772),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_4776),
.Y(n_5024)
);

INVx5_ASAP7_75t_L g5025 ( 
.A(n_4974),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4708),
.Y(n_5026)
);

BUFx6f_ASAP7_75t_L g5027 ( 
.A(n_4644),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4793),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4813),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_SL g5030 ( 
.A(n_4575),
.B(n_2040),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4879),
.A2(n_4952),
.B(n_4580),
.Y(n_5031)
);

AND2x4_ASAP7_75t_L g5032 ( 
.A(n_4629),
.B(n_2048),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4850),
.Y(n_5033)
);

AOI22xp33_ASAP7_75t_L g5034 ( 
.A1(n_4748),
.A2(n_2050),
.B1(n_2053),
.B2(n_2048),
.Y(n_5034)
);

BUFx10_ASAP7_75t_L g5035 ( 
.A(n_4902),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_4686),
.Y(n_5036)
);

OAI22xp5_ASAP7_75t_L g5037 ( 
.A1(n_4617),
.A2(n_4931),
.B1(n_4725),
.B2(n_4963),
.Y(n_5037)
);

CKINVDCx6p67_ASAP7_75t_R g5038 ( 
.A(n_4687),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4580),
.A2(n_2244),
.B(n_2231),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_4585),
.B(n_4956),
.Y(n_5040)
);

NOR2xp67_ASAP7_75t_SL g5041 ( 
.A(n_4812),
.B(n_2048),
.Y(n_5041)
);

BUFx12f_ASAP7_75t_L g5042 ( 
.A(n_4891),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4729),
.Y(n_5043)
);

AOI21xp5_ASAP7_75t_L g5044 ( 
.A1(n_4632),
.A2(n_2244),
.B(n_2231),
.Y(n_5044)
);

A2O1A1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4964),
.A2(n_93),
.B(n_94),
.C(n_92),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4629),
.B(n_4877),
.Y(n_5046)
);

AOI21xp5_ASAP7_75t_L g5047 ( 
.A1(n_4632),
.A2(n_2244),
.B(n_2231),
.Y(n_5047)
);

INVx2_ASAP7_75t_L g5048 ( 
.A(n_4572),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4900),
.B(n_13),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4883),
.B(n_13),
.Y(n_5050)
);

INVx3_ASAP7_75t_L g5051 ( 
.A(n_4887),
.Y(n_5051)
);

NOR2xp33_ASAP7_75t_L g5052 ( 
.A(n_4940),
.B(n_95),
.Y(n_5052)
);

OR2x6_ASAP7_75t_L g5053 ( 
.A(n_4756),
.B(n_2048),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_4895),
.B(n_96),
.Y(n_5054)
);

NAND3xp33_ASAP7_75t_L g5055 ( 
.A(n_4596),
.B(n_2053),
.C(n_2050),
.Y(n_5055)
);

NOR2xp33_ASAP7_75t_L g5056 ( 
.A(n_4626),
.B(n_96),
.Y(n_5056)
);

A2O1A1Ixp33_ASAP7_75t_SL g5057 ( 
.A1(n_4757),
.A2(n_2029),
.B(n_1713),
.C(n_1703),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4628),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4871),
.B(n_97),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4816),
.B(n_97),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4631),
.B(n_14),
.Y(n_5061)
);

NOR2x1_ASAP7_75t_SL g5062 ( 
.A(n_4635),
.B(n_4756),
.Y(n_5062)
);

AOI21xp33_ASAP7_75t_L g5063 ( 
.A1(n_4638),
.A2(n_14),
.B(n_15),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4639),
.Y(n_5064)
);

NAND2x1p5_ASAP7_75t_L g5065 ( 
.A(n_4647),
.B(n_1797),
.Y(n_5065)
);

INVx3_ASAP7_75t_L g5066 ( 
.A(n_4916),
.Y(n_5066)
);

OAI22xp5_ASAP7_75t_L g5067 ( 
.A1(n_4617),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_5067)
);

OR2x6_ASAP7_75t_L g5068 ( 
.A(n_4756),
.B(n_4635),
.Y(n_5068)
);

AOI21xp5_ASAP7_75t_L g5069 ( 
.A1(n_4632),
.A2(n_2244),
.B(n_2231),
.Y(n_5069)
);

INVx3_ASAP7_75t_L g5070 ( 
.A(n_4916),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4651),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4694),
.Y(n_5072)
);

NOR2x1_ASAP7_75t_SL g5073 ( 
.A(n_4635),
.B(n_4719),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4761),
.Y(n_5074)
);

INVx3_ASAP7_75t_L g5075 ( 
.A(n_4644),
.Y(n_5075)
);

INVx2_ASAP7_75t_L g5076 ( 
.A(n_4804),
.Y(n_5076)
);

AND2x4_ASAP7_75t_L g5077 ( 
.A(n_4719),
.B(n_2050),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4567),
.B(n_15),
.Y(n_5078)
);

INVx2_ASAP7_75t_L g5079 ( 
.A(n_4827),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4841),
.Y(n_5080)
);

OA21x2_ASAP7_75t_L g5081 ( 
.A1(n_4982),
.A2(n_2029),
.B(n_1300),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4849),
.Y(n_5082)
);

O2A1O1Ixp5_ASAP7_75t_L g5083 ( 
.A1(n_4959),
.A2(n_1301),
.B(n_1302),
.C(n_1296),
.Y(n_5083)
);

BUFx6f_ASAP7_75t_L g5084 ( 
.A(n_4644),
.Y(n_5084)
);

BUFx12f_ASAP7_75t_L g5085 ( 
.A(n_4891),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4567),
.B(n_16),
.Y(n_5086)
);

O2A1O1Ixp33_ASAP7_75t_L g5087 ( 
.A1(n_4963),
.A2(n_1301),
.B(n_1302),
.C(n_1296),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_4903),
.Y(n_5088)
);

INVx2_ASAP7_75t_SL g5089 ( 
.A(n_4663),
.Y(n_5089)
);

INVx1_ASAP7_75t_SL g5090 ( 
.A(n_4612),
.Y(n_5090)
);

INVx2_ASAP7_75t_L g5091 ( 
.A(n_4878),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_4876),
.B(n_98),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_4878),
.Y(n_5093)
);

AND2x4_ASAP7_75t_L g5094 ( 
.A(n_4719),
.B(n_2050),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_SL g5095 ( 
.A(n_4928),
.B(n_2053),
.Y(n_5095)
);

INVxp67_ASAP7_75t_L g5096 ( 
.A(n_4968),
.Y(n_5096)
);

AND2x4_ASAP7_75t_L g5097 ( 
.A(n_4890),
.B(n_2053),
.Y(n_5097)
);

AOI21xp33_ASAP7_75t_L g5098 ( 
.A1(n_4716),
.A2(n_4839),
.B(n_4599),
.Y(n_5098)
);

AOI22xp33_ASAP7_75t_L g5099 ( 
.A1(n_4633),
.A2(n_1921),
.B1(n_1929),
.B2(n_1914),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4858),
.Y(n_5100)
);

OAI22xp5_ASAP7_75t_L g5101 ( 
.A1(n_4931),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_5101)
);

INVxp67_ASAP7_75t_SL g5102 ( 
.A(n_4783),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4690),
.B(n_17),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_4864),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_4880),
.Y(n_5105)
);

A2O1A1Ixp33_ASAP7_75t_L g5106 ( 
.A1(n_4777),
.A2(n_104),
.B(n_105),
.C(n_103),
.Y(n_5106)
);

O2A1O1Ixp5_ASAP7_75t_L g5107 ( 
.A1(n_4942),
.A2(n_1308),
.B(n_1309),
.C(n_1307),
.Y(n_5107)
);

AOI222xp33_ASAP7_75t_L g5108 ( 
.A1(n_4970),
.A2(n_45),
.B1(n_26),
.B2(n_53),
.C1(n_35),
.C2(n_18),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4932),
.Y(n_5109)
);

INVxp67_ASAP7_75t_SL g5110 ( 
.A(n_4783),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_4568),
.B(n_103),
.Y(n_5111)
);

BUFx6f_ASAP7_75t_L g5112 ( 
.A(n_4663),
.Y(n_5112)
);

NOR2xp67_ASAP7_75t_L g5113 ( 
.A(n_4594),
.B(n_18),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4829),
.A2(n_2244),
.B(n_2231),
.Y(n_5114)
);

AOI22xp5_ASAP7_75t_L g5115 ( 
.A1(n_4778),
.A2(n_1308),
.B1(n_1309),
.B2(n_1307),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4829),
.A2(n_2287),
.B(n_2231),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4690),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4690),
.Y(n_5118)
);

AND2x2_ASAP7_75t_SL g5119 ( 
.A(n_4781),
.B(n_1914),
.Y(n_5119)
);

AND2x2_ASAP7_75t_L g5120 ( 
.A(n_4588),
.B(n_105),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_4641),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4641),
.Y(n_5122)
);

AND2x2_ASAP7_75t_SL g5123 ( 
.A(n_4606),
.B(n_1914),
.Y(n_5123)
);

NOR2x1_ASAP7_75t_SL g5124 ( 
.A(n_4647),
.B(n_1799),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_4643),
.Y(n_5125)
);

HB1xp67_ASAP7_75t_L g5126 ( 
.A(n_4583),
.Y(n_5126)
);

BUFx6f_ASAP7_75t_L g5127 ( 
.A(n_4663),
.Y(n_5127)
);

OR2x6_ASAP7_75t_L g5128 ( 
.A(n_4890),
.B(n_4912),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_4957),
.Y(n_5129)
);

A2O1A1Ixp33_ASAP7_75t_L g5130 ( 
.A1(n_4919),
.A2(n_107),
.B(n_108),
.C(n_106),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4835),
.A2(n_4834),
.B(n_4720),
.Y(n_5131)
);

NOR2xp33_ASAP7_75t_L g5132 ( 
.A(n_4874),
.B(n_106),
.Y(n_5132)
);

INVx5_ASAP7_75t_L g5133 ( 
.A(n_4974),
.Y(n_5133)
);

CKINVDCx20_ASAP7_75t_R g5134 ( 
.A(n_4936),
.Y(n_5134)
);

AOI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_4835),
.A2(n_2289),
.B(n_2287),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4844),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_4643),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_4595),
.B(n_19),
.Y(n_5138)
);

OAI22xp33_ASAP7_75t_L g5139 ( 
.A1(n_4927),
.A2(n_4599),
.B1(n_4979),
.B2(n_4970),
.Y(n_5139)
);

NOR2xp33_ASAP7_75t_L g5140 ( 
.A(n_4807),
.B(n_108),
.Y(n_5140)
);

BUFx6f_ASAP7_75t_L g5141 ( 
.A(n_4606),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4604),
.B(n_19),
.Y(n_5142)
);

O2A1O1Ixp33_ASAP7_75t_L g5143 ( 
.A1(n_4715),
.A2(n_1311),
.B(n_1313),
.C(n_1310),
.Y(n_5143)
);

AOI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_4647),
.A2(n_2289),
.B(n_2287),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4643),
.Y(n_5145)
);

BUFx10_ASAP7_75t_L g5146 ( 
.A(n_4702),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_4645),
.B(n_19),
.Y(n_5147)
);

INVx5_ASAP7_75t_L g5148 ( 
.A(n_4974),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_4616),
.Y(n_5149)
);

AOI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_4647),
.A2(n_2289),
.B(n_2287),
.Y(n_5150)
);

AND2x4_ASAP7_75t_L g5151 ( 
.A(n_4890),
.B(n_1914),
.Y(n_5151)
);

INVx3_ASAP7_75t_L g5152 ( 
.A(n_4616),
.Y(n_5152)
);

NOR2xp33_ASAP7_75t_SL g5153 ( 
.A(n_4854),
.B(n_1799),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_4762),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4723),
.Y(n_5155)
);

BUFx2_ASAP7_75t_L g5156 ( 
.A(n_4863),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4820),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_4645),
.B(n_20),
.Y(n_5158)
);

CKINVDCx5p33_ASAP7_75t_R g5159 ( 
.A(n_4780),
.Y(n_5159)
);

OAI21x1_ASAP7_75t_SL g5160 ( 
.A1(n_4601),
.A2(n_20),
.B(n_21),
.Y(n_5160)
);

INVx3_ASAP7_75t_L g5161 ( 
.A(n_4723),
.Y(n_5161)
);

BUFx6f_ASAP7_75t_L g5162 ( 
.A(n_4723),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4820),
.Y(n_5163)
);

OAI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4697),
.A2(n_1311),
.B(n_1310),
.Y(n_5164)
);

AOI22xp33_ASAP7_75t_L g5165 ( 
.A1(n_4942),
.A2(n_1921),
.B1(n_1929),
.B2(n_1914),
.Y(n_5165)
);

INVx2_ASAP7_75t_SL g5166 ( 
.A(n_4735),
.Y(n_5166)
);

INVx2_ASAP7_75t_SL g5167 ( 
.A(n_4670),
.Y(n_5167)
);

NAND2x1p5_ASAP7_75t_L g5168 ( 
.A(n_4720),
.B(n_1799),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_4740),
.B(n_109),
.Y(n_5169)
);

AND2x4_ASAP7_75t_L g5170 ( 
.A(n_4734),
.B(n_1921),
.Y(n_5170)
);

INVx1_ASAP7_75t_SL g5171 ( 
.A(n_4742),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4820),
.Y(n_5172)
);

NOR2xp33_ASAP7_75t_SL g5173 ( 
.A(n_4854),
.B(n_1799),
.Y(n_5173)
);

INVx5_ASAP7_75t_L g5174 ( 
.A(n_4810),
.Y(n_5174)
);

INVx2_ASAP7_75t_L g5175 ( 
.A(n_4770),
.Y(n_5175)
);

AND2x2_ASAP7_75t_L g5176 ( 
.A(n_4862),
.B(n_109),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4720),
.A2(n_4625),
.B(n_4656),
.Y(n_5177)
);

BUFx6f_ASAP7_75t_L g5178 ( 
.A(n_4770),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4770),
.Y(n_5179)
);

BUFx2_ASAP7_75t_L g5180 ( 
.A(n_4657),
.Y(n_5180)
);

NAND2x1p5_ASAP7_75t_L g5181 ( 
.A(n_4720),
.B(n_1799),
.Y(n_5181)
);

OR2x6_ASAP7_75t_L g5182 ( 
.A(n_4579),
.B(n_1921),
.Y(n_5182)
);

BUFx2_ASAP7_75t_L g5183 ( 
.A(n_4657),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_SL g5184 ( 
.A(n_4928),
.B(n_1921),
.Y(n_5184)
);

OAI22xp5_ASAP7_75t_SL g5185 ( 
.A1(n_4945),
.A2(n_4944),
.B1(n_4915),
.B2(n_4981),
.Y(n_5185)
);

BUFx2_ASAP7_75t_L g5186 ( 
.A(n_4666),
.Y(n_5186)
);

INVx3_ASAP7_75t_L g5187 ( 
.A(n_4821),
.Y(n_5187)
);

AND2x4_ASAP7_75t_L g5188 ( 
.A(n_4734),
.B(n_1929),
.Y(n_5188)
);

NOR2xp33_ASAP7_75t_L g5189 ( 
.A(n_4658),
.B(n_110),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_4645),
.B(n_20),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4744),
.B(n_21),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_4821),
.Y(n_5192)
);

AOI21xp5_ASAP7_75t_L g5193 ( 
.A1(n_4625),
.A2(n_2289),
.B(n_2287),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_L g5194 ( 
.A(n_4744),
.B(n_4745),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4821),
.Y(n_5195)
);

BUFx3_ASAP7_75t_L g5196 ( 
.A(n_4590),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_4745),
.B(n_21),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_4721),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_4751),
.B(n_22),
.Y(n_5199)
);

INVx2_ASAP7_75t_L g5200 ( 
.A(n_4846),
.Y(n_5200)
);

INVx3_ASAP7_75t_SL g5201 ( 
.A(n_4980),
.Y(n_5201)
);

AOI22xp33_ASAP7_75t_L g5202 ( 
.A1(n_4715),
.A2(n_1941),
.B1(n_1947),
.B2(n_1929),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_4846),
.Y(n_5203)
);

AOI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_4656),
.A2(n_2289),
.B(n_2287),
.Y(n_5204)
);

OAI22xp5_ASAP7_75t_L g5205 ( 
.A1(n_4979),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4721),
.Y(n_5206)
);

BUFx6f_ASAP7_75t_L g5207 ( 
.A(n_4846),
.Y(n_5207)
);

OAI21xp33_ASAP7_75t_L g5208 ( 
.A1(n_4981),
.A2(n_23),
.B(n_24),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4732),
.Y(n_5209)
);

INVx2_ASAP7_75t_L g5210 ( 
.A(n_4868),
.Y(n_5210)
);

BUFx4f_ASAP7_75t_SL g5211 ( 
.A(n_4838),
.Y(n_5211)
);

AOI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4589),
.A2(n_2291),
.B(n_2289),
.Y(n_5212)
);

AND2x2_ASAP7_75t_L g5213 ( 
.A(n_4771),
.B(n_4805),
.Y(n_5213)
);

INVx4_ASAP7_75t_L g5214 ( 
.A(n_4810),
.Y(n_5214)
);

AND2x4_ASAP7_75t_L g5215 ( 
.A(n_4734),
.B(n_1929),
.Y(n_5215)
);

AND2x4_ASAP7_75t_L g5216 ( 
.A(n_4734),
.B(n_1941),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_4868),
.Y(n_5217)
);

BUFx12f_ASAP7_75t_L g5218 ( 
.A(n_4714),
.Y(n_5218)
);

OR2x6_ASAP7_75t_SL g5219 ( 
.A(n_4584),
.B(n_1313),
.Y(n_5219)
);

BUFx6f_ASAP7_75t_L g5220 ( 
.A(n_4868),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_4897),
.Y(n_5221)
);

BUFx3_ASAP7_75t_L g5222 ( 
.A(n_4785),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_4768),
.B(n_112),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_4897),
.Y(n_5224)
);

BUFx3_ASAP7_75t_L g5225 ( 
.A(n_4861),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4732),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_L g5227 ( 
.A(n_4662),
.B(n_114),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_4751),
.B(n_25),
.Y(n_5228)
);

AND2x4_ASAP7_75t_L g5229 ( 
.A(n_4800),
.B(n_1941),
.Y(n_5229)
);

OR2x6_ASAP7_75t_L g5230 ( 
.A(n_4958),
.B(n_1941),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4755),
.B(n_25),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4897),
.Y(n_5232)
);

BUFx2_ASAP7_75t_L g5233 ( 
.A(n_4666),
.Y(n_5233)
);

OAI22xp5_ASAP7_75t_L g5234 ( 
.A1(n_4573),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4707),
.Y(n_5235)
);

OAI21xp5_ASAP7_75t_L g5236 ( 
.A1(n_4706),
.A2(n_1320),
.B(n_1316),
.Y(n_5236)
);

INVx5_ASAP7_75t_L g5237 ( 
.A(n_4905),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_4907),
.B(n_115),
.Y(n_5238)
);

BUFx12f_ASAP7_75t_L g5239 ( 
.A(n_4823),
.Y(n_5239)
);

O2A1O1Ixp33_ASAP7_75t_L g5240 ( 
.A1(n_4609),
.A2(n_4622),
.B(n_4630),
.C(n_4603),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4707),
.Y(n_5241)
);

A2O1A1Ixp33_ASAP7_75t_L g5242 ( 
.A1(n_4965),
.A2(n_117),
.B(n_118),
.C(n_116),
.Y(n_5242)
);

AOI21xp5_ASAP7_75t_L g5243 ( 
.A1(n_4589),
.A2(n_2292),
.B(n_2291),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_4905),
.Y(n_5244)
);

OAI22xp5_ASAP7_75t_L g5245 ( 
.A1(n_4584),
.A2(n_4696),
.B1(n_4948),
.B2(n_4693),
.Y(n_5245)
);

INVx5_ASAP7_75t_L g5246 ( 
.A(n_4905),
.Y(n_5246)
);

AOI21xp5_ASAP7_75t_L g5247 ( 
.A1(n_4698),
.A2(n_2292),
.B(n_2291),
.Y(n_5247)
);

BUFx12f_ASAP7_75t_L g5248 ( 
.A(n_4823),
.Y(n_5248)
);

O2A1O1Ixp5_ASAP7_75t_SL g5249 ( 
.A1(n_4696),
.A2(n_1320),
.B(n_1316),
.C(n_1713),
.Y(n_5249)
);

AO31x2_ASAP7_75t_L g5250 ( 
.A1(n_4914),
.A2(n_2228),
.A3(n_2354),
.B(n_2206),
.Y(n_5250)
);

INVxp67_ASAP7_75t_SL g5251 ( 
.A(n_4901),
.Y(n_5251)
);

NOR2xp33_ASAP7_75t_L g5252 ( 
.A(n_4685),
.B(n_4886),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_4707),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_4636),
.B(n_117),
.Y(n_5254)
);

AOI21xp5_ASAP7_75t_L g5255 ( 
.A1(n_4698),
.A2(n_2292),
.B(n_2291),
.Y(n_5255)
);

OAI22xp5_ASAP7_75t_L g5256 ( 
.A1(n_4865),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_4921),
.Y(n_5257)
);

AOI21xp5_ASAP7_75t_L g5258 ( 
.A1(n_4637),
.A2(n_2292),
.B(n_2291),
.Y(n_5258)
);

AOI21xp5_ASAP7_75t_L g5259 ( 
.A1(n_4637),
.A2(n_2292),
.B(n_2291),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_4741),
.Y(n_5260)
);

O2A1O1Ixp33_ASAP7_75t_L g5261 ( 
.A1(n_4923),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_4640),
.B(n_118),
.Y(n_5262)
);

BUFx3_ASAP7_75t_L g5263 ( 
.A(n_4921),
.Y(n_5263)
);

INVx3_ASAP7_75t_L g5264 ( 
.A(n_4921),
.Y(n_5264)
);

AOI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_4906),
.A2(n_2300),
.B(n_2292),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_4961),
.Y(n_5266)
);

NAND2x1p5_ASAP7_75t_L g5267 ( 
.A(n_4800),
.B(n_1941),
.Y(n_5267)
);

AOI21xp5_ASAP7_75t_L g5268 ( 
.A1(n_4930),
.A2(n_2303),
.B(n_2300),
.Y(n_5268)
);

AND2x4_ASAP7_75t_L g5269 ( 
.A(n_4800),
.B(n_1947),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_4961),
.Y(n_5270)
);

BUFx3_ASAP7_75t_L g5271 ( 
.A(n_4961),
.Y(n_5271)
);

CKINVDCx11_ASAP7_75t_R g5272 ( 
.A(n_4737),
.Y(n_5272)
);

INVx1_ASAP7_75t_SL g5273 ( 
.A(n_4984),
.Y(n_5273)
);

BUFx3_ASAP7_75t_L g5274 ( 
.A(n_4938),
.Y(n_5274)
);

AND2x2_ASAP7_75t_L g5275 ( 
.A(n_4718),
.B(n_119),
.Y(n_5275)
);

AOI21xp5_ASAP7_75t_L g5276 ( 
.A1(n_4839),
.A2(n_2303),
.B(n_2300),
.Y(n_5276)
);

AOI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_4706),
.A2(n_4737),
.B1(n_4570),
.B2(n_4758),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_4955),
.A2(n_2303),
.B(n_2300),
.Y(n_5278)
);

AND2x4_ASAP7_75t_L g5279 ( 
.A(n_4800),
.B(n_1947),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_SL g5280 ( 
.A(n_4640),
.B(n_1947),
.Y(n_5280)
);

AOI22xp5_ASAP7_75t_L g5281 ( 
.A1(n_4806),
.A2(n_1948),
.B1(n_1959),
.B2(n_1947),
.Y(n_5281)
);

INVx3_ASAP7_75t_L g5282 ( 
.A(n_4938),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_L g5283 ( 
.A1(n_4955),
.A2(n_2303),
.B(n_2300),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_4966),
.A2(n_2303),
.B(n_2300),
.Y(n_5284)
);

AOI21xp5_ASAP7_75t_L g5285 ( 
.A1(n_4966),
.A2(n_4731),
.B(n_4797),
.Y(n_5285)
);

AOI22xp33_ASAP7_75t_L g5286 ( 
.A1(n_4614),
.A2(n_1948),
.B1(n_1963),
.B2(n_1959),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_4741),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4797),
.A2(n_2313),
.B(n_2303),
.Y(n_5288)
);

INVxp67_ASAP7_75t_SL g5289 ( 
.A(n_4901),
.Y(n_5289)
);

BUFx6f_ASAP7_75t_L g5290 ( 
.A(n_4947),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_4741),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_4747),
.B(n_4619),
.Y(n_5292)
);

O2A1O1Ixp33_ASAP7_75t_L g5293 ( 
.A1(n_4726),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_5293)
);

AND2x2_ASAP7_75t_L g5294 ( 
.A(n_4943),
.B(n_119),
.Y(n_5294)
);

BUFx6f_ASAP7_75t_L g5295 ( 
.A(n_4824),
.Y(n_5295)
);

INVx2_ASAP7_75t_L g5296 ( 
.A(n_4946),
.Y(n_5296)
);

CKINVDCx20_ASAP7_75t_R g5297 ( 
.A(n_4774),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_4593),
.B(n_121),
.Y(n_5298)
);

OA21x2_ASAP7_75t_L g5299 ( 
.A1(n_4592),
.A2(n_42),
.B(n_31),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4975),
.A2(n_2313),
.B(n_2320),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4946),
.Y(n_5301)
);

BUFx2_ASAP7_75t_L g5302 ( 
.A(n_4904),
.Y(n_5302)
);

INVx2_ASAP7_75t_SL g5303 ( 
.A(n_4941),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4946),
.Y(n_5304)
);

AND2x4_ASAP7_75t_L g5305 ( 
.A(n_4904),
.B(n_4973),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4701),
.A2(n_2313),
.B(n_2320),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_L g5307 ( 
.A1(n_4701),
.A2(n_2313),
.B(n_2320),
.Y(n_5307)
);

NOR2xp33_ASAP7_75t_L g5308 ( 
.A(n_4782),
.B(n_122),
.Y(n_5308)
);

BUFx6f_ASAP7_75t_L g5309 ( 
.A(n_4943),
.Y(n_5309)
);

AOI22xp33_ASAP7_75t_L g5310 ( 
.A1(n_4739),
.A2(n_4653),
.B1(n_4949),
.B2(n_4671),
.Y(n_5310)
);

NAND2x2_ASAP7_75t_L g5311 ( 
.A(n_4929),
.B(n_4934),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_4951),
.Y(n_5312)
);

INVx3_ASAP7_75t_L g5313 ( 
.A(n_4904),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_4755),
.B(n_33),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_4746),
.B(n_33),
.Y(n_5315)
);

AOI221xp5_ASAP7_75t_L g5316 ( 
.A1(n_4852),
.A2(n_1963),
.B1(n_1964),
.B2(n_1959),
.C(n_1948),
.Y(n_5316)
);

BUFx2_ASAP7_75t_SL g5317 ( 
.A(n_4904),
.Y(n_5317)
);

AOI22xp33_ASAP7_75t_L g5318 ( 
.A1(n_4569),
.A2(n_1948),
.B1(n_1963),
.B2(n_1959),
.Y(n_5318)
);

NAND2x1p5_ASAP7_75t_L g5319 ( 
.A(n_4960),
.B(n_1948),
.Y(n_5319)
);

OAI22xp5_ASAP7_75t_L g5320 ( 
.A1(n_4675),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_5320)
);

CKINVDCx20_ASAP7_75t_R g5321 ( 
.A(n_4623),
.Y(n_5321)
);

BUFx6f_ASAP7_75t_L g5322 ( 
.A(n_4951),
.Y(n_5322)
);

BUFx3_ASAP7_75t_L g5323 ( 
.A(n_4941),
.Y(n_5323)
);

INVx8_ASAP7_75t_L g5324 ( 
.A(n_4571),
.Y(n_5324)
);

CKINVDCx5p33_ASAP7_75t_R g5325 ( 
.A(n_4920),
.Y(n_5325)
);

INVx2_ASAP7_75t_L g5326 ( 
.A(n_4976),
.Y(n_5326)
);

AND2x2_ASAP7_75t_L g5327 ( 
.A(n_4976),
.B(n_122),
.Y(n_5327)
);

AOI21xp5_ASAP7_75t_L g5328 ( 
.A1(n_4798),
.A2(n_2313),
.B(n_2320),
.Y(n_5328)
);

AOI21xp5_ASAP7_75t_L g5329 ( 
.A1(n_4798),
.A2(n_2313),
.B(n_2320),
.Y(n_5329)
);

AOI21xp5_ASAP7_75t_L g5330 ( 
.A1(n_4796),
.A2(n_2321),
.B(n_2320),
.Y(n_5330)
);

BUFx2_ASAP7_75t_L g5331 ( 
.A(n_4983),
.Y(n_5331)
);

CKINVDCx8_ASAP7_75t_R g5332 ( 
.A(n_4571),
.Y(n_5332)
);

AOI21xp5_ASAP7_75t_L g5333 ( 
.A1(n_4802),
.A2(n_2350),
.B(n_2321),
.Y(n_5333)
);

AOI22xp5_ASAP7_75t_L g5334 ( 
.A1(n_4730),
.A2(n_1963),
.B1(n_1964),
.B2(n_1959),
.Y(n_5334)
);

AND2x4_ASAP7_75t_L g5335 ( 
.A(n_4660),
.B(n_1963),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_4587),
.A2(n_2350),
.B(n_2321),
.Y(n_5336)
);

AND2x2_ASAP7_75t_SL g5337 ( 
.A(n_4764),
.B(n_4836),
.Y(n_5337)
);

BUFx4f_ASAP7_75t_L g5338 ( 
.A(n_4611),
.Y(n_5338)
);

OR2x2_ASAP7_75t_SL g5339 ( 
.A(n_4764),
.B(n_35),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_4648),
.Y(n_5340)
);

AOI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_4856),
.A2(n_2350),
.B(n_2321),
.Y(n_5341)
);

INVx2_ASAP7_75t_L g5342 ( 
.A(n_4983),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4648),
.Y(n_5343)
);

CKINVDCx20_ASAP7_75t_R g5344 ( 
.A(n_4754),
.Y(n_5344)
);

INVxp67_ASAP7_75t_SL g5345 ( 
.A(n_4791),
.Y(n_5345)
);

OAI22xp5_ASAP7_75t_L g5346 ( 
.A1(n_4894),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_5346)
);

HB1xp67_ASAP7_75t_L g5347 ( 
.A(n_4582),
.Y(n_5347)
);

HB1xp67_ASAP7_75t_L g5348 ( 
.A(n_4828),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4648),
.Y(n_5349)
);

A2O1A1Ixp33_ASAP7_75t_L g5350 ( 
.A1(n_4784),
.A2(n_125),
.B(n_127),
.C(n_124),
.Y(n_5350)
);

AND2x4_ASAP7_75t_L g5351 ( 
.A(n_4660),
.B(n_1964),
.Y(n_5351)
);

BUFx12f_ASAP7_75t_L g5352 ( 
.A(n_4896),
.Y(n_5352)
);

CKINVDCx5p33_ASAP7_75t_R g5353 ( 
.A(n_4607),
.Y(n_5353)
);

AOI22xp33_ASAP7_75t_L g5354 ( 
.A1(n_4872),
.A2(n_4950),
.B1(n_4917),
.B2(n_4852),
.Y(n_5354)
);

NOR2xp67_ASAP7_75t_R g5355 ( 
.A(n_4925),
.B(n_1964),
.Y(n_5355)
);

AND2x2_ASAP7_75t_SL g5356 ( 
.A(n_4836),
.B(n_4746),
.Y(n_5356)
);

OR2x2_ASAP7_75t_L g5357 ( 
.A(n_4750),
.B(n_124),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_4926),
.Y(n_5358)
);

BUFx3_ASAP7_75t_L g5359 ( 
.A(n_4896),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_4750),
.B(n_36),
.Y(n_5360)
);

INVx6_ASAP7_75t_L g5361 ( 
.A(n_4759),
.Y(n_5361)
);

INVx2_ASAP7_75t_L g5362 ( 
.A(n_4969),
.Y(n_5362)
);

OR2x2_ASAP7_75t_L g5363 ( 
.A(n_4894),
.B(n_127),
.Y(n_5363)
);

AOI22xp5_ASAP7_75t_L g5364 ( 
.A1(n_4857),
.A2(n_1972),
.B1(n_1975),
.B2(n_1964),
.Y(n_5364)
);

AND2x2_ASAP7_75t_L g5365 ( 
.A(n_4620),
.B(n_131),
.Y(n_5365)
);

BUFx2_ASAP7_75t_L g5366 ( 
.A(n_4611),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_4608),
.Y(n_5367)
);

INVxp67_ASAP7_75t_L g5368 ( 
.A(n_4610),
.Y(n_5368)
);

INVx2_ASAP7_75t_L g5369 ( 
.A(n_4969),
.Y(n_5369)
);

NAND2xp5_ASAP7_75t_L g5370 ( 
.A(n_4795),
.B(n_37),
.Y(n_5370)
);

AND2x6_ASAP7_75t_L g5371 ( 
.A(n_4791),
.B(n_1972),
.Y(n_5371)
);

AND2x2_ASAP7_75t_L g5372 ( 
.A(n_4795),
.B(n_131),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_4837),
.B(n_132),
.Y(n_5373)
);

INVx2_ASAP7_75t_L g5374 ( 
.A(n_4969),
.Y(n_5374)
);

AND2x4_ASAP7_75t_L g5375 ( 
.A(n_4711),
.B(n_1972),
.Y(n_5375)
);

INVx3_ASAP7_75t_L g5376 ( 
.A(n_4953),
.Y(n_5376)
);

O2A1O1Ixp33_ASAP7_75t_L g5377 ( 
.A1(n_4790),
.A2(n_42),
.B(n_39),
.C(n_40),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_4837),
.B(n_39),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_SL g5379 ( 
.A(n_4842),
.B(n_4799),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_4842),
.B(n_39),
.Y(n_5380)
);

OAI22xp5_ASAP7_75t_L g5381 ( 
.A1(n_4848),
.A2(n_45),
.B1(n_40),
.B2(n_43),
.Y(n_5381)
);

AND2x4_ASAP7_75t_L g5382 ( 
.A(n_4743),
.B(n_1972),
.Y(n_5382)
);

BUFx8_ASAP7_75t_SL g5383 ( 
.A(n_4909),
.Y(n_5383)
);

OAI22xp5_ASAP7_75t_L g5384 ( 
.A1(n_4848),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_5384)
);

CKINVDCx20_ASAP7_75t_R g5385 ( 
.A(n_4808),
.Y(n_5385)
);

CKINVDCx5p33_ASAP7_75t_R g5386 ( 
.A(n_4831),
.Y(n_5386)
);

AND2x2_ASAP7_75t_L g5387 ( 
.A(n_4845),
.B(n_132),
.Y(n_5387)
);

BUFx2_ASAP7_75t_L g5388 ( 
.A(n_4962),
.Y(n_5388)
);

AND2x2_ASAP7_75t_L g5389 ( 
.A(n_4845),
.B(n_133),
.Y(n_5389)
);

OAI21x1_ASAP7_75t_L g5390 ( 
.A1(n_4760),
.A2(n_2066),
.B(n_2060),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_4799),
.B(n_46),
.Y(n_5391)
);

BUFx2_ASAP7_75t_SL g5392 ( 
.A(n_4999),
.Y(n_5392)
);

INVx1_ASAP7_75t_SL g5393 ( 
.A(n_5018),
.Y(n_5393)
);

AOI22xp5_ASAP7_75t_L g5394 ( 
.A1(n_4989),
.A2(n_4679),
.B1(n_4811),
.B2(n_4717),
.Y(n_5394)
);

BUFx12f_ASAP7_75t_L g5395 ( 
.A(n_5020),
.Y(n_5395)
);

AOI22xp33_ASAP7_75t_SL g5396 ( 
.A1(n_5185),
.A2(n_4826),
.B1(n_4925),
.B2(n_4811),
.Y(n_5396)
);

OAI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5339),
.A2(n_4815),
.B1(n_4925),
.B2(n_4576),
.Y(n_5397)
);

OAI22xp33_ASAP7_75t_L g5398 ( 
.A1(n_4991),
.A2(n_4649),
.B1(n_4676),
.B2(n_4817),
.Y(n_5398)
);

AOI22xp33_ASAP7_75t_SL g5399 ( 
.A1(n_5185),
.A2(n_4826),
.B1(n_4866),
.B2(n_4843),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_4988),
.Y(n_5400)
);

AOI21xp33_ASAP7_75t_L g5401 ( 
.A1(n_4991),
.A2(n_4913),
.B(n_4700),
.Y(n_5401)
);

OAI22xp33_ASAP7_75t_L g5402 ( 
.A1(n_5182),
.A2(n_4668),
.B1(n_4885),
.B2(n_4971),
.Y(n_5402)
);

OAI22xp5_ASAP7_75t_L g5403 ( 
.A1(n_5130),
.A2(n_5045),
.B1(n_5277),
.B2(n_5139),
.Y(n_5403)
);

INVx2_ASAP7_75t_L g5404 ( 
.A(n_5005),
.Y(n_5404)
);

AOI22xp33_ASAP7_75t_SL g5405 ( 
.A1(n_5037),
.A2(n_4866),
.B1(n_4843),
.B2(n_4578),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_L g5406 ( 
.A(n_4987),
.B(n_4853),
.Y(n_5406)
);

INVx8_ASAP7_75t_L g5407 ( 
.A(n_5239),
.Y(n_5407)
);

INVx1_ASAP7_75t_SL g5408 ( 
.A(n_5018),
.Y(n_5408)
);

INVx1_ASAP7_75t_SL g5409 ( 
.A(n_5090),
.Y(n_5409)
);

CKINVDCx6p67_ASAP7_75t_R g5410 ( 
.A(n_5007),
.Y(n_5410)
);

AOI22xp33_ASAP7_75t_L g5411 ( 
.A1(n_5272),
.A2(n_4847),
.B1(n_4855),
.B2(n_4978),
.Y(n_5411)
);

BUFx3_ASAP7_75t_L g5412 ( 
.A(n_5154),
.Y(n_5412)
);

AOI22xp33_ASAP7_75t_L g5413 ( 
.A1(n_5056),
.A2(n_4847),
.B1(n_4855),
.B2(n_4978),
.Y(n_5413)
);

INVx4_ASAP7_75t_L g5414 ( 
.A(n_5237),
.Y(n_5414)
);

INVxp67_ASAP7_75t_SL g5415 ( 
.A(n_4987),
.Y(n_5415)
);

AOI22xp33_ASAP7_75t_L g5416 ( 
.A1(n_5140),
.A2(n_4728),
.B1(n_4937),
.B2(n_4699),
.Y(n_5416)
);

AOI22xp33_ASAP7_75t_L g5417 ( 
.A1(n_5208),
.A2(n_4728),
.B1(n_4699),
.B2(n_4688),
.Y(n_5417)
);

INVx1_ASAP7_75t_SL g5418 ( 
.A(n_5090),
.Y(n_5418)
);

BUFx3_ASAP7_75t_L g5419 ( 
.A(n_5038),
.Y(n_5419)
);

BUFx4_ASAP7_75t_R g5420 ( 
.A(n_5383),
.Y(n_5420)
);

CKINVDCx20_ASAP7_75t_R g5421 ( 
.A(n_5134),
.Y(n_5421)
);

INVxp67_ASAP7_75t_SL g5422 ( 
.A(n_5016),
.Y(n_5422)
);

INVx6_ASAP7_75t_L g5423 ( 
.A(n_5035),
.Y(n_5423)
);

BUFx4f_ASAP7_75t_SL g5424 ( 
.A(n_5042),
.Y(n_5424)
);

BUFx3_ASAP7_75t_L g5425 ( 
.A(n_5085),
.Y(n_5425)
);

INVx4_ASAP7_75t_L g5426 ( 
.A(n_5237),
.Y(n_5426)
);

INVx1_ASAP7_75t_SL g5427 ( 
.A(n_5273),
.Y(n_5427)
);

AOI22xp33_ASAP7_75t_SL g5428 ( 
.A1(n_5037),
.A2(n_4591),
.B1(n_4705),
.B2(n_4860),
.Y(n_5428)
);

INVx6_ASAP7_75t_L g5429 ( 
.A(n_5035),
.Y(n_5429)
);

BUFx2_ASAP7_75t_L g5430 ( 
.A(n_5013),
.Y(n_5430)
);

INVx4_ASAP7_75t_L g5431 ( 
.A(n_5237),
.Y(n_5431)
);

AOI22xp33_ASAP7_75t_SL g5432 ( 
.A1(n_5245),
.A2(n_5014),
.B1(n_5101),
.B2(n_5205),
.Y(n_5432)
);

CKINVDCx20_ASAP7_75t_R g5433 ( 
.A(n_5036),
.Y(n_5433)
);

CKINVDCx11_ASAP7_75t_R g5434 ( 
.A(n_5201),
.Y(n_5434)
);

BUFx3_ASAP7_75t_L g5435 ( 
.A(n_5222),
.Y(n_5435)
);

BUFx2_ASAP7_75t_L g5436 ( 
.A(n_4990),
.Y(n_5436)
);

BUFx2_ASAP7_75t_L g5437 ( 
.A(n_5046),
.Y(n_5437)
);

AOI22xp5_ASAP7_75t_L g5438 ( 
.A1(n_5208),
.A2(n_4860),
.B1(n_4688),
.B2(n_4705),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_4998),
.Y(n_5439)
);

CKINVDCx20_ASAP7_75t_R g5440 ( 
.A(n_5211),
.Y(n_5440)
);

OAI22xp5_ASAP7_75t_SL g5441 ( 
.A1(n_5344),
.A2(n_5321),
.B1(n_5385),
.B2(n_5325),
.Y(n_5441)
);

BUFx8_ASAP7_75t_L g5442 ( 
.A(n_5218),
.Y(n_5442)
);

BUFx12f_ASAP7_75t_L g5443 ( 
.A(n_5159),
.Y(n_5443)
);

OAI22xp33_ASAP7_75t_L g5444 ( 
.A1(n_5182),
.A2(n_4738),
.B1(n_4727),
.B2(n_4888),
.Y(n_5444)
);

OAI22xp33_ASAP7_75t_L g5445 ( 
.A1(n_5182),
.A2(n_5277),
.B1(n_5311),
.B2(n_5205),
.Y(n_5445)
);

BUFx3_ASAP7_75t_L g5446 ( 
.A(n_5196),
.Y(n_5446)
);

INVx6_ASAP7_75t_L g5447 ( 
.A(n_5146),
.Y(n_5447)
);

INVx1_ASAP7_75t_SL g5448 ( 
.A(n_5273),
.Y(n_5448)
);

INVx2_ASAP7_75t_L g5449 ( 
.A(n_5006),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_L g5450 ( 
.A(n_5040),
.B(n_5096),
.Y(n_5450)
);

AOI22xp5_ASAP7_75t_L g5451 ( 
.A1(n_5108),
.A2(n_4899),
.B1(n_4892),
.B2(n_4692),
.Y(n_5451)
);

INVx6_ASAP7_75t_L g5452 ( 
.A(n_5146),
.Y(n_5452)
);

BUFx3_ASAP7_75t_L g5453 ( 
.A(n_5225),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5002),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_5026),
.Y(n_5455)
);

INVx2_ASAP7_75t_L g5456 ( 
.A(n_5129),
.Y(n_5456)
);

BUFx6f_ASAP7_75t_L g5457 ( 
.A(n_5141),
.Y(n_5457)
);

AOI22xp33_ASAP7_75t_L g5458 ( 
.A1(n_5108),
.A2(n_4875),
.B1(n_4692),
.B2(n_4691),
.Y(n_5458)
);

AOI22xp5_ASAP7_75t_L g5459 ( 
.A1(n_5320),
.A2(n_4691),
.B1(n_4779),
.B2(n_4908),
.Y(n_5459)
);

OAI22xp5_ASAP7_75t_L g5460 ( 
.A1(n_5219),
.A2(n_5242),
.B1(n_5106),
.B2(n_5354),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_SL g5461 ( 
.A1(n_5245),
.A2(n_4922),
.B1(n_4924),
.B2(n_4634),
.Y(n_5461)
);

AOI22xp33_ASAP7_75t_L g5462 ( 
.A1(n_5256),
.A2(n_5189),
.B1(n_5095),
.B2(n_5098),
.Y(n_5462)
);

BUFx2_ASAP7_75t_SL g5463 ( 
.A(n_5166),
.Y(n_5463)
);

BUFx10_ASAP7_75t_L g5464 ( 
.A(n_5361),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5004),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_5353),
.Y(n_5466)
);

AOI22xp33_ASAP7_75t_L g5467 ( 
.A1(n_5256),
.A2(n_4954),
.B1(n_4779),
.B2(n_4766),
.Y(n_5467)
);

INVx1_ASAP7_75t_SL g5468 ( 
.A(n_5171),
.Y(n_5468)
);

INVx6_ASAP7_75t_L g5469 ( 
.A(n_5141),
.Y(n_5469)
);

AOI22xp5_ASAP7_75t_L g5470 ( 
.A1(n_5320),
.A2(n_4922),
.B1(n_4972),
.B2(n_4977),
.Y(n_5470)
);

BUFx12f_ASAP7_75t_L g5471 ( 
.A(n_5361),
.Y(n_5471)
);

AOI22xp33_ASAP7_75t_SL g5472 ( 
.A1(n_5101),
.A2(n_4634),
.B1(n_4851),
.B2(n_4840),
.Y(n_5472)
);

INVx4_ASAP7_75t_L g5473 ( 
.A(n_5246),
.Y(n_5473)
);

AOI22xp5_ASAP7_75t_L g5474 ( 
.A1(n_5067),
.A2(n_4704),
.B1(n_4703),
.B2(n_4712),
.Y(n_5474)
);

AOI22xp33_ASAP7_75t_SL g5475 ( 
.A1(n_5067),
.A2(n_5356),
.B1(n_5337),
.B2(n_5346),
.Y(n_5475)
);

INVx11_ASAP7_75t_L g5476 ( 
.A(n_5248),
.Y(n_5476)
);

CKINVDCx14_ASAP7_75t_R g5477 ( 
.A(n_5156),
.Y(n_5477)
);

AOI22xp33_ASAP7_75t_SL g5478 ( 
.A1(n_5346),
.A2(n_5384),
.B1(n_5381),
.B2(n_5119),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5008),
.Y(n_5479)
);

OAI22xp33_ASAP7_75t_L g5480 ( 
.A1(n_5098),
.A2(n_4713),
.B1(n_4870),
.B2(n_4655),
.Y(n_5480)
);

INVxp67_ASAP7_75t_SL g5481 ( 
.A(n_4996),
.Y(n_5481)
);

AOI22x1_ASAP7_75t_L g5482 ( 
.A1(n_5345),
.A2(n_4749),
.B1(n_4724),
.B2(n_4667),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5331),
.B(n_4608),
.Y(n_5483)
);

CKINVDCx6p67_ASAP7_75t_R g5484 ( 
.A(n_5010),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5017),
.Y(n_5485)
);

INVx1_ASAP7_75t_SL g5486 ( 
.A(n_5171),
.Y(n_5486)
);

INVx2_ASAP7_75t_SL g5487 ( 
.A(n_5167),
.Y(n_5487)
);

INVx1_ASAP7_75t_SL g5488 ( 
.A(n_4996),
.Y(n_5488)
);

NAND2x1p5_ASAP7_75t_L g5489 ( 
.A(n_5025),
.B(n_4832),
.Y(n_5489)
);

INVx1_ASAP7_75t_SL g5490 ( 
.A(n_5109),
.Y(n_5490)
);

INVx3_ASAP7_75t_SL g5491 ( 
.A(n_5386),
.Y(n_5491)
);

INVx1_ASAP7_75t_L g5492 ( 
.A(n_5023),
.Y(n_5492)
);

AOI22xp33_ASAP7_75t_L g5493 ( 
.A1(n_5009),
.A2(n_4682),
.B1(n_4689),
.B2(n_4672),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5011),
.B(n_4608),
.Y(n_5494)
);

AOI22xp33_ASAP7_75t_L g5495 ( 
.A1(n_5009),
.A2(n_4893),
.B1(n_4586),
.B2(n_4985),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_5024),
.Y(n_5496)
);

AOI22xp33_ASAP7_75t_SL g5497 ( 
.A1(n_5381),
.A2(n_4967),
.B1(n_4581),
.B2(n_4574),
.Y(n_5497)
);

AOI22xp33_ASAP7_75t_L g5498 ( 
.A1(n_5184),
.A2(n_4825),
.B1(n_4881),
.B2(n_4787),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5029),
.Y(n_5499)
);

AOI22xp33_ASAP7_75t_L g5500 ( 
.A1(n_5227),
.A2(n_5308),
.B1(n_5298),
.B2(n_5309),
.Y(n_5500)
);

AOI22xp5_ASAP7_75t_L g5501 ( 
.A1(n_5234),
.A2(n_5384),
.B1(n_5052),
.B2(n_5252),
.Y(n_5501)
);

INVx2_ASAP7_75t_SL g5502 ( 
.A(n_4986),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5033),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_5297),
.Y(n_5504)
);

AOI22xp33_ASAP7_75t_SL g5505 ( 
.A1(n_5234),
.A2(n_4678),
.B1(n_4621),
.B2(n_4884),
.Y(n_5505)
);

INVx1_ASAP7_75t_SL g5506 ( 
.A(n_5180),
.Y(n_5506)
);

INVx1_ASAP7_75t_SL g5507 ( 
.A(n_5183),
.Y(n_5507)
);

CKINVDCx11_ASAP7_75t_R g5508 ( 
.A(n_5010),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_5028),
.Y(n_5509)
);

NAND2x1p5_ASAP7_75t_L g5510 ( 
.A(n_5025),
.B(n_4819),
.Y(n_5510)
);

AOI22xp33_ASAP7_75t_L g5511 ( 
.A1(n_5309),
.A2(n_5322),
.B1(n_5063),
.B2(n_5323),
.Y(n_5511)
);

BUFx6f_ASAP7_75t_L g5512 ( 
.A(n_5141),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5100),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5104),
.Y(n_5514)
);

OAI21xp5_ASAP7_75t_SL g5515 ( 
.A1(n_5293),
.A2(n_4933),
.B(n_4910),
.Y(n_5515)
);

OAI22xp33_ASAP7_75t_L g5516 ( 
.A1(n_5078),
.A2(n_4867),
.B1(n_4753),
.B2(n_4935),
.Y(n_5516)
);

BUFx3_ASAP7_75t_L g5517 ( 
.A(n_5263),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5043),
.Y(n_5518)
);

AND2x2_ASAP7_75t_L g5519 ( 
.A(n_5126),
.B(n_4828),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_SL g5520 ( 
.A1(n_5062),
.A2(n_4889),
.B1(n_4767),
.B2(n_4803),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_5058),
.Y(n_5521)
);

OAI22xp33_ASAP7_75t_L g5522 ( 
.A1(n_5078),
.A2(n_4627),
.B1(n_4828),
.B2(n_4833),
.Y(n_5522)
);

BUFx6f_ASAP7_75t_SL g5523 ( 
.A(n_5032),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5064),
.Y(n_5524)
);

BUFx8_ASAP7_75t_SL g5525 ( 
.A(n_5066),
.Y(n_5525)
);

CKINVDCx11_ASAP7_75t_R g5526 ( 
.A(n_5332),
.Y(n_5526)
);

AOI22xp33_ASAP7_75t_L g5527 ( 
.A1(n_5309),
.A2(n_4873),
.B1(n_4882),
.B2(n_4869),
.Y(n_5527)
);

AOI22xp33_ASAP7_75t_L g5528 ( 
.A1(n_5322),
.A2(n_4859),
.B1(n_4822),
.B2(n_4794),
.Y(n_5528)
);

AND2x2_ASAP7_75t_L g5529 ( 
.A(n_5292),
.B(n_4615),
.Y(n_5529)
);

OAI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_5055),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5326),
.B(n_4833),
.Y(n_5531)
);

AOI22xp33_ASAP7_75t_SL g5532 ( 
.A1(n_5131),
.A2(n_4789),
.B1(n_4618),
.B2(n_4669),
.Y(n_5532)
);

BUFx6f_ASAP7_75t_L g5533 ( 
.A(n_4986),
.Y(n_5533)
);

AOI22xp33_ASAP7_75t_L g5534 ( 
.A1(n_5322),
.A2(n_4683),
.B1(n_4677),
.B2(n_4792),
.Y(n_5534)
);

BUFx12f_ASAP7_75t_L g5535 ( 
.A(n_5111),
.Y(n_5535)
);

AOI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_5063),
.A2(n_1972),
.B1(n_1976),
.B2(n_1975),
.Y(n_5536)
);

CKINVDCx11_ASAP7_75t_R g5537 ( 
.A(n_4986),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5071),
.Y(n_5538)
);

OAI22xp5_ASAP7_75t_L g5539 ( 
.A1(n_5055),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_5539)
);

AND2x4_ASAP7_75t_SL g5540 ( 
.A(n_5213),
.B(n_1975),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5072),
.Y(n_5541)
);

INVx3_ASAP7_75t_L g5542 ( 
.A(n_5066),
.Y(n_5542)
);

INVx6_ASAP7_75t_L g5543 ( 
.A(n_4995),
.Y(n_5543)
);

AOI22xp33_ASAP7_75t_L g5544 ( 
.A1(n_5132),
.A2(n_1975),
.B1(n_1987),
.B2(n_1976),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_5074),
.Y(n_5545)
);

CKINVDCx6p67_ASAP7_75t_R g5546 ( 
.A(n_5271),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5080),
.Y(n_5547)
);

AND2x2_ASAP7_75t_L g5548 ( 
.A(n_5303),
.B(n_4615),
.Y(n_5548)
);

AOI22xp33_ASAP7_75t_L g5549 ( 
.A1(n_5368),
.A2(n_1975),
.B1(n_1987),
.B2(n_1976),
.Y(n_5549)
);

AOI22xp33_ASAP7_75t_L g5550 ( 
.A1(n_5012),
.A2(n_5136),
.B1(n_5312),
.B2(n_5342),
.Y(n_5550)
);

INVx8_ASAP7_75t_L g5551 ( 
.A(n_5032),
.Y(n_5551)
);

CKINVDCx11_ASAP7_75t_R g5552 ( 
.A(n_4995),
.Y(n_5552)
);

INVx3_ASAP7_75t_L g5553 ( 
.A(n_5070),
.Y(n_5553)
);

BUFx2_ASAP7_75t_L g5554 ( 
.A(n_5070),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_5082),
.Y(n_5555)
);

OAI22xp5_ASAP7_75t_L g5556 ( 
.A1(n_5310),
.A2(n_4833),
.B1(n_58),
.B2(n_66),
.Y(n_5556)
);

INVx2_ASAP7_75t_L g5557 ( 
.A(n_5048),
.Y(n_5557)
);

AOI21xp5_ASAP7_75t_L g5558 ( 
.A1(n_5031),
.A2(n_4710),
.B(n_4709),
.Y(n_5558)
);

NAND2xp5_ASAP7_75t_L g5559 ( 
.A(n_5121),
.B(n_4615),
.Y(n_5559)
);

CKINVDCx11_ASAP7_75t_R g5560 ( 
.A(n_4995),
.Y(n_5560)
);

BUFx6f_ASAP7_75t_L g5561 ( 
.A(n_5027),
.Y(n_5561)
);

AND2x2_ASAP7_75t_L g5562 ( 
.A(n_5051),
.B(n_4597),
.Y(n_5562)
);

BUFx6f_ASAP7_75t_L g5563 ( 
.A(n_5027),
.Y(n_5563)
);

BUFx10_ASAP7_75t_L g5564 ( 
.A(n_5347),
.Y(n_5564)
);

BUFx6f_ASAP7_75t_L g5565 ( 
.A(n_5027),
.Y(n_5565)
);

CKINVDCx16_ASAP7_75t_R g5566 ( 
.A(n_5176),
.Y(n_5566)
);

INVx1_ASAP7_75t_SL g5567 ( 
.A(n_5186),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5076),
.Y(n_5568)
);

BUFx3_ASAP7_75t_L g5569 ( 
.A(n_5084),
.Y(n_5569)
);

BUFx3_ASAP7_75t_L g5570 ( 
.A(n_5084),
.Y(n_5570)
);

AOI22xp33_ASAP7_75t_L g5571 ( 
.A1(n_5128),
.A2(n_1976),
.B1(n_1987),
.B2(n_4674),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_5079),
.Y(n_5572)
);

BUFx12f_ASAP7_75t_L g5573 ( 
.A(n_5238),
.Y(n_5573)
);

BUFx4f_ASAP7_75t_L g5574 ( 
.A(n_5123),
.Y(n_5574)
);

BUFx10_ASAP7_75t_L g5575 ( 
.A(n_5122),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_5088),
.Y(n_5576)
);

BUFx3_ASAP7_75t_L g5577 ( 
.A(n_5084),
.Y(n_5577)
);

CKINVDCx20_ASAP7_75t_R g5578 ( 
.A(n_5324),
.Y(n_5578)
);

BUFx12f_ASAP7_75t_L g5579 ( 
.A(n_5120),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5103),
.Y(n_5580)
);

AOI22xp33_ASAP7_75t_L g5581 ( 
.A1(n_5128),
.A2(n_1976),
.B1(n_1987),
.B2(n_4646),
.Y(n_5581)
);

BUFx10_ASAP7_75t_L g5582 ( 
.A(n_5335),
.Y(n_5582)
);

AOI22xp5_ASAP7_75t_L g5583 ( 
.A1(n_5086),
.A2(n_4898),
.B1(n_4911),
.B2(n_4918),
.Y(n_5583)
);

BUFx8_ASAP7_75t_L g5584 ( 
.A(n_5169),
.Y(n_5584)
);

INVx5_ASAP7_75t_L g5585 ( 
.A(n_5230),
.Y(n_5585)
);

BUFx3_ASAP7_75t_L g5586 ( 
.A(n_5112),
.Y(n_5586)
);

BUFx3_ASAP7_75t_L g5587 ( 
.A(n_5112),
.Y(n_5587)
);

BUFx3_ASAP7_75t_L g5588 ( 
.A(n_5112),
.Y(n_5588)
);

INVx1_ASAP7_75t_SL g5589 ( 
.A(n_5233),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5103),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5149),
.Y(n_5591)
);

AOI22xp33_ASAP7_75t_L g5592 ( 
.A1(n_5128),
.A2(n_1987),
.B1(n_4652),
.B2(n_4722),
.Y(n_5592)
);

AOI22xp33_ASAP7_75t_L g5593 ( 
.A1(n_5294),
.A2(n_4765),
.B1(n_4659),
.B2(n_4664),
.Y(n_5593)
);

BUFx6f_ASAP7_75t_L g5594 ( 
.A(n_5127),
.Y(n_5594)
);

AOI22xp33_ASAP7_75t_L g5595 ( 
.A1(n_5327),
.A2(n_4773),
.B1(n_4775),
.B2(n_4642),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5147),
.Y(n_5596)
);

BUFx6f_ASAP7_75t_L g5597 ( 
.A(n_5127),
.Y(n_5597)
);

HB1xp67_ASAP7_75t_L g5598 ( 
.A(n_5105),
.Y(n_5598)
);

AOI22xp33_ASAP7_75t_L g5599 ( 
.A1(n_5086),
.A2(n_4769),
.B1(n_2014),
.B2(n_2021),
.Y(n_5599)
);

INVx6_ASAP7_75t_L g5600 ( 
.A(n_5127),
.Y(n_5600)
);

OAI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5061),
.A2(n_51),
.B1(n_47),
.B2(n_50),
.Y(n_5601)
);

AOI22xp33_ASAP7_75t_L g5602 ( 
.A1(n_5387),
.A2(n_2014),
.B1(n_2021),
.B2(n_2009),
.Y(n_5602)
);

BUFx8_ASAP7_75t_L g5603 ( 
.A(n_5054),
.Y(n_5603)
);

AOI22xp33_ASAP7_75t_SL g5604 ( 
.A1(n_5061),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_5604)
);

BUFx8_ASAP7_75t_L g5605 ( 
.A(n_5223),
.Y(n_5605)
);

AOI22xp33_ASAP7_75t_L g5606 ( 
.A1(n_5389),
.A2(n_2014),
.B1(n_2021),
.B2(n_2009),
.Y(n_5606)
);

CKINVDCx5p33_ASAP7_75t_R g5607 ( 
.A(n_5162),
.Y(n_5607)
);

OAI22xp33_ASAP7_75t_L g5608 ( 
.A1(n_5068),
.A2(n_56),
.B1(n_52),
.B2(n_54),
.Y(n_5608)
);

AOI22xp5_ASAP7_75t_L g5609 ( 
.A1(n_5379),
.A2(n_57),
.B1(n_58),
.B2(n_56),
.Y(n_5609)
);

INVx6_ASAP7_75t_L g5610 ( 
.A(n_5162),
.Y(n_5610)
);

NAND2xp5_ASAP7_75t_L g5611 ( 
.A(n_5194),
.B(n_133),
.Y(n_5611)
);

HB1xp67_ASAP7_75t_L g5612 ( 
.A(n_5147),
.Y(n_5612)
);

AOI22xp33_ASAP7_75t_SL g5613 ( 
.A1(n_5073),
.A2(n_57),
.B1(n_52),
.B2(n_56),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5158),
.Y(n_5614)
);

CKINVDCx11_ASAP7_75t_R g5615 ( 
.A(n_5290),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_L g5616 ( 
.A(n_5194),
.B(n_134),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5158),
.Y(n_5617)
);

INVx2_ASAP7_75t_L g5618 ( 
.A(n_5091),
.Y(n_5618)
);

CKINVDCx6p67_ASAP7_75t_R g5619 ( 
.A(n_5246),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5190),
.Y(n_5620)
);

INVx2_ASAP7_75t_L g5621 ( 
.A(n_5093),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5190),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_L g5623 ( 
.A1(n_5041),
.A2(n_2014),
.B1(n_2021),
.B2(n_2009),
.Y(n_5623)
);

INVx5_ASAP7_75t_L g5624 ( 
.A(n_5230),
.Y(n_5624)
);

CKINVDCx20_ASAP7_75t_R g5625 ( 
.A(n_5324),
.Y(n_5625)
);

INVx6_ASAP7_75t_L g5626 ( 
.A(n_5162),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5117),
.Y(n_5627)
);

OAI22xp5_ASAP7_75t_L g5628 ( 
.A1(n_5350),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_5628)
);

AOI22xp33_ASAP7_75t_L g5629 ( 
.A1(n_5160),
.A2(n_2014),
.B1(n_2021),
.B2(n_2009),
.Y(n_5629)
);

BUFx2_ASAP7_75t_L g5630 ( 
.A(n_5051),
.Y(n_5630)
);

CKINVDCx6p67_ASAP7_75t_R g5631 ( 
.A(n_5246),
.Y(n_5631)
);

NAND2xp5_ASAP7_75t_L g5632 ( 
.A(n_5198),
.B(n_134),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5152),
.Y(n_5633)
);

OAI22xp33_ASAP7_75t_L g5634 ( 
.A1(n_5068),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5118),
.Y(n_5635)
);

CKINVDCx16_ASAP7_75t_R g5636 ( 
.A(n_5274),
.Y(n_5636)
);

INVx5_ASAP7_75t_L g5637 ( 
.A(n_5230),
.Y(n_5637)
);

BUFx4f_ASAP7_75t_L g5638 ( 
.A(n_5290),
.Y(n_5638)
);

AOI22xp5_ASAP7_75t_L g5639 ( 
.A1(n_5206),
.A2(n_62),
.B1(n_63),
.B2(n_61),
.Y(n_5639)
);

BUFx4f_ASAP7_75t_SL g5640 ( 
.A(n_5075),
.Y(n_5640)
);

OAI22xp5_ASAP7_75t_L g5641 ( 
.A1(n_5357),
.A2(n_63),
.B1(n_59),
.B2(n_62),
.Y(n_5641)
);

AOI22xp33_ASAP7_75t_L g5642 ( 
.A1(n_5371),
.A2(n_2030),
.B1(n_2009),
.B2(n_2321),
.Y(n_5642)
);

NAND2xp5_ASAP7_75t_L g5643 ( 
.A(n_5209),
.B(n_135),
.Y(n_5643)
);

AND2x2_ASAP7_75t_L g5644 ( 
.A(n_5305),
.B(n_137),
.Y(n_5644)
);

INVxp67_ASAP7_75t_L g5645 ( 
.A(n_5021),
.Y(n_5645)
);

AOI22xp5_ASAP7_75t_SL g5646 ( 
.A1(n_5317),
.A2(n_71),
.B1(n_79),
.B2(n_63),
.Y(n_5646)
);

AOI22xp33_ASAP7_75t_L g5647 ( 
.A1(n_5371),
.A2(n_2030),
.B1(n_2350),
.B2(n_2321),
.Y(n_5647)
);

HB1xp67_ASAP7_75t_L g5648 ( 
.A(n_5102),
.Y(n_5648)
);

INVx3_ASAP7_75t_L g5649 ( 
.A(n_5282),
.Y(n_5649)
);

INVx2_ASAP7_75t_L g5650 ( 
.A(n_5152),
.Y(n_5650)
);

AOI22xp33_ASAP7_75t_SL g5651 ( 
.A1(n_4994),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_5651)
);

INVx6_ASAP7_75t_L g5652 ( 
.A(n_5178),
.Y(n_5652)
);

BUFx2_ASAP7_75t_L g5653 ( 
.A(n_5305),
.Y(n_5653)
);

CKINVDCx11_ASAP7_75t_R g5654 ( 
.A(n_5290),
.Y(n_5654)
);

AOI22xp33_ASAP7_75t_L g5655 ( 
.A1(n_5371),
.A2(n_2030),
.B1(n_2364),
.B2(n_2350),
.Y(n_5655)
);

BUFx12f_ASAP7_75t_L g5656 ( 
.A(n_5275),
.Y(n_5656)
);

OAI22xp33_ASAP7_75t_L g5657 ( 
.A1(n_5068),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_5657)
);

INVx4_ASAP7_75t_L g5658 ( 
.A(n_5178),
.Y(n_5658)
);

OAI22xp5_ASAP7_75t_L g5659 ( 
.A1(n_5262),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_5659)
);

AOI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5371),
.A2(n_2030),
.B1(n_2364),
.B2(n_2350),
.Y(n_5660)
);

AOI22xp5_ASAP7_75t_L g5661 ( 
.A1(n_5226),
.A2(n_70),
.B1(n_72),
.B2(n_69),
.Y(n_5661)
);

AOI22xp5_ASAP7_75t_L g5662 ( 
.A1(n_5365),
.A2(n_70),
.B1(n_72),
.B2(n_69),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5155),
.Y(n_5663)
);

INVx2_ASAP7_75t_SL g5664 ( 
.A(n_5178),
.Y(n_5664)
);

BUFx2_ASAP7_75t_L g5665 ( 
.A(n_5110),
.Y(n_5665)
);

CKINVDCx5p33_ASAP7_75t_R g5666 ( 
.A(n_5207),
.Y(n_5666)
);

INVx6_ASAP7_75t_L g5667 ( 
.A(n_5207),
.Y(n_5667)
);

NAND2xp5_ASAP7_75t_L g5668 ( 
.A(n_5015),
.B(n_139),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_5175),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_5372),
.A2(n_2030),
.B1(n_2372),
.B2(n_2364),
.Y(n_5670)
);

OAI22xp33_ASAP7_75t_L g5671 ( 
.A1(n_4993),
.A2(n_73),
.B1(n_68),
.B2(n_70),
.Y(n_5671)
);

AOI22xp33_ASAP7_75t_L g5672 ( 
.A1(n_5373),
.A2(n_2372),
.B1(n_2384),
.B2(n_2364),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5157),
.Y(n_5673)
);

INVx4_ASAP7_75t_L g5674 ( 
.A(n_5207),
.Y(n_5674)
);

BUFx10_ASAP7_75t_L g5675 ( 
.A(n_5335),
.Y(n_5675)
);

AOI22xp33_ASAP7_75t_L g5676 ( 
.A1(n_5254),
.A2(n_2372),
.B1(n_2384),
.B2(n_2364),
.Y(n_5676)
);

CKINVDCx11_ASAP7_75t_R g5677 ( 
.A(n_5220),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_5019),
.B(n_139),
.Y(n_5678)
);

NAND2x1p5_ASAP7_75t_L g5679 ( 
.A(n_5025),
.B(n_2364),
.Y(n_5679)
);

AOI22xp33_ASAP7_75t_L g5680 ( 
.A1(n_5053),
.A2(n_2384),
.B1(n_2388),
.B2(n_2372),
.Y(n_5680)
);

CKINVDCx11_ASAP7_75t_R g5681 ( 
.A(n_5220),
.Y(n_5681)
);

CKINVDCx11_ASAP7_75t_R g5682 ( 
.A(n_5220),
.Y(n_5682)
);

INVx1_ASAP7_75t_SL g5683 ( 
.A(n_5302),
.Y(n_5683)
);

BUFx2_ASAP7_75t_L g5684 ( 
.A(n_5282),
.Y(n_5684)
);

BUFx3_ASAP7_75t_L g5685 ( 
.A(n_5075),
.Y(n_5685)
);

INVx6_ASAP7_75t_L g5686 ( 
.A(n_5352),
.Y(n_5686)
);

AOI22xp33_ASAP7_75t_SL g5687 ( 
.A1(n_4993),
.A2(n_74),
.B1(n_68),
.B2(n_73),
.Y(n_5687)
);

INVx2_ASAP7_75t_L g5688 ( 
.A(n_5179),
.Y(n_5688)
);

INVx3_ASAP7_75t_L g5689 ( 
.A(n_5214),
.Y(n_5689)
);

AOI22xp33_ASAP7_75t_L g5690 ( 
.A1(n_5053),
.A2(n_2384),
.B1(n_2388),
.B2(n_2372),
.Y(n_5690)
);

CKINVDCx5p33_ASAP7_75t_R g5691 ( 
.A(n_5000),
.Y(n_5691)
);

CKINVDCx6p67_ASAP7_75t_R g5692 ( 
.A(n_5138),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5192),
.Y(n_5693)
);

INVx2_ASAP7_75t_L g5694 ( 
.A(n_5195),
.Y(n_5694)
);

AOI22xp33_ASAP7_75t_SL g5695 ( 
.A1(n_5177),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_5695)
);

OAI22xp5_ASAP7_75t_L g5696 ( 
.A1(n_5377),
.A2(n_82),
.B1(n_74),
.B2(n_76),
.Y(n_5696)
);

INVx3_ASAP7_75t_L g5697 ( 
.A(n_5214),
.Y(n_5697)
);

AOI22xp33_ASAP7_75t_SL g5698 ( 
.A1(n_4992),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_5698)
);

CKINVDCx20_ASAP7_75t_R g5699 ( 
.A(n_5324),
.Y(n_5699)
);

CKINVDCx11_ASAP7_75t_R g5700 ( 
.A(n_5200),
.Y(n_5700)
);

AOI22xp33_ASAP7_75t_SL g5701 ( 
.A1(n_5191),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5203),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5059),
.B(n_5021),
.Y(n_5703)
);

NAND2xp5_ASAP7_75t_L g5704 ( 
.A(n_5060),
.B(n_140),
.Y(n_5704)
);

OAI21xp5_ASAP7_75t_SL g5705 ( 
.A1(n_5261),
.A2(n_79),
.B(n_80),
.Y(n_5705)
);

AOI22xp33_ASAP7_75t_SL g5706 ( 
.A1(n_5191),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5163),
.Y(n_5707)
);

OAI22xp33_ASAP7_75t_L g5708 ( 
.A1(n_5053),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5172),
.Y(n_5709)
);

BUFx10_ASAP7_75t_L g5710 ( 
.A(n_5351),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5301),
.Y(n_5711)
);

OAI22xp5_ASAP7_75t_L g5712 ( 
.A1(n_5197),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5304),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5348),
.Y(n_5714)
);

BUFx3_ASAP7_75t_L g5715 ( 
.A(n_5161),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_5125),
.Y(n_5716)
);

OAI22xp5_ASAP7_75t_L g5717 ( 
.A1(n_5197),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5137),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5210),
.Y(n_5719)
);

CKINVDCx20_ASAP7_75t_R g5720 ( 
.A(n_5089),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5145),
.Y(n_5721)
);

AOI22xp33_ASAP7_75t_L g5722 ( 
.A1(n_5316),
.A2(n_2384),
.B1(n_2388),
.B2(n_2372),
.Y(n_5722)
);

BUFx2_ASAP7_75t_L g5723 ( 
.A(n_5217),
.Y(n_5723)
);

AOI22xp33_ASAP7_75t_L g5724 ( 
.A1(n_5363),
.A2(n_2388),
.B1(n_2398),
.B2(n_2384),
.Y(n_5724)
);

INVx6_ASAP7_75t_L g5725 ( 
.A(n_5295),
.Y(n_5725)
);

INVx5_ASAP7_75t_L g5726 ( 
.A(n_5174),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_5340),
.Y(n_5727)
);

AOI22xp5_ASAP7_75t_L g5728 ( 
.A1(n_5199),
.A2(n_88),
.B1(n_89),
.B2(n_87),
.Y(n_5728)
);

AOI22xp33_ASAP7_75t_L g5729 ( 
.A1(n_5280),
.A2(n_2398),
.B1(n_2426),
.B2(n_2388),
.Y(n_5729)
);

AOI22xp33_ASAP7_75t_SL g5730 ( 
.A1(n_5199),
.A2(n_88),
.B1(n_84),
.B2(n_87),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5343),
.Y(n_5731)
);

AOI22xp33_ASAP7_75t_L g5732 ( 
.A1(n_5097),
.A2(n_2398),
.B1(n_2426),
.B2(n_2388),
.Y(n_5732)
);

AOI22xp33_ASAP7_75t_L g5733 ( 
.A1(n_5097),
.A2(n_2426),
.B1(n_2428),
.B2(n_2398),
.Y(n_5733)
);

BUFx3_ASAP7_75t_L g5734 ( 
.A(n_5161),
.Y(n_5734)
);

NAND2x1p5_ASAP7_75t_L g5735 ( 
.A(n_5133),
.B(n_2398),
.Y(n_5735)
);

INVx1_ASAP7_75t_L g5736 ( 
.A(n_5349),
.Y(n_5736)
);

AND2x2_ASAP7_75t_L g5737 ( 
.A(n_5221),
.B(n_141),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_5224),
.Y(n_5738)
);

AOI22xp33_ASAP7_75t_SL g5739 ( 
.A1(n_5228),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_5739)
);

CKINVDCx20_ASAP7_75t_R g5740 ( 
.A(n_5421),
.Y(n_5740)
);

O2A1O1Ixp5_ASAP7_75t_L g5741 ( 
.A1(n_5403),
.A2(n_5001),
.B(n_5231),
.C(n_5228),
.Y(n_5741)
);

A2O1A1Ixp33_ASAP7_75t_L g5742 ( 
.A1(n_5705),
.A2(n_5646),
.B(n_5399),
.C(n_5501),
.Y(n_5742)
);

AND2x2_ASAP7_75t_L g5743 ( 
.A(n_5437),
.B(n_5313),
.Y(n_5743)
);

AND2x2_ASAP7_75t_L g5744 ( 
.A(n_5653),
.B(n_5313),
.Y(n_5744)
);

OAI22xp5_ASAP7_75t_L g5745 ( 
.A1(n_5396),
.A2(n_5240),
.B1(n_5315),
.B2(n_5314),
.Y(n_5745)
);

O2A1O1Ixp5_ASAP7_75t_L g5746 ( 
.A1(n_5712),
.A2(n_5231),
.B(n_5315),
.C(n_5314),
.Y(n_5746)
);

NAND2xp5_ASAP7_75t_L g5747 ( 
.A(n_5415),
.B(n_5367),
.Y(n_5747)
);

AND2x4_ASAP7_75t_L g5748 ( 
.A(n_5542),
.B(n_5244),
.Y(n_5748)
);

OAI22xp5_ASAP7_75t_L g5749 ( 
.A1(n_5478),
.A2(n_5360),
.B1(n_5391),
.B2(n_5165),
.Y(n_5749)
);

BUFx3_ASAP7_75t_L g5750 ( 
.A(n_5440),
.Y(n_5750)
);

AOI21x1_ASAP7_75t_SL g5751 ( 
.A1(n_5494),
.A2(n_5142),
.B(n_5138),
.Y(n_5751)
);

NOR2xp33_ASAP7_75t_L g5752 ( 
.A(n_5491),
.B(n_5142),
.Y(n_5752)
);

BUFx6f_ASAP7_75t_L g5753 ( 
.A(n_5434),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_SL g5754 ( 
.A1(n_5460),
.A2(n_5124),
.B(n_5065),
.Y(n_5754)
);

A2O1A1Ixp33_ASAP7_75t_SL g5755 ( 
.A1(n_5401),
.A2(n_5360),
.B(n_5391),
.C(n_5378),
.Y(n_5755)
);

AOI21xp5_ASAP7_75t_L g5756 ( 
.A1(n_5398),
.A2(n_5276),
.B(n_5039),
.Y(n_5756)
);

AND2x2_ASAP7_75t_L g5757 ( 
.A(n_5430),
.B(n_5257),
.Y(n_5757)
);

AOI21x1_ASAP7_75t_SL g5758 ( 
.A1(n_5483),
.A2(n_5050),
.B(n_5049),
.Y(n_5758)
);

NAND2xp5_ASAP7_75t_L g5759 ( 
.A(n_5481),
.B(n_5049),
.Y(n_5759)
);

AND2x2_ASAP7_75t_L g5760 ( 
.A(n_5436),
.B(n_5266),
.Y(n_5760)
);

A2O1A1Ixp33_ASAP7_75t_L g5761 ( 
.A1(n_5705),
.A2(n_5083),
.B(n_5113),
.C(n_5370),
.Y(n_5761)
);

HB1xp67_ASAP7_75t_L g5762 ( 
.A(n_5427),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5400),
.Y(n_5763)
);

AND2x2_ASAP7_75t_L g5764 ( 
.A(n_5409),
.B(n_5270),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5683),
.Y(n_5765)
);

HB1xp67_ASAP7_75t_L g5766 ( 
.A(n_5427),
.Y(n_5766)
);

OR2x2_ASAP7_75t_L g5767 ( 
.A(n_5612),
.B(n_5235),
.Y(n_5767)
);

BUFx6f_ASAP7_75t_L g5768 ( 
.A(n_5464),
.Y(n_5768)
);

OAI22xp5_ASAP7_75t_L g5769 ( 
.A1(n_5432),
.A2(n_5370),
.B1(n_5380),
.B2(n_5378),
.Y(n_5769)
);

AND2x4_ASAP7_75t_L g5770 ( 
.A(n_5542),
.B(n_5388),
.Y(n_5770)
);

AOI221x1_ASAP7_75t_SL g5771 ( 
.A1(n_5712),
.A2(n_5380),
.B1(n_5050),
.B2(n_89),
.C(n_5355),
.Y(n_5771)
);

AND2x2_ASAP7_75t_L g5772 ( 
.A(n_5409),
.B(n_5174),
.Y(n_5772)
);

AND2x2_ASAP7_75t_L g5773 ( 
.A(n_5418),
.B(n_5174),
.Y(n_5773)
);

OAI22xp5_ASAP7_75t_L g5774 ( 
.A1(n_5501),
.A2(n_5034),
.B1(n_5148),
.B2(n_5133),
.Y(n_5774)
);

INVx1_ASAP7_75t_SL g5775 ( 
.A(n_5683),
.Y(n_5775)
);

AOI21x1_ASAP7_75t_SL g5776 ( 
.A1(n_5611),
.A2(n_5092),
.B(n_5151),
.Y(n_5776)
);

AOI221x1_ASAP7_75t_SL g5777 ( 
.A1(n_5717),
.A2(n_5355),
.B1(n_145),
.B2(n_150),
.C(n_144),
.Y(n_5777)
);

CKINVDCx5p33_ASAP7_75t_R g5778 ( 
.A(n_5395),
.Y(n_5778)
);

AND2x2_ASAP7_75t_SL g5779 ( 
.A(n_5636),
.B(n_5338),
.Y(n_5779)
);

INVxp67_ASAP7_75t_SL g5780 ( 
.A(n_5648),
.Y(n_5780)
);

OR2x2_ASAP7_75t_L g5781 ( 
.A(n_5488),
.B(n_5241),
.Y(n_5781)
);

HB1xp67_ASAP7_75t_L g5782 ( 
.A(n_5448),
.Y(n_5782)
);

CKINVDCx16_ASAP7_75t_R g5783 ( 
.A(n_5433),
.Y(n_5783)
);

AOI21xp5_ASAP7_75t_L g5784 ( 
.A1(n_5413),
.A2(n_5116),
.B(n_5114),
.Y(n_5784)
);

AND2x2_ASAP7_75t_L g5785 ( 
.A(n_5418),
.B(n_5187),
.Y(n_5785)
);

BUFx6f_ASAP7_75t_L g5786 ( 
.A(n_5464),
.Y(n_5786)
);

BUFx2_ASAP7_75t_L g5787 ( 
.A(n_5477),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5630),
.B(n_5187),
.Y(n_5788)
);

O2A1O1Ixp33_ASAP7_75t_L g5789 ( 
.A1(n_5460),
.A2(n_5003),
.B(n_5030),
.C(n_5057),
.Y(n_5789)
);

NAND2xp5_ASAP7_75t_L g5790 ( 
.A(n_5488),
.B(n_5358),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5439),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5575),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_5448),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_5454),
.Y(n_5794)
);

AOI21xp5_ASAP7_75t_SL g5795 ( 
.A1(n_5397),
.A2(n_5402),
.B(n_5530),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5465),
.Y(n_5796)
);

O2A1O1Ixp5_ASAP7_75t_L g5797 ( 
.A1(n_5717),
.A2(n_5289),
.B(n_5251),
.C(n_5338),
.Y(n_5797)
);

OA21x2_ASAP7_75t_L g5798 ( 
.A1(n_5627),
.A2(n_5265),
.B(n_5260),
.Y(n_5798)
);

AND2x4_ASAP7_75t_L g5799 ( 
.A(n_5553),
.B(n_5232),
.Y(n_5799)
);

HB1xp67_ASAP7_75t_L g5800 ( 
.A(n_5468),
.Y(n_5800)
);

A2O1A1Ixp33_ASAP7_75t_L g5801 ( 
.A1(n_5646),
.A2(n_5258),
.B(n_5259),
.C(n_5285),
.Y(n_5801)
);

NOR2xp33_ASAP7_75t_R g5802 ( 
.A(n_5504),
.B(n_5232),
.Y(n_5802)
);

INVx1_ASAP7_75t_SL g5803 ( 
.A(n_5506),
.Y(n_5803)
);

OAI22xp5_ASAP7_75t_L g5804 ( 
.A1(n_5462),
.A2(n_5148),
.B1(n_5133),
.B2(n_5281),
.Y(n_5804)
);

AOI21xp5_ASAP7_75t_SL g5805 ( 
.A1(n_5397),
.A2(n_5168),
.B(n_5065),
.Y(n_5805)
);

OR2x2_ASAP7_75t_L g5806 ( 
.A(n_5596),
.B(n_5253),
.Y(n_5806)
);

HB1xp67_ASAP7_75t_L g5807 ( 
.A(n_5468),
.Y(n_5807)
);

NOR2xp67_ASAP7_75t_L g5808 ( 
.A(n_5726),
.B(n_5148),
.Y(n_5808)
);

O2A1O1Ixp5_ASAP7_75t_L g5809 ( 
.A1(n_5659),
.A2(n_5144),
.B(n_5150),
.C(n_5264),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5575),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5479),
.Y(n_5811)
);

OR2x2_ASAP7_75t_L g5812 ( 
.A(n_5614),
.B(n_5287),
.Y(n_5812)
);

OR2x2_ASAP7_75t_L g5813 ( 
.A(n_5617),
.B(n_5291),
.Y(n_5813)
);

INVxp67_ASAP7_75t_L g5814 ( 
.A(n_5422),
.Y(n_5814)
);

INVx2_ASAP7_75t_L g5815 ( 
.A(n_5513),
.Y(n_5815)
);

INVx1_ASAP7_75t_SL g5816 ( 
.A(n_5506),
.Y(n_5816)
);

AND2x2_ASAP7_75t_L g5817 ( 
.A(n_5490),
.B(n_5264),
.Y(n_5817)
);

AOI21xp5_ASAP7_75t_L g5818 ( 
.A1(n_5515),
.A2(n_5135),
.B(n_5204),
.Y(n_5818)
);

O2A1O1Ixp5_ASAP7_75t_L g5819 ( 
.A1(n_5659),
.A2(n_5445),
.B(n_5641),
.C(n_5601),
.Y(n_5819)
);

AND2x2_ASAP7_75t_L g5820 ( 
.A(n_5490),
.B(n_5366),
.Y(n_5820)
);

AOI21x1_ASAP7_75t_SL g5821 ( 
.A1(n_5616),
.A2(n_5151),
.B(n_5375),
.Y(n_5821)
);

A2O1A1Ixp33_ASAP7_75t_L g5822 ( 
.A1(n_5475),
.A2(n_5212),
.B(n_5243),
.C(n_5193),
.Y(n_5822)
);

NOR2xp67_ASAP7_75t_L g5823 ( 
.A(n_5726),
.B(n_5376),
.Y(n_5823)
);

NAND2xp5_ASAP7_75t_L g5824 ( 
.A(n_5620),
.B(n_5296),
.Y(n_5824)
);

OA21x2_ASAP7_75t_L g5825 ( 
.A1(n_5635),
.A2(n_5390),
.B(n_5329),
.Y(n_5825)
);

NAND2xp5_ASAP7_75t_L g5826 ( 
.A(n_5622),
.B(n_5362),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_5665),
.Y(n_5827)
);

AND2x2_ASAP7_75t_L g5828 ( 
.A(n_5486),
.B(n_5376),
.Y(n_5828)
);

AND2x2_ASAP7_75t_L g5829 ( 
.A(n_5486),
.B(n_5168),
.Y(n_5829)
);

AND2x4_ASAP7_75t_L g5830 ( 
.A(n_5553),
.B(n_5359),
.Y(n_5830)
);

NAND2xp5_ASAP7_75t_L g5831 ( 
.A(n_5393),
.B(n_5278),
.Y(n_5831)
);

NOR2xp67_ASAP7_75t_L g5832 ( 
.A(n_5726),
.B(n_5044),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5393),
.B(n_5283),
.Y(n_5833)
);

NAND2xp5_ASAP7_75t_L g5834 ( 
.A(n_5408),
.B(n_5306),
.Y(n_5834)
);

O2A1O1Ixp33_ASAP7_75t_L g5835 ( 
.A1(n_5628),
.A2(n_5087),
.B(n_5255),
.C(n_5247),
.Y(n_5835)
);

HB1xp67_ASAP7_75t_L g5836 ( 
.A(n_5408),
.Y(n_5836)
);

OA21x2_ASAP7_75t_L g5837 ( 
.A1(n_5673),
.A2(n_5328),
.B(n_5369),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5564),
.Y(n_5838)
);

INVxp67_ASAP7_75t_L g5839 ( 
.A(n_5703),
.Y(n_5839)
);

AOI21x1_ASAP7_75t_SL g5840 ( 
.A1(n_5406),
.A2(n_5382),
.B(n_5375),
.Y(n_5840)
);

BUFx2_ASAP7_75t_L g5841 ( 
.A(n_5554),
.Y(n_5841)
);

AOI21xp5_ASAP7_75t_SL g5842 ( 
.A1(n_5530),
.A2(n_5181),
.B(n_5267),
.Y(n_5842)
);

OA21x2_ASAP7_75t_L g5843 ( 
.A1(n_5707),
.A2(n_5374),
.B(n_5288),
.Y(n_5843)
);

HB1xp67_ASAP7_75t_L g5844 ( 
.A(n_5580),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5485),
.Y(n_5845)
);

AOI21x1_ASAP7_75t_SL g5846 ( 
.A1(n_5559),
.A2(n_5382),
.B(n_5094),
.Y(n_5846)
);

OAI22xp5_ASAP7_75t_L g5847 ( 
.A1(n_5411),
.A2(n_5281),
.B1(n_5115),
.B2(n_5181),
.Y(n_5847)
);

A2O1A1Ixp33_ASAP7_75t_L g5848 ( 
.A1(n_5662),
.A2(n_5115),
.B(n_5173),
.C(n_5153),
.Y(n_5848)
);

INVx1_ASAP7_75t_SL g5849 ( 
.A(n_5507),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5492),
.Y(n_5850)
);

OA21x2_ASAP7_75t_L g5851 ( 
.A1(n_5709),
.A2(n_5341),
.B(n_4997),
.Y(n_5851)
);

O2A1O1Ixp5_ASAP7_75t_L g5852 ( 
.A1(n_5641),
.A2(n_5047),
.B(n_5069),
.C(n_5077),
.Y(n_5852)
);

NOR3xp33_ASAP7_75t_L g5853 ( 
.A(n_5405),
.B(n_5107),
.C(n_5022),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5723),
.B(n_5267),
.Y(n_5854)
);

INVx2_ASAP7_75t_L g5855 ( 
.A(n_5564),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5684),
.B(n_5170),
.Y(n_5856)
);

BUFx2_ASAP7_75t_L g5857 ( 
.A(n_5685),
.Y(n_5857)
);

AOI21xp5_ASAP7_75t_L g5858 ( 
.A1(n_5515),
.A2(n_5307),
.B(n_5284),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5499),
.Y(n_5859)
);

O2A1O1Ixp33_ASAP7_75t_L g5860 ( 
.A1(n_5628),
.A2(n_5351),
.B(n_5077),
.C(n_5094),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5507),
.B(n_5170),
.Y(n_5861)
);

AND2x4_ASAP7_75t_L g5862 ( 
.A(n_5567),
.B(n_5188),
.Y(n_5862)
);

OAI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_5662),
.A2(n_5099),
.B1(n_5364),
.B2(n_5334),
.Y(n_5863)
);

NAND2xp5_ASAP7_75t_L g5864 ( 
.A(n_5590),
.B(n_5299),
.Y(n_5864)
);

NOR2xp67_ASAP7_75t_L g5865 ( 
.A(n_5471),
.B(n_5300),
.Y(n_5865)
);

O2A1O1Ixp33_ASAP7_75t_L g5866 ( 
.A1(n_5696),
.A2(n_5153),
.B(n_5173),
.C(n_5330),
.Y(n_5866)
);

BUFx3_ASAP7_75t_L g5867 ( 
.A(n_5443),
.Y(n_5867)
);

NAND2xp5_ASAP7_75t_L g5868 ( 
.A(n_5518),
.B(n_5299),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5633),
.Y(n_5869)
);

BUFx3_ASAP7_75t_L g5870 ( 
.A(n_5412),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5567),
.B(n_5188),
.Y(n_5871)
);

AND2x2_ASAP7_75t_L g5872 ( 
.A(n_5589),
.B(n_5215),
.Y(n_5872)
);

AOI21x1_ASAP7_75t_SL g5873 ( 
.A1(n_5632),
.A2(n_5216),
.B(n_5215),
.Y(n_5873)
);

HB1xp67_ASAP7_75t_L g5874 ( 
.A(n_5598),
.Y(n_5874)
);

AND2x2_ASAP7_75t_L g5875 ( 
.A(n_5589),
.B(n_5216),
.Y(n_5875)
);

BUFx3_ASAP7_75t_L g5876 ( 
.A(n_5442),
.Y(n_5876)
);

OA22x2_ASAP7_75t_L g5877 ( 
.A1(n_5728),
.A2(n_5364),
.B1(n_5334),
.B2(n_5229),
.Y(n_5877)
);

AOI21xp5_ASAP7_75t_SL g5878 ( 
.A1(n_5539),
.A2(n_5269),
.B(n_5229),
.Y(n_5878)
);

OAI22xp5_ASAP7_75t_L g5879 ( 
.A1(n_5695),
.A2(n_5286),
.B1(n_5202),
.B2(n_5318),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5463),
.B(n_5269),
.Y(n_5880)
);

HB1xp67_ASAP7_75t_L g5881 ( 
.A(n_5519),
.Y(n_5881)
);

AND2x2_ASAP7_75t_L g5882 ( 
.A(n_5450),
.B(n_5279),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5503),
.Y(n_5883)
);

O2A1O1Ixp5_ASAP7_75t_L g5884 ( 
.A1(n_5608),
.A2(n_5657),
.B(n_5634),
.C(n_5671),
.Y(n_5884)
);

OAI22xp5_ASAP7_75t_L g5885 ( 
.A1(n_5728),
.A2(n_5295),
.B1(n_5333),
.B2(n_5279),
.Y(n_5885)
);

BUFx3_ASAP7_75t_L g5886 ( 
.A(n_5442),
.Y(n_5886)
);

NAND2xp5_ASAP7_75t_L g5887 ( 
.A(n_5645),
.B(n_5081),
.Y(n_5887)
);

INVx4_ASAP7_75t_L g5888 ( 
.A(n_5423),
.Y(n_5888)
);

AND2x2_ASAP7_75t_L g5889 ( 
.A(n_5529),
.B(n_5295),
.Y(n_5889)
);

NOR2xp33_ASAP7_75t_L g5890 ( 
.A(n_5484),
.B(n_142),
.Y(n_5890)
);

AND2x2_ASAP7_75t_L g5891 ( 
.A(n_5692),
.B(n_5319),
.Y(n_5891)
);

NAND2xp5_ASAP7_75t_L g5892 ( 
.A(n_5568),
.B(n_5572),
.Y(n_5892)
);

O2A1O1Ixp33_ASAP7_75t_L g5893 ( 
.A1(n_5708),
.A2(n_5022),
.B(n_5236),
.C(n_5336),
.Y(n_5893)
);

OAI22xp5_ASAP7_75t_L g5894 ( 
.A1(n_5394),
.A2(n_5236),
.B1(n_5319),
.B2(n_5268),
.Y(n_5894)
);

OA21x2_ASAP7_75t_L g5895 ( 
.A1(n_5716),
.A2(n_5164),
.B(n_5081),
.Y(n_5895)
);

AOI21xp5_ASAP7_75t_L g5896 ( 
.A1(n_5417),
.A2(n_5164),
.B(n_5143),
.Y(n_5896)
);

AOI211xp5_ASAP7_75t_L g5897 ( 
.A1(n_5639),
.A2(n_148),
.B(n_142),
.C(n_145),
.Y(n_5897)
);

AND2x2_ASAP7_75t_L g5898 ( 
.A(n_5650),
.B(n_5250),
.Y(n_5898)
);

CKINVDCx5p33_ASAP7_75t_R g5899 ( 
.A(n_5392),
.Y(n_5899)
);

CKINVDCx5p33_ASAP7_75t_R g5900 ( 
.A(n_5410),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5455),
.Y(n_5901)
);

AND2x2_ASAP7_75t_L g5902 ( 
.A(n_5663),
.B(n_5250),
.Y(n_5902)
);

INVxp67_ASAP7_75t_L g5903 ( 
.A(n_5669),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_5496),
.B(n_5249),
.Y(n_5904)
);

AOI21xp5_ASAP7_75t_L g5905 ( 
.A1(n_5574),
.A2(n_5250),
.B(n_2066),
.Y(n_5905)
);

AOI221xp5_ASAP7_75t_L g5906 ( 
.A1(n_5604),
.A2(n_5730),
.B1(n_5706),
.B2(n_5701),
.C(n_5739),
.Y(n_5906)
);

CKINVDCx5p33_ASAP7_75t_R g5907 ( 
.A(n_5466),
.Y(n_5907)
);

HB1xp67_ASAP7_75t_L g5908 ( 
.A(n_5548),
.Y(n_5908)
);

AOI21xp5_ASAP7_75t_SL g5909 ( 
.A1(n_5539),
.A2(n_5394),
.B(n_5735),
.Y(n_5909)
);

BUFx2_ASAP7_75t_L g5910 ( 
.A(n_5715),
.Y(n_5910)
);

AOI21xp5_ASAP7_75t_L g5911 ( 
.A1(n_5574),
.A2(n_2132),
.B(n_2060),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5514),
.Y(n_5912)
);

OR2x2_ASAP7_75t_L g5913 ( 
.A(n_5404),
.B(n_148),
.Y(n_5913)
);

O2A1O1Ixp33_ASAP7_75t_L g5914 ( 
.A1(n_5556),
.A2(n_154),
.B(n_151),
.C(n_152),
.Y(n_5914)
);

O2A1O1Ixp33_ASAP7_75t_L g5915 ( 
.A1(n_5704),
.A2(n_158),
.B(n_152),
.C(n_155),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5688),
.B(n_155),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5524),
.Y(n_5917)
);

AND2x2_ASAP7_75t_L g5918 ( 
.A(n_5693),
.B(n_158),
.Y(n_5918)
);

OAI22xp5_ASAP7_75t_SL g5919 ( 
.A1(n_5441),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_5919)
);

OR2x2_ASAP7_75t_L g5920 ( 
.A(n_5449),
.B(n_159),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5538),
.Y(n_5921)
);

BUFx2_ASAP7_75t_L g5922 ( 
.A(n_5734),
.Y(n_5922)
);

OR2x2_ASAP7_75t_L g5923 ( 
.A(n_5456),
.B(n_162),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5694),
.B(n_163),
.Y(n_5924)
);

OAI22xp5_ASAP7_75t_L g5925 ( 
.A1(n_5609),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5702),
.B(n_165),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5719),
.B(n_166),
.Y(n_5927)
);

AND2x4_ASAP7_75t_L g5928 ( 
.A(n_5649),
.B(n_166),
.Y(n_5928)
);

OAI22xp5_ASAP7_75t_L g5929 ( 
.A1(n_5609),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5541),
.Y(n_5930)
);

OA21x2_ASAP7_75t_L g5931 ( 
.A1(n_5718),
.A2(n_167),
.B(n_169),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5509),
.B(n_171),
.Y(n_5932)
);

CKINVDCx5p33_ASAP7_75t_R g5933 ( 
.A(n_5420),
.Y(n_5933)
);

OA21x2_ASAP7_75t_L g5934 ( 
.A1(n_5721),
.A2(n_171),
.B(n_172),
.Y(n_5934)
);

OR2x2_ASAP7_75t_L g5935 ( 
.A(n_5521),
.B(n_172),
.Y(n_5935)
);

O2A1O1Ixp5_ASAP7_75t_L g5936 ( 
.A1(n_5643),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_5936)
);

CKINVDCx20_ASAP7_75t_R g5937 ( 
.A(n_5424),
.Y(n_5937)
);

AOI21x1_ASAP7_75t_SL g5938 ( 
.A1(n_5531),
.A2(n_174),
.B(n_175),
.Y(n_5938)
);

NOR2xp67_ASAP7_75t_R g5939 ( 
.A(n_5585),
.B(n_177),
.Y(n_5939)
);

O2A1O1Ixp33_ASAP7_75t_L g5940 ( 
.A1(n_5500),
.A2(n_182),
.B(n_178),
.C(n_180),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5738),
.Y(n_5941)
);

OAI22xp5_ASAP7_75t_L g5942 ( 
.A1(n_5639),
.A2(n_184),
.B1(n_180),
.B2(n_183),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5591),
.B(n_184),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5545),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5618),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5547),
.Y(n_5946)
);

AND2x2_ASAP7_75t_SL g5947 ( 
.A(n_5566),
.B(n_185),
.Y(n_5947)
);

OAI22xp5_ASAP7_75t_L g5948 ( 
.A1(n_5661),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5557),
.B(n_186),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5555),
.Y(n_5950)
);

NAND2xp5_ASAP7_75t_L g5951 ( 
.A(n_5576),
.B(n_188),
.Y(n_5951)
);

BUFx2_ASAP7_75t_L g5952 ( 
.A(n_5525),
.Y(n_5952)
);

HB1xp67_ASAP7_75t_L g5953 ( 
.A(n_5621),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5711),
.Y(n_5954)
);

NAND2xp5_ASAP7_75t_L g5955 ( 
.A(n_5714),
.B(n_190),
.Y(n_5955)
);

OAI22xp5_ASAP7_75t_L g5956 ( 
.A1(n_5661),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_5956)
);

O2A1O1Ixp33_ASAP7_75t_L g5957 ( 
.A1(n_5480),
.A2(n_196),
.B(n_191),
.C(n_195),
.Y(n_5957)
);

HB1xp67_ASAP7_75t_L g5958 ( 
.A(n_5649),
.Y(n_5958)
);

AND2x2_ASAP7_75t_L g5959 ( 
.A(n_5517),
.B(n_195),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_SL g5960 ( 
.A(n_5419),
.B(n_1995),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5435),
.B(n_196),
.Y(n_5961)
);

AND2x2_ASAP7_75t_L g5962 ( 
.A(n_5700),
.B(n_197),
.Y(n_5962)
);

AND2x2_ASAP7_75t_L g5963 ( 
.A(n_5550),
.B(n_198),
.Y(n_5963)
);

INVx3_ASAP7_75t_L g5964 ( 
.A(n_5689),
.Y(n_5964)
);

OR2x2_ASAP7_75t_L g5965 ( 
.A(n_5727),
.B(n_199),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5713),
.Y(n_5966)
);

OAI22xp5_ASAP7_75t_L g5967 ( 
.A1(n_5651),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_5967)
);

BUFx2_ASAP7_75t_R g5968 ( 
.A(n_5425),
.Y(n_5968)
);

AND2x4_ASAP7_75t_L g5969 ( 
.A(n_5689),
.B(n_5697),
.Y(n_5969)
);

AND2x2_ASAP7_75t_L g5970 ( 
.A(n_5446),
.B(n_201),
.Y(n_5970)
);

OAI22xp5_ASAP7_75t_L g5971 ( 
.A1(n_5698),
.A2(n_205),
.B1(n_202),
.B2(n_203),
.Y(n_5971)
);

OA21x2_ASAP7_75t_L g5972 ( 
.A1(n_5731),
.A2(n_207),
.B(n_208),
.Y(n_5972)
);

INVx2_ASAP7_75t_L g5973 ( 
.A(n_5736),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5562),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_5537),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5697),
.Y(n_5976)
);

AND2x2_ASAP7_75t_L g5977 ( 
.A(n_5487),
.B(n_207),
.Y(n_5977)
);

NAND2xp5_ASAP7_75t_L g5978 ( 
.A(n_5511),
.B(n_208),
.Y(n_5978)
);

OAI22xp5_ASAP7_75t_L g5979 ( 
.A1(n_5613),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_5979)
);

BUFx2_ASAP7_75t_L g5980 ( 
.A(n_5578),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5569),
.Y(n_5981)
);

O2A1O1Ixp33_ASAP7_75t_L g5982 ( 
.A1(n_5668),
.A2(n_5678),
.B(n_5516),
.C(n_5644),
.Y(n_5982)
);

OR2x2_ASAP7_75t_L g5983 ( 
.A(n_5510),
.B(n_210),
.Y(n_5983)
);

AND2x2_ASAP7_75t_L g5984 ( 
.A(n_5546),
.B(n_212),
.Y(n_5984)
);

OAI22xp5_ASAP7_75t_L g5985 ( 
.A1(n_5687),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_5985)
);

OAI22xp5_ASAP7_75t_L g5986 ( 
.A1(n_5459),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.Y(n_5986)
);

AOI21x1_ASAP7_75t_SL g5987 ( 
.A1(n_5737),
.A2(n_216),
.B(n_217),
.Y(n_5987)
);

AOI21xp5_ASAP7_75t_L g5988 ( 
.A1(n_5459),
.A2(n_2135),
.B(n_2132),
.Y(n_5988)
);

OR2x2_ASAP7_75t_L g5989 ( 
.A(n_5510),
.B(n_217),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5583),
.B(n_218),
.Y(n_5990)
);

OAI22xp5_ASAP7_75t_L g5991 ( 
.A1(n_5451),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_5570),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5453),
.B(n_5615),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5654),
.B(n_221),
.Y(n_5994)
);

AOI21x1_ASAP7_75t_SL g5995 ( 
.A1(n_5508),
.A2(n_222),
.B(n_223),
.Y(n_5995)
);

OAI31xp33_ASAP7_75t_SL g5996 ( 
.A1(n_5428),
.A2(n_227),
.A3(n_223),
.B(n_226),
.Y(n_5996)
);

INVx2_ASAP7_75t_SL g5997 ( 
.A(n_5447),
.Y(n_5997)
);

O2A1O1Ixp33_ASAP7_75t_L g5998 ( 
.A1(n_5444),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_5998)
);

AND2x4_ASAP7_75t_L g5999 ( 
.A(n_5658),
.B(n_228),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_L g6000 ( 
.A(n_5583),
.B(n_229),
.Y(n_6000)
);

BUFx3_ASAP7_75t_L g6001 ( 
.A(n_5423),
.Y(n_6001)
);

OA21x2_ASAP7_75t_L g6002 ( 
.A1(n_5558),
.A2(n_231),
.B(n_233),
.Y(n_6002)
);

AOI21xp5_ASAP7_75t_L g6003 ( 
.A1(n_5416),
.A2(n_2135),
.B(n_2132),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5438),
.B(n_5522),
.Y(n_6004)
);

AOI21xp5_ASAP7_75t_L g6005 ( 
.A1(n_5467),
.A2(n_2135),
.B(n_2132),
.Y(n_6005)
);

CKINVDCx5p33_ASAP7_75t_R g6006 ( 
.A(n_5552),
.Y(n_6006)
);

NAND2xp5_ASAP7_75t_L g6007 ( 
.A(n_5438),
.B(n_231),
.Y(n_6007)
);

O2A1O1Ixp33_ASAP7_75t_L g6008 ( 
.A1(n_5458),
.A2(n_238),
.B(n_235),
.C(n_237),
.Y(n_6008)
);

INVxp67_ASAP7_75t_L g6009 ( 
.A(n_5603),
.Y(n_6009)
);

A2O1A1Ixp33_ASAP7_75t_L g6010 ( 
.A1(n_5451),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_6010)
);

O2A1O1Ixp33_ASAP7_75t_L g6011 ( 
.A1(n_5629),
.A2(n_244),
.B(n_239),
.C(n_241),
.Y(n_6011)
);

O2A1O1Ixp33_ASAP7_75t_L g6012 ( 
.A1(n_5493),
.A2(n_5495),
.B(n_5724),
.C(n_5606),
.Y(n_6012)
);

BUFx6f_ASAP7_75t_L g6013 ( 
.A(n_5560),
.Y(n_6013)
);

HB1xp67_ASAP7_75t_L g6014 ( 
.A(n_5502),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5447),
.B(n_245),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5577),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5452),
.B(n_245),
.Y(n_6017)
);

AOI21xp5_ASAP7_75t_L g6018 ( 
.A1(n_5482),
.A2(n_2144),
.B(n_2135),
.Y(n_6018)
);

AOI21xp5_ASAP7_75t_L g6019 ( 
.A1(n_5474),
.A2(n_2184),
.B(n_2144),
.Y(n_6019)
);

AND2x2_ASAP7_75t_L g6020 ( 
.A(n_5452),
.B(n_246),
.Y(n_6020)
);

AND2x6_ASAP7_75t_L g6021 ( 
.A(n_5457),
.B(n_246),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5586),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5677),
.B(n_5681),
.Y(n_6023)
);

CKINVDCx20_ASAP7_75t_R g6024 ( 
.A(n_5526),
.Y(n_6024)
);

OR2x6_ASAP7_75t_L g6025 ( 
.A(n_5754),
.B(n_5407),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5954),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5743),
.B(n_5429),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5966),
.Y(n_6028)
);

CKINVDCx16_ASAP7_75t_R g6029 ( 
.A(n_5783),
.Y(n_6029)
);

AND2x4_ASAP7_75t_L g6030 ( 
.A(n_5838),
.B(n_5587),
.Y(n_6030)
);

AOI21xp5_ASAP7_75t_SL g6031 ( 
.A1(n_5742),
.A2(n_5426),
.B(n_5414),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5828),
.Y(n_6032)
);

OR2x2_ASAP7_75t_L g6033 ( 
.A(n_5874),
.B(n_5664),
.Y(n_6033)
);

OR2x2_ASAP7_75t_L g6034 ( 
.A(n_5831),
.B(n_5588),
.Y(n_6034)
);

NOR2xp33_ASAP7_75t_R g6035 ( 
.A(n_6024),
.B(n_5933),
.Y(n_6035)
);

INVx2_ASAP7_75t_L g6036 ( 
.A(n_5792),
.Y(n_6036)
);

AO21x2_ASAP7_75t_L g6037 ( 
.A1(n_6004),
.A2(n_5470),
.B(n_5474),
.Y(n_6037)
);

OR2x2_ASAP7_75t_L g6038 ( 
.A(n_5833),
.B(n_5489),
.Y(n_6038)
);

NAND2xp5_ASAP7_75t_L g6039 ( 
.A(n_5839),
.B(n_5472),
.Y(n_6039)
);

OR2x2_ASAP7_75t_L g6040 ( 
.A(n_5800),
.B(n_5489),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5744),
.B(n_5429),
.Y(n_6041)
);

BUFx3_ASAP7_75t_L g6042 ( 
.A(n_5753),
.Y(n_6042)
);

NAND2xp5_ASAP7_75t_L g6043 ( 
.A(n_5762),
.B(n_5540),
.Y(n_6043)
);

AND2x2_ASAP7_75t_L g6044 ( 
.A(n_5787),
.B(n_5691),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5889),
.B(n_5607),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5772),
.B(n_5666),
.Y(n_6046)
);

AND2x2_ASAP7_75t_L g6047 ( 
.A(n_5773),
.B(n_5686),
.Y(n_6047)
);

CKINVDCx16_ASAP7_75t_R g6048 ( 
.A(n_5802),
.Y(n_6048)
);

AND2x4_ASAP7_75t_L g6049 ( 
.A(n_5855),
.B(n_5658),
.Y(n_6049)
);

AND2x4_ASAP7_75t_L g6050 ( 
.A(n_5969),
.B(n_5674),
.Y(n_6050)
);

OR2x2_ASAP7_75t_L g6051 ( 
.A(n_5807),
.B(n_5551),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5973),
.Y(n_6052)
);

NAND2x1p5_ASAP7_75t_L g6053 ( 
.A(n_5779),
.B(n_5585),
.Y(n_6053)
);

INVx1_ASAP7_75t_L g6054 ( 
.A(n_5844),
.Y(n_6054)
);

AND2x4_ASAP7_75t_L g6055 ( 
.A(n_5969),
.B(n_5674),
.Y(n_6055)
);

NOR2xp33_ASAP7_75t_R g6056 ( 
.A(n_5778),
.B(n_5625),
.Y(n_6056)
);

NOR2xp33_ASAP7_75t_R g6057 ( 
.A(n_5900),
.B(n_5699),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5810),
.Y(n_6058)
);

NOR2xp33_ASAP7_75t_R g6059 ( 
.A(n_5937),
.B(n_5720),
.Y(n_6059)
);

OR2x6_ASAP7_75t_L g6060 ( 
.A(n_5805),
.B(n_5407),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5892),
.Y(n_6061)
);

AND2x4_ASAP7_75t_SL g6062 ( 
.A(n_5753),
.B(n_5619),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5892),
.Y(n_6063)
);

AOI22xp33_ASAP7_75t_L g6064 ( 
.A1(n_5853),
.A2(n_5535),
.B1(n_5656),
.B2(n_5579),
.Y(n_6064)
);

AND2x2_ASAP7_75t_L g6065 ( 
.A(n_5857),
.B(n_5686),
.Y(n_6065)
);

CKINVDCx5p33_ASAP7_75t_R g6066 ( 
.A(n_5740),
.Y(n_6066)
);

AND2x2_ASAP7_75t_L g6067 ( 
.A(n_5910),
.B(n_5682),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_5763),
.Y(n_6068)
);

AND2x4_ASAP7_75t_L g6069 ( 
.A(n_5830),
.B(n_5414),
.Y(n_6069)
);

CKINVDCx8_ASAP7_75t_R g6070 ( 
.A(n_5753),
.Y(n_6070)
);

CKINVDCx16_ASAP7_75t_R g6071 ( 
.A(n_6023),
.Y(n_6071)
);

BUFx6f_ASAP7_75t_L g6072 ( 
.A(n_5876),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5791),
.Y(n_6073)
);

INVxp67_ASAP7_75t_L g6074 ( 
.A(n_5766),
.Y(n_6074)
);

CKINVDCx16_ASAP7_75t_R g6075 ( 
.A(n_6013),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5794),
.Y(n_6076)
);

CKINVDCx16_ASAP7_75t_R g6077 ( 
.A(n_6013),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5782),
.B(n_5461),
.Y(n_6078)
);

O2A1O1Ixp33_ASAP7_75t_L g6079 ( 
.A1(n_5745),
.A2(n_5735),
.B(n_5679),
.C(n_5544),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_5841),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_5922),
.B(n_5582),
.Y(n_6081)
);

INVx5_ASAP7_75t_L g6082 ( 
.A(n_6021),
.Y(n_6082)
);

OR2x2_ASAP7_75t_L g6083 ( 
.A(n_5864),
.B(n_5551),
.Y(n_6083)
);

INVx1_ASAP7_75t_SL g6084 ( 
.A(n_5968),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_5793),
.B(n_5725),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5824),
.Y(n_6086)
);

OR2x2_ASAP7_75t_L g6087 ( 
.A(n_5834),
.B(n_5551),
.Y(n_6087)
);

CKINVDCx5p33_ASAP7_75t_R g6088 ( 
.A(n_5907),
.Y(n_6088)
);

OR2x6_ASAP7_75t_L g6089 ( 
.A(n_5795),
.B(n_5407),
.Y(n_6089)
);

AND2x2_ASAP7_75t_L g6090 ( 
.A(n_5861),
.B(n_5582),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_5871),
.B(n_5675),
.Y(n_6091)
);

INVx3_ASAP7_75t_L g6092 ( 
.A(n_5888),
.Y(n_6092)
);

AND2x4_ASAP7_75t_L g6093 ( 
.A(n_5830),
.B(n_5426),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5759),
.B(n_5725),
.Y(n_6094)
);

AOI22xp33_ASAP7_75t_SL g6095 ( 
.A1(n_5745),
.A2(n_5441),
.B1(n_5624),
.B2(n_5585),
.Y(n_6095)
);

OR2x2_ASAP7_75t_L g6096 ( 
.A(n_5836),
.B(n_5533),
.Y(n_6096)
);

AND2x4_ASAP7_75t_L g6097 ( 
.A(n_5770),
.B(n_5431),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5824),
.Y(n_6098)
);

NAND2xp33_ASAP7_75t_R g6099 ( 
.A(n_5952),
.B(n_247),
.Y(n_6099)
);

AO31x2_ASAP7_75t_L g6100 ( 
.A1(n_6004),
.A2(n_5473),
.A3(n_5431),
.B(n_5631),
.Y(n_6100)
);

NAND2xp33_ASAP7_75t_R g6101 ( 
.A(n_5975),
.B(n_247),
.Y(n_6101)
);

HB1xp67_ASAP7_75t_L g6102 ( 
.A(n_5881),
.Y(n_6102)
);

CKINVDCx20_ASAP7_75t_R g6103 ( 
.A(n_5750),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5796),
.Y(n_6104)
);

OR2x6_ASAP7_75t_L g6105 ( 
.A(n_5909),
.B(n_5473),
.Y(n_6105)
);

OR2x6_ASAP7_75t_L g6106 ( 
.A(n_5878),
.B(n_5469),
.Y(n_6106)
);

CKINVDCx20_ASAP7_75t_R g6107 ( 
.A(n_5899),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_5811),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5872),
.B(n_5675),
.Y(n_6109)
);

CKINVDCx5p33_ASAP7_75t_R g6110 ( 
.A(n_6006),
.Y(n_6110)
);

OAI21x1_ASAP7_75t_L g6111 ( 
.A1(n_5868),
.A2(n_5846),
.B(n_5840),
.Y(n_6111)
);

NOR2xp33_ASAP7_75t_L g6112 ( 
.A(n_5888),
.B(n_5476),
.Y(n_6112)
);

CKINVDCx16_ASAP7_75t_R g6113 ( 
.A(n_6013),
.Y(n_6113)
);

NOR2x1_ASAP7_75t_SL g6114 ( 
.A(n_5765),
.B(n_5624),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5875),
.B(n_5710),
.Y(n_6115)
);

OR2x2_ASAP7_75t_L g6116 ( 
.A(n_5868),
.B(n_5533),
.Y(n_6116)
);

AOI22xp5_ASAP7_75t_L g6117 ( 
.A1(n_5986),
.A2(n_5523),
.B1(n_5469),
.B2(n_5672),
.Y(n_6117)
);

INVx2_ASAP7_75t_L g6118 ( 
.A(n_5976),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5845),
.Y(n_6119)
);

AND2x2_ASAP7_75t_L g6120 ( 
.A(n_5820),
.B(n_5710),
.Y(n_6120)
);

AOI22xp5_ASAP7_75t_L g6121 ( 
.A1(n_5986),
.A2(n_5523),
.B1(n_5670),
.B2(n_5573),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_5814),
.B(n_5470),
.Y(n_6122)
);

INVxp67_ASAP7_75t_L g6123 ( 
.A(n_5939),
.Y(n_6123)
);

NOR2xp33_ASAP7_75t_R g6124 ( 
.A(n_5947),
.B(n_5603),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_5780),
.B(n_5533),
.Y(n_6125)
);

INVx2_ASAP7_75t_L g6126 ( 
.A(n_5958),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_5850),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5964),
.Y(n_6128)
);

INVx2_ASAP7_75t_L g6129 ( 
.A(n_5964),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_5974),
.Y(n_6130)
);

INVxp67_ASAP7_75t_L g6131 ( 
.A(n_5939),
.Y(n_6131)
);

AND2x2_ASAP7_75t_L g6132 ( 
.A(n_5785),
.B(n_5638),
.Y(n_6132)
);

INVxp67_ASAP7_75t_L g6133 ( 
.A(n_5955),
.Y(n_6133)
);

AND2x2_ASAP7_75t_L g6134 ( 
.A(n_5788),
.B(n_5638),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_5886),
.Y(n_6135)
);

NAND2xp33_ASAP7_75t_R g6136 ( 
.A(n_5962),
.B(n_248),
.Y(n_6136)
);

BUFx2_ASAP7_75t_L g6137 ( 
.A(n_6001),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_5870),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_5803),
.B(n_5561),
.Y(n_6139)
);

NOR2xp33_ASAP7_75t_R g6140 ( 
.A(n_6021),
.B(n_5584),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_L g6141 ( 
.A(n_5803),
.B(n_5816),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5859),
.Y(n_6142)
);

INVx2_ASAP7_75t_L g6143 ( 
.A(n_5827),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_5817),
.B(n_5760),
.Y(n_6144)
);

OAI21xp5_ASAP7_75t_SL g6145 ( 
.A1(n_5996),
.A2(n_5906),
.B(n_5769),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5883),
.Y(n_6146)
);

NAND3xp33_ASAP7_75t_SL g6147 ( 
.A(n_5819),
.B(n_5741),
.C(n_5897),
.Y(n_6147)
);

INVx1_ASAP7_75t_SL g6148 ( 
.A(n_5816),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_5757),
.B(n_5543),
.Y(n_6149)
);

HB1xp67_ASAP7_75t_L g6150 ( 
.A(n_5767),
.Y(n_6150)
);

CKINVDCx5p33_ASAP7_75t_R g6151 ( 
.A(n_5867),
.Y(n_6151)
);

NAND3xp33_ASAP7_75t_L g6152 ( 
.A(n_5996),
.B(n_5602),
.C(n_5676),
.Y(n_6152)
);

INVx2_ASAP7_75t_SL g6153 ( 
.A(n_5768),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_5912),
.Y(n_6154)
);

O2A1O1Ixp33_ASAP7_75t_SL g6155 ( 
.A1(n_5848),
.A2(n_5584),
.B(n_5605),
.C(n_5624),
.Y(n_6155)
);

CKINVDCx16_ASAP7_75t_R g6156 ( 
.A(n_5994),
.Y(n_6156)
);

BUFx6f_ASAP7_75t_L g6157 ( 
.A(n_5768),
.Y(n_6157)
);

OR2x6_ASAP7_75t_L g6158 ( 
.A(n_5842),
.B(n_5457),
.Y(n_6158)
);

OR2x6_ASAP7_75t_L g6159 ( 
.A(n_5768),
.B(n_5457),
.Y(n_6159)
);

OR2x2_ASAP7_75t_L g6160 ( 
.A(n_5887),
.B(n_5561),
.Y(n_6160)
);

A2O1A1Ixp33_ASAP7_75t_L g6161 ( 
.A1(n_5915),
.A2(n_5637),
.B(n_5512),
.C(n_5536),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5826),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_5826),
.Y(n_6163)
);

OAI21x1_ASAP7_75t_L g6164 ( 
.A1(n_5747),
.A2(n_5679),
.B(n_5592),
.Y(n_6164)
);

CKINVDCx5p33_ASAP7_75t_R g6165 ( 
.A(n_5980),
.Y(n_6165)
);

AND2x2_ASAP7_75t_L g6166 ( 
.A(n_5882),
.B(n_5543),
.Y(n_6166)
);

CKINVDCx5p33_ASAP7_75t_R g6167 ( 
.A(n_5786),
.Y(n_6167)
);

OR2x6_ASAP7_75t_L g6168 ( 
.A(n_5786),
.B(n_5993),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_5856),
.B(n_5600),
.Y(n_6169)
);

NOR2xp33_ASAP7_75t_R g6170 ( 
.A(n_6021),
.B(n_5605),
.Y(n_6170)
);

INVx3_ASAP7_75t_L g6171 ( 
.A(n_5786),
.Y(n_6171)
);

CKINVDCx5p33_ASAP7_75t_R g6172 ( 
.A(n_5849),
.Y(n_6172)
);

NOR3xp33_ASAP7_75t_SL g6173 ( 
.A(n_5919),
.B(n_5640),
.C(n_5512),
.Y(n_6173)
);

NOR2xp33_ASAP7_75t_R g6174 ( 
.A(n_6021),
.B(n_5512),
.Y(n_6174)
);

AND2x2_ASAP7_75t_L g6175 ( 
.A(n_5775),
.B(n_5600),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5775),
.B(n_5610),
.Y(n_6176)
);

INVx2_ASAP7_75t_L g6177 ( 
.A(n_5869),
.Y(n_6177)
);

NAND2xp5_ASAP7_75t_L g6178 ( 
.A(n_5849),
.B(n_5561),
.Y(n_6178)
);

OA21x2_ASAP7_75t_L g6179 ( 
.A1(n_5747),
.A2(n_5581),
.B(n_5571),
.Y(n_6179)
);

CKINVDCx20_ASAP7_75t_R g6180 ( 
.A(n_6009),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_5997),
.Y(n_6181)
);

AO21x2_ASAP7_75t_L g6182 ( 
.A1(n_5990),
.A2(n_6000),
.B(n_6007),
.Y(n_6182)
);

CKINVDCx16_ASAP7_75t_R g6183 ( 
.A(n_5984),
.Y(n_6183)
);

OR2x2_ASAP7_75t_L g6184 ( 
.A(n_5953),
.B(n_5563),
.Y(n_6184)
);

NAND2xp33_ASAP7_75t_SL g6185 ( 
.A(n_5999),
.B(n_5563),
.Y(n_6185)
);

AND2x2_ASAP7_75t_SL g6186 ( 
.A(n_6007),
.B(n_5563),
.Y(n_6186)
);

NOR2xp33_ASAP7_75t_L g6187 ( 
.A(n_5752),
.B(n_5610),
.Y(n_6187)
);

OR2x6_ASAP7_75t_L g6188 ( 
.A(n_5808),
.B(n_5626),
.Y(n_6188)
);

AND2x2_ASAP7_75t_L g6189 ( 
.A(n_5764),
.B(n_5626),
.Y(n_6189)
);

NOR2xp33_ASAP7_75t_R g6190 ( 
.A(n_5890),
.B(n_6015),
.Y(n_6190)
);

AO31x2_ASAP7_75t_L g6191 ( 
.A1(n_5801),
.A2(n_5637),
.A3(n_5667),
.B(n_5652),
.Y(n_6191)
);

CKINVDCx5p33_ASAP7_75t_R g6192 ( 
.A(n_6014),
.Y(n_6192)
);

INVx2_ASAP7_75t_L g6193 ( 
.A(n_5815),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_5917),
.Y(n_6194)
);

INVx2_ASAP7_75t_L g6195 ( 
.A(n_5901),
.Y(n_6195)
);

INVx3_ASAP7_75t_L g6196 ( 
.A(n_5799),
.Y(n_6196)
);

NAND2xp33_ASAP7_75t_R g6197 ( 
.A(n_5999),
.B(n_250),
.Y(n_6197)
);

OAI22xp5_ASAP7_75t_L g6198 ( 
.A1(n_6010),
.A2(n_5637),
.B1(n_5690),
.B2(n_5680),
.Y(n_6198)
);

NAND2xp5_ASAP7_75t_L g6199 ( 
.A(n_5903),
.B(n_5921),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_5981),
.B(n_5652),
.Y(n_6200)
);

NAND2xp33_ASAP7_75t_SL g6201 ( 
.A(n_5769),
.B(n_5565),
.Y(n_6201)
);

CKINVDCx16_ASAP7_75t_R g6202 ( 
.A(n_5880),
.Y(n_6202)
);

NAND2xp5_ASAP7_75t_L g6203 ( 
.A(n_5930),
.B(n_5944),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_L g6204 ( 
.A(n_5946),
.B(n_5565),
.Y(n_6204)
);

NAND2xp33_ASAP7_75t_SL g6205 ( 
.A(n_5928),
.B(n_5565),
.Y(n_6205)
);

BUFx3_ASAP7_75t_L g6206 ( 
.A(n_6022),
.Y(n_6206)
);

BUFx6f_ASAP7_75t_L g6207 ( 
.A(n_5928),
.Y(n_6207)
);

OR2x6_ASAP7_75t_L g6208 ( 
.A(n_5860),
.B(n_5667),
.Y(n_6208)
);

INVxp67_ASAP7_75t_L g6209 ( 
.A(n_5955),
.Y(n_6209)
);

NAND2xp5_ASAP7_75t_L g6210 ( 
.A(n_5950),
.B(n_5594),
.Y(n_6210)
);

AND2x4_ASAP7_75t_L g6211 ( 
.A(n_5770),
.B(n_5594),
.Y(n_6211)
);

CKINVDCx5p33_ASAP7_75t_R g6212 ( 
.A(n_6017),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_5806),
.Y(n_6213)
);

A2O1A1Ixp33_ASAP7_75t_L g6214 ( 
.A1(n_5771),
.A2(n_5498),
.B(n_5623),
.C(n_5722),
.Y(n_6214)
);

AOI22xp33_ASAP7_75t_L g6215 ( 
.A1(n_5877),
.A2(n_5497),
.B1(n_5532),
.B2(n_5520),
.Y(n_6215)
);

OR2x2_ASAP7_75t_L g6216 ( 
.A(n_5790),
.B(n_5594),
.Y(n_6216)
);

AND3x1_ASAP7_75t_L g6217 ( 
.A(n_6020),
.B(n_5655),
.C(n_5647),
.Y(n_6217)
);

INVxp67_ASAP7_75t_L g6218 ( 
.A(n_5983),
.Y(n_6218)
);

INVx2_ASAP7_75t_L g6219 ( 
.A(n_5941),
.Y(n_6219)
);

NAND2xp5_ASAP7_75t_L g6220 ( 
.A(n_5990),
.B(n_5597),
.Y(n_6220)
);

OAI22xp5_ASAP7_75t_SL g6221 ( 
.A1(n_5749),
.A2(n_5597),
.B1(n_5660),
.B2(n_5642),
.Y(n_6221)
);

AND2x2_ASAP7_75t_L g6222 ( 
.A(n_5799),
.B(n_5597),
.Y(n_6222)
);

NAND2x1p5_ASAP7_75t_L g6223 ( 
.A(n_5862),
.B(n_5829),
.Y(n_6223)
);

AO31x2_ASAP7_75t_L g6224 ( 
.A1(n_6000),
.A2(n_5822),
.A3(n_5756),
.B(n_5818),
.Y(n_6224)
);

OR2x2_ASAP7_75t_SL g6225 ( 
.A(n_5989),
.B(n_251),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_5862),
.Y(n_6226)
);

AND3x2_ASAP7_75t_L g6227 ( 
.A(n_5963),
.B(n_253),
.C(n_254),
.Y(n_6227)
);

HB1xp67_ASAP7_75t_L g6228 ( 
.A(n_5812),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_5945),
.Y(n_6229)
);

OR2x6_ASAP7_75t_L g6230 ( 
.A(n_5877),
.B(n_5505),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5813),
.Y(n_6231)
);

OR2x2_ASAP7_75t_L g6232 ( 
.A(n_5781),
.B(n_5599),
.Y(n_6232)
);

INVx2_ASAP7_75t_L g6233 ( 
.A(n_5748),
.Y(n_6233)
);

NOR2xp33_ASAP7_75t_R g6234 ( 
.A(n_5961),
.B(n_253),
.Y(n_6234)
);

AND2x2_ASAP7_75t_L g6235 ( 
.A(n_5992),
.B(n_5595),
.Y(n_6235)
);

OAI22xp5_ASAP7_75t_SL g6236 ( 
.A1(n_5749),
.A2(n_5991),
.B1(n_5948),
.B2(n_5956),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_5908),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_5932),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6016),
.B(n_5593),
.Y(n_6239)
);

NAND3xp33_ASAP7_75t_SL g6240 ( 
.A(n_5797),
.B(n_5549),
.C(n_5732),
.Y(n_6240)
);

CKINVDCx5p33_ASAP7_75t_R g6241 ( 
.A(n_5970),
.Y(n_6241)
);

NAND2xp33_ASAP7_75t_R g6242 ( 
.A(n_5931),
.B(n_255),
.Y(n_6242)
);

NOR2x1p5_ASAP7_75t_L g6243 ( 
.A(n_5978),
.B(n_5949),
.Y(n_6243)
);

NAND2xp5_ASAP7_75t_L g6244 ( 
.A(n_5982),
.B(n_5527),
.Y(n_6244)
);

AND2x2_ASAP7_75t_L g6245 ( 
.A(n_5854),
.B(n_5534),
.Y(n_6245)
);

AND2x4_ASAP7_75t_SL g6246 ( 
.A(n_5891),
.B(n_5733),
.Y(n_6246)
);

CKINVDCx5p33_ASAP7_75t_R g6247 ( 
.A(n_5959),
.Y(n_6247)
);

NAND2xp5_ASAP7_75t_L g6248 ( 
.A(n_5784),
.B(n_5528),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_5932),
.Y(n_6249)
);

CKINVDCx20_ASAP7_75t_R g6250 ( 
.A(n_5977),
.Y(n_6250)
);

AOI22xp33_ASAP7_75t_L g6251 ( 
.A1(n_5991),
.A2(n_5729),
.B1(n_2426),
.B2(n_2428),
.Y(n_6251)
);

AND2x2_ASAP7_75t_L g6252 ( 
.A(n_5748),
.B(n_256),
.Y(n_6252)
);

BUFx10_ASAP7_75t_L g6253 ( 
.A(n_5995),
.Y(n_6253)
);

INVx3_ASAP7_75t_L g6254 ( 
.A(n_5913),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_5965),
.Y(n_6255)
);

INVx2_ASAP7_75t_L g6256 ( 
.A(n_5935),
.Y(n_6256)
);

NAND2xp33_ASAP7_75t_R g6257 ( 
.A(n_5931),
.B(n_256),
.Y(n_6257)
);

HB1xp67_ASAP7_75t_L g6258 ( 
.A(n_5902),
.Y(n_6258)
);

HB1xp67_ASAP7_75t_L g6259 ( 
.A(n_5898),
.Y(n_6259)
);

AOI22xp33_ASAP7_75t_L g6260 ( 
.A1(n_5896),
.A2(n_2426),
.B1(n_2428),
.B2(n_2398),
.Y(n_6260)
);

BUFx6f_ASAP7_75t_L g6261 ( 
.A(n_5920),
.Y(n_6261)
);

HB1xp67_ASAP7_75t_L g6262 ( 
.A(n_5934),
.Y(n_6262)
);

CKINVDCx5p33_ASAP7_75t_R g6263 ( 
.A(n_5916),
.Y(n_6263)
);

AOI22xp33_ASAP7_75t_L g6264 ( 
.A1(n_5942),
.A2(n_2428),
.B1(n_2432),
.B2(n_2426),
.Y(n_6264)
);

BUFx2_ASAP7_75t_L g6265 ( 
.A(n_5923),
.Y(n_6265)
);

OAI21xp5_ASAP7_75t_L g6266 ( 
.A1(n_5957),
.A2(n_257),
.B(n_260),
.Y(n_6266)
);

CKINVDCx16_ASAP7_75t_R g6267 ( 
.A(n_5979),
.Y(n_6267)
);

NOR2xp33_ASAP7_75t_R g6268 ( 
.A(n_5918),
.B(n_260),
.Y(n_6268)
);

OAI21xp5_ASAP7_75t_SL g6269 ( 
.A1(n_5940),
.A2(n_261),
.B(n_262),
.Y(n_6269)
);

INVx2_ASAP7_75t_L g6270 ( 
.A(n_5943),
.Y(n_6270)
);

HB1xp67_ASAP7_75t_L g6271 ( 
.A(n_5934),
.Y(n_6271)
);

CKINVDCx16_ASAP7_75t_R g6272 ( 
.A(n_5979),
.Y(n_6272)
);

A2O1A1Ixp33_ASAP7_75t_L g6273 ( 
.A1(n_5771),
.A2(n_264),
.B(n_261),
.C(n_263),
.Y(n_6273)
);

OR2x2_ASAP7_75t_L g6274 ( 
.A(n_5904),
.B(n_5949),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5972),
.Y(n_6275)
);

NOR2xp33_ASAP7_75t_R g6276 ( 
.A(n_5924),
.B(n_263),
.Y(n_6276)
);

AND2x2_ASAP7_75t_L g6277 ( 
.A(n_5823),
.B(n_264),
.Y(n_6277)
);

AOI22xp33_ASAP7_75t_SL g6278 ( 
.A1(n_6267),
.A2(n_5948),
.B1(n_5956),
.B2(n_5942),
.Y(n_6278)
);

NAND2xp5_ASAP7_75t_L g6279 ( 
.A(n_6182),
.B(n_5755),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_6026),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6026),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_6261),
.Y(n_6282)
);

INVx2_ASAP7_75t_L g6283 ( 
.A(n_6160),
.Y(n_6283)
);

OA21x2_ASAP7_75t_L g6284 ( 
.A1(n_6275),
.A2(n_5858),
.B(n_5746),
.Y(n_6284)
);

OR2x2_ASAP7_75t_L g6285 ( 
.A(n_6122),
.B(n_5951),
.Y(n_6285)
);

AND2x4_ASAP7_75t_L g6286 ( 
.A(n_6092),
.B(n_5865),
.Y(n_6286)
);

NAND2xp5_ASAP7_75t_L g6287 ( 
.A(n_6262),
.B(n_5972),
.Y(n_6287)
);

OAI211xp5_ASAP7_75t_L g6288 ( 
.A1(n_6145),
.A2(n_5761),
.B(n_5998),
.C(n_6008),
.Y(n_6288)
);

AND2x2_ASAP7_75t_L g6289 ( 
.A(n_6050),
.B(n_6055),
.Y(n_6289)
);

OR2x2_ASAP7_75t_L g6290 ( 
.A(n_6116),
.B(n_6232),
.Y(n_6290)
);

OR2x6_ASAP7_75t_L g6291 ( 
.A(n_6025),
.B(n_5835),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6028),
.Y(n_6292)
);

OA21x2_ASAP7_75t_L g6293 ( 
.A1(n_6275),
.A2(n_5809),
.B(n_5951),
.Y(n_6293)
);

NOR2xp33_ASAP7_75t_L g6294 ( 
.A(n_6272),
.B(n_5925),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6050),
.B(n_5926),
.Y(n_6295)
);

OAI21xp5_ASAP7_75t_L g6296 ( 
.A1(n_6147),
.A2(n_5884),
.B(n_5936),
.Y(n_6296)
);

OR2x6_ASAP7_75t_L g6297 ( 
.A(n_6025),
.B(n_5789),
.Y(n_6297)
);

HB1xp67_ASAP7_75t_L g6298 ( 
.A(n_6271),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6028),
.Y(n_6299)
);

INVx4_ASAP7_75t_L g6300 ( 
.A(n_6072),
.Y(n_6300)
);

OA21x2_ASAP7_75t_L g6301 ( 
.A1(n_6248),
.A2(n_5852),
.B(n_5904),
.Y(n_6301)
);

AOI221xp5_ASAP7_75t_L g6302 ( 
.A1(n_6236),
.A2(n_5925),
.B1(n_5929),
.B2(n_5777),
.C(n_5967),
.Y(n_6302)
);

OR2x2_ASAP7_75t_L g6303 ( 
.A(n_6078),
.B(n_6002),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_6068),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6073),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_6261),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_6261),
.Y(n_6307)
);

NAND4xp25_ASAP7_75t_L g6308 ( 
.A(n_6273),
.B(n_5777),
.C(n_5914),
.D(n_5929),
.Y(n_6308)
);

OR2x2_ASAP7_75t_L g6309 ( 
.A(n_6037),
.B(n_6002),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6076),
.Y(n_6310)
);

INVx2_ASAP7_75t_SL g6311 ( 
.A(n_6062),
.Y(n_6311)
);

INVx2_ASAP7_75t_L g6312 ( 
.A(n_6184),
.Y(n_6312)
);

AND2x2_ASAP7_75t_L g6313 ( 
.A(n_6055),
.B(n_5927),
.Y(n_6313)
);

OAI211xp5_ASAP7_75t_SL g6314 ( 
.A1(n_6244),
.A2(n_6012),
.B(n_5971),
.C(n_5967),
.Y(n_6314)
);

AO21x2_ASAP7_75t_L g6315 ( 
.A1(n_6114),
.A2(n_5832),
.B(n_5905),
.Y(n_6315)
);

NOR2xp33_ASAP7_75t_L g6316 ( 
.A(n_6071),
.B(n_5971),
.Y(n_6316)
);

BUFx2_ASAP7_75t_L g6317 ( 
.A(n_6168),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6104),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_6202),
.B(n_5885),
.Y(n_6319)
);

AO21x2_ASAP7_75t_L g6320 ( 
.A1(n_6114),
.A2(n_5985),
.B(n_5804),
.Y(n_6320)
);

OA21x2_ASAP7_75t_L g6321 ( 
.A1(n_6123),
.A2(n_5988),
.B(n_6019),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_6069),
.B(n_5885),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_6102),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_6233),
.Y(n_6324)
);

OA21x2_ASAP7_75t_L g6325 ( 
.A1(n_6131),
.A2(n_5960),
.B(n_5894),
.Y(n_6325)
);

OAI322xp33_ASAP7_75t_L g6326 ( 
.A1(n_6242),
.A2(n_5985),
.A3(n_5863),
.B1(n_5804),
.B2(n_5774),
.C1(n_5894),
.C2(n_6011),
.Y(n_6326)
);

AO21x2_ASAP7_75t_L g6327 ( 
.A1(n_6031),
.A2(n_5774),
.B(n_5863),
.Y(n_6327)
);

OR2x2_ASAP7_75t_L g6328 ( 
.A(n_6274),
.B(n_5895),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_SL g6329 ( 
.A(n_6095),
.B(n_5847),
.Y(n_6329)
);

AOI22xp33_ASAP7_75t_L g6330 ( 
.A1(n_6266),
.A2(n_5847),
.B1(n_5879),
.B2(n_5895),
.Y(n_6330)
);

BUFx3_ASAP7_75t_L g6331 ( 
.A(n_6070),
.Y(n_6331)
);

AO21x2_ASAP7_75t_L g6332 ( 
.A1(n_6277),
.A2(n_6018),
.B(n_6003),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_6108),
.Y(n_6333)
);

AOI21xp5_ASAP7_75t_SL g6334 ( 
.A1(n_6089),
.A2(n_5866),
.B(n_5893),
.Y(n_6334)
);

INVx2_ASAP7_75t_L g6335 ( 
.A(n_6223),
.Y(n_6335)
);

OAI21xp5_ASAP7_75t_L g6336 ( 
.A1(n_6161),
.A2(n_5879),
.B(n_5987),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6040),
.Y(n_6337)
);

OA21x2_ASAP7_75t_L g6338 ( 
.A1(n_6111),
.A2(n_6005),
.B(n_5911),
.Y(n_6338)
);

AND2x4_ASAP7_75t_L g6339 ( 
.A(n_6092),
.B(n_5873),
.Y(n_6339)
);

AND2x2_ASAP7_75t_L g6340 ( 
.A(n_6069),
.B(n_5798),
.Y(n_6340)
);

INVx2_ASAP7_75t_L g6341 ( 
.A(n_6083),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_6119),
.Y(n_6342)
);

HB1xp67_ASAP7_75t_L g6343 ( 
.A(n_6150),
.Y(n_6343)
);

BUFx6f_ASAP7_75t_L g6344 ( 
.A(n_6072),
.Y(n_6344)
);

AO21x2_ASAP7_75t_L g6345 ( 
.A1(n_6234),
.A2(n_5751),
.B(n_5758),
.Y(n_6345)
);

AND2x2_ASAP7_75t_L g6346 ( 
.A(n_6093),
.B(n_5798),
.Y(n_6346)
);

OR2x6_ASAP7_75t_L g6347 ( 
.A(n_6060),
.B(n_5821),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_6127),
.Y(n_6348)
);

INVx4_ASAP7_75t_L g6349 ( 
.A(n_6072),
.Y(n_6349)
);

AND2x2_ASAP7_75t_L g6350 ( 
.A(n_6093),
.B(n_5837),
.Y(n_6350)
);

OR2x2_ASAP7_75t_SL g6351 ( 
.A(n_6029),
.B(n_5776),
.Y(n_6351)
);

OAI21x1_ASAP7_75t_L g6352 ( 
.A1(n_6196),
.A2(n_5837),
.B(n_5843),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6118),
.Y(n_6353)
);

HB1xp67_ASAP7_75t_L g6354 ( 
.A(n_6228),
.Y(n_6354)
);

INVx2_ASAP7_75t_L g6355 ( 
.A(n_6126),
.Y(n_6355)
);

OA21x2_ASAP7_75t_L g6356 ( 
.A1(n_6215),
.A2(n_5843),
.B(n_5938),
.Y(n_6356)
);

INVx1_ASAP7_75t_L g6357 ( 
.A(n_6142),
.Y(n_6357)
);

AND2x2_ASAP7_75t_L g6358 ( 
.A(n_6222),
.B(n_5825),
.Y(n_6358)
);

OAI22xp33_ASAP7_75t_L g6359 ( 
.A1(n_6230),
.A2(n_6099),
.B1(n_6257),
.B2(n_6269),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6245),
.B(n_5825),
.Y(n_6360)
);

INVx4_ASAP7_75t_L g6361 ( 
.A(n_6075),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_6047),
.B(n_5851),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6053),
.B(n_5851),
.Y(n_6363)
);

HB1xp67_ASAP7_75t_L g6364 ( 
.A(n_6086),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6146),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6154),
.Y(n_6366)
);

BUFx6f_ASAP7_75t_L g6367 ( 
.A(n_6042),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6087),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_6194),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6203),
.Y(n_6370)
);

AND2x2_ASAP7_75t_L g6371 ( 
.A(n_6196),
.B(n_265),
.Y(n_6371)
);

OR2x2_ASAP7_75t_L g6372 ( 
.A(n_6039),
.B(n_265),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_6254),
.Y(n_6373)
);

BUFx3_ASAP7_75t_L g6374 ( 
.A(n_6168),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_6254),
.Y(n_6375)
);

OR2x6_ASAP7_75t_L g6376 ( 
.A(n_6060),
.B(n_267),
.Y(n_6376)
);

INVx2_ASAP7_75t_L g6377 ( 
.A(n_6128),
.Y(n_6377)
);

CKINVDCx5p33_ASAP7_75t_R g6378 ( 
.A(n_6066),
.Y(n_6378)
);

NOR2xp33_ASAP7_75t_L g6379 ( 
.A(n_6077),
.B(n_267),
.Y(n_6379)
);

AND2x2_ASAP7_75t_L g6380 ( 
.A(n_6097),
.B(n_268),
.Y(n_6380)
);

AO21x2_ASAP7_75t_L g6381 ( 
.A1(n_6124),
.A2(n_269),
.B(n_270),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6199),
.Y(n_6382)
);

OAI21xp5_ASAP7_75t_L g6383 ( 
.A1(n_6201),
.A2(n_273),
.B(n_274),
.Y(n_6383)
);

OAI31xp33_ASAP7_75t_L g6384 ( 
.A1(n_6155),
.A2(n_275),
.A3(n_273),
.B(n_274),
.Y(n_6384)
);

NAND2xp5_ASAP7_75t_L g6385 ( 
.A(n_6061),
.B(n_275),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_6097),
.B(n_276),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6054),
.Y(n_6387)
);

HB1xp67_ASAP7_75t_L g6388 ( 
.A(n_6086),
.Y(n_6388)
);

OA21x2_ASAP7_75t_L g6389 ( 
.A1(n_6164),
.A2(n_276),
.B(n_280),
.Y(n_6389)
);

AO21x2_ASAP7_75t_L g6390 ( 
.A1(n_6141),
.A2(n_281),
.B(n_283),
.Y(n_6390)
);

OA21x2_ASAP7_75t_L g6391 ( 
.A1(n_6098),
.A2(n_283),
.B(n_285),
.Y(n_6391)
);

OAI21x1_ASAP7_75t_L g6392 ( 
.A1(n_6129),
.A2(n_285),
.B(n_286),
.Y(n_6392)
);

INVxp67_ASAP7_75t_SL g6393 ( 
.A(n_6133),
.Y(n_6393)
);

AO21x2_ASAP7_75t_L g6394 ( 
.A1(n_6098),
.A2(n_6163),
.B(n_6162),
.Y(n_6394)
);

INVx3_ASAP7_75t_L g6395 ( 
.A(n_6157),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_6137),
.Y(n_6396)
);

NOR2xp67_ASAP7_75t_SL g6397 ( 
.A(n_6082),
.B(n_286),
.Y(n_6397)
);

OR2x2_ASAP7_75t_L g6398 ( 
.A(n_6265),
.B(n_287),
.Y(n_6398)
);

INVx2_ASAP7_75t_L g6399 ( 
.A(n_6216),
.Y(n_6399)
);

NAND3xp33_ASAP7_75t_L g6400 ( 
.A(n_6230),
.B(n_288),
.C(n_289),
.Y(n_6400)
);

HB1xp67_ASAP7_75t_L g6401 ( 
.A(n_6162),
.Y(n_6401)
);

INVx2_ASAP7_75t_L g6402 ( 
.A(n_6207),
.Y(n_6402)
);

AOI21xp5_ASAP7_75t_SL g6403 ( 
.A1(n_6089),
.A2(n_290),
.B(n_291),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6052),
.Y(n_6404)
);

INVx2_ASAP7_75t_SL g6405 ( 
.A(n_6113),
.Y(n_6405)
);

OR2x2_ASAP7_75t_L g6406 ( 
.A(n_6074),
.B(n_290),
.Y(n_6406)
);

OR2x6_ASAP7_75t_L g6407 ( 
.A(n_6105),
.B(n_292),
.Y(n_6407)
);

OA21x2_ASAP7_75t_L g6408 ( 
.A1(n_6163),
.A2(n_292),
.B(n_293),
.Y(n_6408)
);

INVx2_ASAP7_75t_L g6409 ( 
.A(n_6207),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6063),
.Y(n_6410)
);

OAI221xp5_ASAP7_75t_L g6411 ( 
.A1(n_6101),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.C(n_296),
.Y(n_6411)
);

OR2x2_ASAP7_75t_L g6412 ( 
.A(n_6256),
.B(n_294),
.Y(n_6412)
);

HB1xp67_ASAP7_75t_L g6413 ( 
.A(n_6213),
.Y(n_6413)
);

OAI22xp5_ASAP7_75t_L g6414 ( 
.A1(n_6082),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_6414)
);

AND2x2_ASAP7_75t_L g6415 ( 
.A(n_6186),
.B(n_299),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_6238),
.Y(n_6416)
);

OA21x2_ASAP7_75t_L g6417 ( 
.A1(n_6220),
.A2(n_299),
.B(n_300),
.Y(n_6417)
);

HB1xp67_ASAP7_75t_L g6418 ( 
.A(n_6213),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_6249),
.Y(n_6419)
);

OA21x2_ASAP7_75t_L g6420 ( 
.A1(n_6064),
.A2(n_300),
.B(n_301),
.Y(n_6420)
);

AO21x2_ASAP7_75t_L g6421 ( 
.A1(n_6190),
.A2(n_302),
.B(n_303),
.Y(n_6421)
);

NAND2xp5_ASAP7_75t_L g6422 ( 
.A(n_6209),
.B(n_304),
.Y(n_6422)
);

NAND2xp5_ASAP7_75t_L g6423 ( 
.A(n_6231),
.B(n_304),
.Y(n_6423)
);

OR2x2_ASAP7_75t_L g6424 ( 
.A(n_6148),
.B(n_305),
.Y(n_6424)
);

OAI21x1_ASAP7_75t_L g6425 ( 
.A1(n_6038),
.A2(n_6080),
.B(n_6085),
.Y(n_6425)
);

OR2x2_ASAP7_75t_L g6426 ( 
.A(n_6255),
.B(n_305),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_6032),
.Y(n_6427)
);

AOI22xp33_ASAP7_75t_L g6428 ( 
.A1(n_6221),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_6428)
);

INVx2_ASAP7_75t_L g6429 ( 
.A(n_6207),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6193),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6195),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_6036),
.Y(n_6432)
);

INVx2_ASAP7_75t_L g6433 ( 
.A(n_6058),
.Y(n_6433)
);

OR2x2_ASAP7_75t_L g6434 ( 
.A(n_6218),
.B(n_306),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_6171),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6219),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_6208),
.B(n_6235),
.Y(n_6437)
);

AND2x4_ASAP7_75t_L g6438 ( 
.A(n_6188),
.B(n_307),
.Y(n_6438)
);

HB1xp67_ASAP7_75t_L g6439 ( 
.A(n_6237),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6171),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_6157),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_6229),
.Y(n_6442)
);

OA21x2_ASAP7_75t_L g6443 ( 
.A1(n_6239),
.A2(n_308),
.B(n_310),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_6243),
.B(n_311),
.Y(n_6444)
);

OA21x2_ASAP7_75t_L g6445 ( 
.A1(n_6125),
.A2(n_312),
.B(n_313),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6208),
.B(n_313),
.Y(n_6446)
);

AO21x2_ASAP7_75t_L g6447 ( 
.A1(n_6268),
.A2(n_315),
.B(n_316),
.Y(n_6447)
);

INVx4_ASAP7_75t_L g6448 ( 
.A(n_6082),
.Y(n_6448)
);

OAI21xp5_ASAP7_75t_L g6449 ( 
.A1(n_6173),
.A2(n_6152),
.B(n_6079),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6177),
.Y(n_6450)
);

OAI321xp33_ASAP7_75t_L g6451 ( 
.A1(n_6198),
.A2(n_319),
.A3(n_321),
.B1(n_315),
.B2(n_318),
.C(n_320),
.Y(n_6451)
);

OA21x2_ASAP7_75t_L g6452 ( 
.A1(n_6130),
.A2(n_318),
.B(n_319),
.Y(n_6452)
);

AO21x2_ASAP7_75t_L g6453 ( 
.A1(n_6276),
.A2(n_322),
.B(n_323),
.Y(n_6453)
);

AOI21xp5_ASAP7_75t_SL g6454 ( 
.A1(n_6105),
.A2(n_324),
.B(n_325),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_6224),
.B(n_324),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6204),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_6210),
.Y(n_6457)
);

OR2x2_ASAP7_75t_L g6458 ( 
.A(n_6143),
.B(n_325),
.Y(n_6458)
);

AND2x2_ASAP7_75t_L g6459 ( 
.A(n_6041),
.B(n_326),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6270),
.Y(n_6460)
);

OAI21xp5_ASAP7_75t_L g6461 ( 
.A1(n_6214),
.A2(n_328),
.B(n_329),
.Y(n_6461)
);

AND2x2_ASAP7_75t_L g6462 ( 
.A(n_6027),
.B(n_330),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_6034),
.Y(n_6463)
);

NAND4xp25_ASAP7_75t_L g6464 ( 
.A(n_6197),
.B(n_334),
.C(n_332),
.D(n_333),
.Y(n_6464)
);

HB1xp67_ASAP7_75t_L g6465 ( 
.A(n_6191),
.Y(n_6465)
);

OA21x2_ASAP7_75t_L g6466 ( 
.A1(n_6139),
.A2(n_332),
.B(n_335),
.Y(n_6466)
);

BUFx3_ASAP7_75t_L g6467 ( 
.A(n_6180),
.Y(n_6467)
);

INVx2_ASAP7_75t_L g6468 ( 
.A(n_6157),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_6094),
.Y(n_6469)
);

INVx2_ASAP7_75t_L g6470 ( 
.A(n_6096),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_6033),
.Y(n_6471)
);

AND2x2_ASAP7_75t_L g6472 ( 
.A(n_6144),
.B(n_336),
.Y(n_6472)
);

OAI22xp5_ASAP7_75t_L g6473 ( 
.A1(n_6225),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_6473)
);

AND2x2_ASAP7_75t_L g6474 ( 
.A(n_6065),
.B(n_340),
.Y(n_6474)
);

INVx2_ASAP7_75t_L g6475 ( 
.A(n_6049),
.Y(n_6475)
);

OA21x2_ASAP7_75t_L g6476 ( 
.A1(n_6178),
.A2(n_340),
.B(n_341),
.Y(n_6476)
);

INVx2_ASAP7_75t_SL g6477 ( 
.A(n_6067),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_6175),
.Y(n_6478)
);

AOI221xp5_ASAP7_75t_L g6479 ( 
.A1(n_6240),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_6479)
);

OR2x2_ASAP7_75t_L g6480 ( 
.A(n_6224),
.B(n_343),
.Y(n_6480)
);

INVx3_ASAP7_75t_L g6481 ( 
.A(n_6188),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_6049),
.Y(n_6482)
);

INVx2_ASAP7_75t_L g6483 ( 
.A(n_6211),
.Y(n_6483)
);

NOR2xp33_ASAP7_75t_L g6484 ( 
.A(n_6183),
.B(n_344),
.Y(n_6484)
);

AND2x2_ASAP7_75t_L g6485 ( 
.A(n_6081),
.B(n_346),
.Y(n_6485)
);

HB1xp67_ASAP7_75t_L g6486 ( 
.A(n_6191),
.Y(n_6486)
);

AND2x4_ASAP7_75t_L g6487 ( 
.A(n_6106),
.B(n_6158),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_6211),
.Y(n_6488)
);

OA21x2_ASAP7_75t_L g6489 ( 
.A1(n_6258),
.A2(n_347),
.B(n_350),
.Y(n_6489)
);

INVx2_ASAP7_75t_SL g6490 ( 
.A(n_6167),
.Y(n_6490)
);

OAI211xp5_ASAP7_75t_L g6491 ( 
.A1(n_6170),
.A2(n_352),
.B(n_347),
.C(n_350),
.Y(n_6491)
);

INVx1_ASAP7_75t_L g6492 ( 
.A(n_6176),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6224),
.B(n_352),
.Y(n_6493)
);

AO21x2_ASAP7_75t_L g6494 ( 
.A1(n_6140),
.A2(n_353),
.B(n_354),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6043),
.Y(n_6495)
);

CKINVDCx5p33_ASAP7_75t_R g6496 ( 
.A(n_6035),
.Y(n_6496)
);

AND2x4_ASAP7_75t_L g6497 ( 
.A(n_6106),
.B(n_6158),
.Y(n_6497)
);

AOI21xp5_ASAP7_75t_SL g6498 ( 
.A1(n_6112),
.A2(n_353),
.B(n_355),
.Y(n_6498)
);

NAND2xp5_ASAP7_75t_L g6499 ( 
.A(n_6259),
.B(n_355),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_6051),
.Y(n_6500)
);

AND2x2_ASAP7_75t_L g6501 ( 
.A(n_6120),
.B(n_356),
.Y(n_6501)
);

BUFx2_ASAP7_75t_L g6502 ( 
.A(n_6185),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6252),
.Y(n_6503)
);

INVx2_ASAP7_75t_SL g6504 ( 
.A(n_6192),
.Y(n_6504)
);

AO21x2_ASAP7_75t_L g6505 ( 
.A1(n_6174),
.A2(n_357),
.B(n_359),
.Y(n_6505)
);

AO21x2_ASAP7_75t_L g6506 ( 
.A1(n_6057),
.A2(n_357),
.B(n_359),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_6100),
.Y(n_6507)
);

CKINVDCx6p67_ASAP7_75t_R g6508 ( 
.A(n_6048),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_SL g6509 ( 
.A(n_6156),
.B(n_360),
.Y(n_6509)
);

AO21x2_ASAP7_75t_L g6510 ( 
.A1(n_6056),
.A2(n_360),
.B(n_361),
.Y(n_6510)
);

AOI22xp33_ASAP7_75t_L g6511 ( 
.A1(n_6253),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_6159),
.Y(n_6512)
);

AND2x2_ASAP7_75t_L g6513 ( 
.A(n_6132),
.B(n_362),
.Y(n_6513)
);

OA21x2_ASAP7_75t_L g6514 ( 
.A1(n_6172),
.A2(n_6260),
.B(n_6117),
.Y(n_6514)
);

HB1xp67_ASAP7_75t_L g6515 ( 
.A(n_6191),
.Y(n_6515)
);

AND2x2_ASAP7_75t_L g6516 ( 
.A(n_6134),
.B(n_363),
.Y(n_6516)
);

OAI22xp5_ASAP7_75t_L g6517 ( 
.A1(n_6121),
.A2(n_6217),
.B1(n_6251),
.B2(n_6264),
.Y(n_6517)
);

AND2x2_ASAP7_75t_L g6518 ( 
.A(n_6090),
.B(n_364),
.Y(n_6518)
);

NOR2x1_ASAP7_75t_R g6519 ( 
.A(n_6135),
.B(n_365),
.Y(n_6519)
);

INVx3_ASAP7_75t_L g6520 ( 
.A(n_6159),
.Y(n_6520)
);

BUFx3_ASAP7_75t_L g6521 ( 
.A(n_6107),
.Y(n_6521)
);

AO21x2_ASAP7_75t_L g6522 ( 
.A1(n_6044),
.A2(n_366),
.B(n_368),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_6354),
.Y(n_6523)
);

INVx2_ASAP7_75t_L g6524 ( 
.A(n_6405),
.Y(n_6524)
);

AND2x2_ASAP7_75t_L g6525 ( 
.A(n_6317),
.B(n_6100),
.Y(n_6525)
);

OAI22xp5_ASAP7_75t_L g6526 ( 
.A1(n_6278),
.A2(n_6084),
.B1(n_6250),
.B2(n_6263),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_6354),
.Y(n_6527)
);

AND2x2_ASAP7_75t_L g6528 ( 
.A(n_6289),
.B(n_6361),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_6367),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6294),
.B(n_6100),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6343),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6361),
.B(n_6153),
.Y(n_6532)
);

BUFx3_ASAP7_75t_L g6533 ( 
.A(n_6467),
.Y(n_6533)
);

AOI22xp5_ASAP7_75t_L g6534 ( 
.A1(n_6359),
.A2(n_6136),
.B1(n_6253),
.B2(n_6227),
.Y(n_6534)
);

AOI221xp5_ASAP7_75t_L g6535 ( 
.A1(n_6294),
.A2(n_6205),
.B1(n_6165),
.B2(n_6212),
.C(n_6241),
.Y(n_6535)
);

AND2x2_ASAP7_75t_L g6536 ( 
.A(n_6374),
.B(n_6189),
.Y(n_6536)
);

BUFx3_ASAP7_75t_L g6537 ( 
.A(n_6467),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_6343),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_6374),
.B(n_6091),
.Y(n_6539)
);

BUFx3_ASAP7_75t_L g6540 ( 
.A(n_6331),
.Y(n_6540)
);

AND2x4_ASAP7_75t_SL g6541 ( 
.A(n_6508),
.B(n_6103),
.Y(n_6541)
);

OR2x2_ASAP7_75t_L g6542 ( 
.A(n_6290),
.B(n_6179),
.Y(n_6542)
);

AND2x2_ASAP7_75t_L g6543 ( 
.A(n_6481),
.B(n_6109),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_6280),
.Y(n_6544)
);

NAND2xp5_ASAP7_75t_L g6545 ( 
.A(n_6279),
.B(n_6206),
.Y(n_6545)
);

OAI22xp5_ASAP7_75t_L g6546 ( 
.A1(n_6278),
.A2(n_6179),
.B1(n_6247),
.B2(n_6226),
.Y(n_6546)
);

NOR3xp33_ASAP7_75t_L g6547 ( 
.A(n_6411),
.B(n_6151),
.C(n_6187),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_6367),
.Y(n_6548)
);

INVxp67_ASAP7_75t_SL g6549 ( 
.A(n_6359),
.Y(n_6549)
);

INVx2_ASAP7_75t_L g6550 ( 
.A(n_6367),
.Y(n_6550)
);

OR2x2_ASAP7_75t_L g6551 ( 
.A(n_6285),
.B(n_6030),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_6281),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6292),
.Y(n_6553)
);

INVx2_ASAP7_75t_SL g6554 ( 
.A(n_6344),
.Y(n_6554)
);

AND2x4_ASAP7_75t_L g6555 ( 
.A(n_6448),
.B(n_6046),
.Y(n_6555)
);

CKINVDCx6p67_ASAP7_75t_R g6556 ( 
.A(n_6331),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_6279),
.B(n_6030),
.Y(n_6557)
);

INVx1_ASAP7_75t_L g6558 ( 
.A(n_6299),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6481),
.B(n_6115),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6413),
.Y(n_6560)
);

INVx1_ASAP7_75t_L g6561 ( 
.A(n_6413),
.Y(n_6561)
);

INVx3_ASAP7_75t_L g6562 ( 
.A(n_6300),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6418),
.Y(n_6563)
);

OR2x2_ASAP7_75t_L g6564 ( 
.A(n_6283),
.B(n_6246),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_6418),
.Y(n_6565)
);

HB1xp67_ASAP7_75t_L g6566 ( 
.A(n_6298),
.Y(n_6566)
);

NOR2xp67_ASAP7_75t_L g6567 ( 
.A(n_6448),
.B(n_6110),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_6393),
.B(n_6200),
.Y(n_6568)
);

OR2x2_ASAP7_75t_L g6569 ( 
.A(n_6283),
.B(n_6470),
.Y(n_6569)
);

OR2x2_ASAP7_75t_L g6570 ( 
.A(n_6470),
.B(n_6166),
.Y(n_6570)
);

OR2x2_ASAP7_75t_L g6571 ( 
.A(n_6373),
.B(n_6149),
.Y(n_6571)
);

INVx2_ASAP7_75t_L g6572 ( 
.A(n_6367),
.Y(n_6572)
);

NAND2xp5_ASAP7_75t_L g6573 ( 
.A(n_6393),
.B(n_6169),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_6437),
.B(n_6045),
.Y(n_6574)
);

AND2x2_ASAP7_75t_L g6575 ( 
.A(n_6502),
.B(n_6181),
.Y(n_6575)
);

OR2x2_ASAP7_75t_L g6576 ( 
.A(n_6375),
.B(n_6138),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_6443),
.B(n_6059),
.Y(n_6577)
);

OR2x2_ASAP7_75t_L g6578 ( 
.A(n_6282),
.B(n_6088),
.Y(n_6578)
);

AND2x4_ASAP7_75t_SL g6579 ( 
.A(n_6300),
.B(n_366),
.Y(n_6579)
);

BUFx2_ASAP7_75t_L g6580 ( 
.A(n_6344),
.Y(n_6580)
);

NAND2xp67_ASAP7_75t_L g6581 ( 
.A(n_6446),
.B(n_368),
.Y(n_6581)
);

AND2x2_ASAP7_75t_L g6582 ( 
.A(n_6319),
.B(n_369),
.Y(n_6582)
);

INVx2_ASAP7_75t_L g6583 ( 
.A(n_6344),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6443),
.B(n_369),
.Y(n_6584)
);

INVx2_ASAP7_75t_L g6585 ( 
.A(n_6344),
.Y(n_6585)
);

INVx2_ASAP7_75t_L g6586 ( 
.A(n_6349),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6298),
.Y(n_6587)
);

OR2x2_ASAP7_75t_L g6588 ( 
.A(n_6306),
.B(n_372),
.Y(n_6588)
);

OR2x2_ASAP7_75t_L g6589 ( 
.A(n_6307),
.B(n_372),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6349),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_6322),
.B(n_376),
.Y(n_6591)
);

NAND2xp5_ASAP7_75t_L g6592 ( 
.A(n_6443),
.B(n_378),
.Y(n_6592)
);

OR2x2_ASAP7_75t_L g6593 ( 
.A(n_6396),
.B(n_378),
.Y(n_6593)
);

AND2x2_ASAP7_75t_L g6594 ( 
.A(n_6487),
.B(n_381),
.Y(n_6594)
);

AOI22xp33_ASAP7_75t_L g6595 ( 
.A1(n_6329),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_6595)
);

AND2x2_ASAP7_75t_L g6596 ( 
.A(n_6487),
.B(n_383),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_L g6597 ( 
.A(n_6416),
.B(n_384),
.Y(n_6597)
);

NAND2xp5_ASAP7_75t_L g6598 ( 
.A(n_6419),
.B(n_6301),
.Y(n_6598)
);

AND2x4_ASAP7_75t_L g6599 ( 
.A(n_6497),
.B(n_387),
.Y(n_6599)
);

INVx1_ASAP7_75t_SL g6600 ( 
.A(n_6407),
.Y(n_6600)
);

AND2x2_ASAP7_75t_L g6601 ( 
.A(n_6497),
.B(n_387),
.Y(n_6601)
);

OAI22xp5_ASAP7_75t_L g6602 ( 
.A1(n_6302),
.A2(n_392),
.B1(n_389),
.B2(n_390),
.Y(n_6602)
);

OR2x2_ASAP7_75t_L g6603 ( 
.A(n_6382),
.B(n_390),
.Y(n_6603)
);

INVx2_ASAP7_75t_L g6604 ( 
.A(n_6477),
.Y(n_6604)
);

INVx2_ASAP7_75t_L g6605 ( 
.A(n_6395),
.Y(n_6605)
);

NAND2xp5_ASAP7_75t_SL g6606 ( 
.A(n_6449),
.B(n_1995),
.Y(n_6606)
);

OR2x2_ASAP7_75t_L g6607 ( 
.A(n_6399),
.B(n_392),
.Y(n_6607)
);

HB1xp67_ASAP7_75t_L g6608 ( 
.A(n_6323),
.Y(n_6608)
);

OR2x2_ASAP7_75t_L g6609 ( 
.A(n_6312),
.B(n_6471),
.Y(n_6609)
);

AND2x2_ASAP7_75t_L g6610 ( 
.A(n_6483),
.B(n_394),
.Y(n_6610)
);

OR2x2_ASAP7_75t_L g6611 ( 
.A(n_6427),
.B(n_6460),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_6323),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6304),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6305),
.Y(n_6614)
);

AND2x4_ASAP7_75t_SL g6615 ( 
.A(n_6438),
.B(n_395),
.Y(n_6615)
);

INVx2_ASAP7_75t_L g6616 ( 
.A(n_6395),
.Y(n_6616)
);

INVx5_ASAP7_75t_L g6617 ( 
.A(n_6376),
.Y(n_6617)
);

HB1xp67_ASAP7_75t_L g6618 ( 
.A(n_6489),
.Y(n_6618)
);

HB1xp67_ASAP7_75t_L g6619 ( 
.A(n_6489),
.Y(n_6619)
);

AND2x2_ASAP7_75t_L g6620 ( 
.A(n_6488),
.B(n_395),
.Y(n_6620)
);

AOI22xp33_ASAP7_75t_L g6621 ( 
.A1(n_6329),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_6621)
);

OR2x2_ASAP7_75t_L g6622 ( 
.A(n_6427),
.B(n_396),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6520),
.Y(n_6623)
);

AND2x2_ASAP7_75t_L g6624 ( 
.A(n_6475),
.B(n_397),
.Y(n_6624)
);

NAND2xp5_ASAP7_75t_L g6625 ( 
.A(n_6301),
.B(n_399),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6482),
.B(n_400),
.Y(n_6626)
);

AND2x2_ASAP7_75t_L g6627 ( 
.A(n_6402),
.B(n_400),
.Y(n_6627)
);

AOI22xp33_ASAP7_75t_L g6628 ( 
.A1(n_6302),
.A2(n_404),
.B1(n_401),
.B2(n_402),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6310),
.Y(n_6629)
);

INVx2_ASAP7_75t_L g6630 ( 
.A(n_6520),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6318),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_6295),
.Y(n_6632)
);

INVx1_ASAP7_75t_SL g6633 ( 
.A(n_6407),
.Y(n_6633)
);

INVx2_ASAP7_75t_L g6634 ( 
.A(n_6313),
.Y(n_6634)
);

NAND2xp5_ASAP7_75t_L g6635 ( 
.A(n_6301),
.B(n_402),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6441),
.Y(n_6636)
);

AND2x2_ASAP7_75t_L g6637 ( 
.A(n_6409),
.B(n_404),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6333),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_6512),
.B(n_405),
.Y(n_6639)
);

AOI22xp33_ASAP7_75t_L g6640 ( 
.A1(n_6314),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_6640)
);

OR2x2_ASAP7_75t_L g6641 ( 
.A(n_6463),
.B(n_406),
.Y(n_6641)
);

NAND2xp5_ASAP7_75t_L g6642 ( 
.A(n_6370),
.B(n_407),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6342),
.Y(n_6643)
);

AND2x2_ASAP7_75t_L g6644 ( 
.A(n_6429),
.B(n_409),
.Y(n_6644)
);

AND2x2_ASAP7_75t_L g6645 ( 
.A(n_6468),
.B(n_409),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6348),
.Y(n_6646)
);

AND2x2_ASAP7_75t_L g6647 ( 
.A(n_6478),
.B(n_410),
.Y(n_6647)
);

AOI22xp33_ASAP7_75t_L g6648 ( 
.A1(n_6327),
.A2(n_413),
.B1(n_410),
.B2(n_411),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6357),
.Y(n_6649)
);

HB1xp67_ASAP7_75t_L g6650 ( 
.A(n_6489),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6492),
.B(n_414),
.Y(n_6651)
);

INVxp67_ASAP7_75t_L g6652 ( 
.A(n_6421),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_L g6653 ( 
.A(n_6439),
.B(n_415),
.Y(n_6653)
);

INVx2_ASAP7_75t_L g6654 ( 
.A(n_6339),
.Y(n_6654)
);

OR2x2_ASAP7_75t_L g6655 ( 
.A(n_6355),
.B(n_415),
.Y(n_6655)
);

INVx8_ASAP7_75t_L g6656 ( 
.A(n_6376),
.Y(n_6656)
);

OAI222xp33_ASAP7_75t_L g6657 ( 
.A1(n_6330),
.A2(n_417),
.B1(n_419),
.B2(n_420),
.C1(n_421),
.C2(n_422),
.Y(n_6657)
);

AND2x2_ASAP7_75t_L g6658 ( 
.A(n_6335),
.B(n_417),
.Y(n_6658)
);

AND2x4_ASAP7_75t_L g6659 ( 
.A(n_6435),
.B(n_422),
.Y(n_6659)
);

AND2x2_ASAP7_75t_L g6660 ( 
.A(n_6440),
.B(n_423),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6368),
.B(n_423),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6365),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6366),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6369),
.Y(n_6664)
);

INVxp67_ASAP7_75t_L g6665 ( 
.A(n_6421),
.Y(n_6665)
);

NAND2xp5_ASAP7_75t_L g6666 ( 
.A(n_6439),
.B(n_6387),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6404),
.Y(n_6667)
);

AOI22xp33_ASAP7_75t_L g6668 ( 
.A1(n_6314),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6364),
.Y(n_6669)
);

HB1xp67_ASAP7_75t_L g6670 ( 
.A(n_6394),
.Y(n_6670)
);

AND2x2_ASAP7_75t_L g6671 ( 
.A(n_6286),
.B(n_424),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6364),
.Y(n_6672)
);

BUFx3_ASAP7_75t_L g6673 ( 
.A(n_6521),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6286),
.B(n_425),
.Y(n_6674)
);

INVxp67_ASAP7_75t_SL g6675 ( 
.A(n_6480),
.Y(n_6675)
);

INVx2_ASAP7_75t_L g6676 ( 
.A(n_6339),
.Y(n_6676)
);

INVxp33_ASAP7_75t_SL g6677 ( 
.A(n_6519),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6500),
.B(n_426),
.Y(n_6678)
);

AND2x2_ASAP7_75t_L g6679 ( 
.A(n_6341),
.B(n_428),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6388),
.Y(n_6680)
);

AND2x2_ASAP7_75t_SL g6681 ( 
.A(n_6316),
.B(n_428),
.Y(n_6681)
);

AND2x2_ASAP7_75t_L g6682 ( 
.A(n_6337),
.B(n_429),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_6388),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6401),
.Y(n_6684)
);

AND2x4_ASAP7_75t_L g6685 ( 
.A(n_6407),
.B(n_431),
.Y(n_6685)
);

NOR2xp67_ASAP7_75t_L g6686 ( 
.A(n_6309),
.B(n_431),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6401),
.Y(n_6687)
);

INVxp67_ASAP7_75t_L g6688 ( 
.A(n_6316),
.Y(n_6688)
);

INVx2_ASAP7_75t_L g6689 ( 
.A(n_6311),
.Y(n_6689)
);

INVx3_ASAP7_75t_L g6690 ( 
.A(n_6438),
.Y(n_6690)
);

OR2x2_ASAP7_75t_L g6691 ( 
.A(n_6355),
.B(n_432),
.Y(n_6691)
);

OR2x2_ASAP7_75t_L g6692 ( 
.A(n_6303),
.B(n_6324),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6410),
.Y(n_6693)
);

BUFx2_ASAP7_75t_L g6694 ( 
.A(n_6376),
.Y(n_6694)
);

AND2x4_ASAP7_75t_L g6695 ( 
.A(n_6347),
.B(n_432),
.Y(n_6695)
);

BUFx6f_ASAP7_75t_L g6696 ( 
.A(n_6371),
.Y(n_6696)
);

INVx2_ASAP7_75t_L g6697 ( 
.A(n_6315),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6452),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6452),
.Y(n_6699)
);

CKINVDCx20_ASAP7_75t_R g6700 ( 
.A(n_6496),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6315),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6469),
.B(n_433),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6452),
.Y(n_6703)
);

INVx2_ASAP7_75t_L g6704 ( 
.A(n_6350),
.Y(n_6704)
);

INVxp67_ASAP7_75t_SL g6705 ( 
.A(n_6455),
.Y(n_6705)
);

AND2x2_ASAP7_75t_L g6706 ( 
.A(n_6456),
.B(n_435),
.Y(n_6706)
);

BUFx2_ASAP7_75t_L g6707 ( 
.A(n_6347),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6457),
.B(n_436),
.Y(n_6708)
);

OAI22xp5_ASAP7_75t_L g6709 ( 
.A1(n_6330),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_6709)
);

NAND2xp5_ASAP7_75t_L g6710 ( 
.A(n_6296),
.B(n_437),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6347),
.B(n_438),
.Y(n_6711)
);

HB1xp67_ASAP7_75t_L g6712 ( 
.A(n_6394),
.Y(n_6712)
);

INVx1_ASAP7_75t_L g6713 ( 
.A(n_6430),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6431),
.Y(n_6714)
);

AOI22xp33_ASAP7_75t_L g6715 ( 
.A1(n_6327),
.A2(n_442),
.B1(n_439),
.B2(n_441),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_6432),
.Y(n_6716)
);

BUFx2_ASAP7_75t_L g6717 ( 
.A(n_6505),
.Y(n_6717)
);

OR2x2_ASAP7_75t_L g6718 ( 
.A(n_6433),
.B(n_439),
.Y(n_6718)
);

NAND2xp5_ASAP7_75t_L g6719 ( 
.A(n_6296),
.B(n_441),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6436),
.Y(n_6720)
);

INVx1_ASAP7_75t_SL g6721 ( 
.A(n_6505),
.Y(n_6721)
);

OR2x2_ASAP7_75t_L g6722 ( 
.A(n_6351),
.B(n_443),
.Y(n_6722)
);

AND2x4_ASAP7_75t_L g6723 ( 
.A(n_6495),
.B(n_6504),
.Y(n_6723)
);

OR2x2_ASAP7_75t_L g6724 ( 
.A(n_6293),
.B(n_443),
.Y(n_6724)
);

AOI22xp33_ASAP7_75t_SL g6725 ( 
.A1(n_6288),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_6725)
);

NOR2xp33_ASAP7_75t_L g6726 ( 
.A(n_6521),
.B(n_6372),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_6291),
.B(n_445),
.Y(n_6727)
);

AND2x4_ASAP7_75t_L g6728 ( 
.A(n_6320),
.B(n_447),
.Y(n_6728)
);

INVx1_ASAP7_75t_SL g6729 ( 
.A(n_6494),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6442),
.Y(n_6730)
);

AND2x2_ASAP7_75t_L g6731 ( 
.A(n_6291),
.B(n_449),
.Y(n_6731)
);

INVx2_ASAP7_75t_L g6732 ( 
.A(n_6380),
.Y(n_6732)
);

AND2x2_ASAP7_75t_L g6733 ( 
.A(n_6291),
.B(n_450),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6450),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_6499),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6503),
.B(n_451),
.Y(n_6736)
);

INVx2_ASAP7_75t_SL g6737 ( 
.A(n_6490),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6499),
.Y(n_6738)
);

INVx2_ASAP7_75t_L g6739 ( 
.A(n_6386),
.Y(n_6739)
);

BUFx2_ASAP7_75t_L g6740 ( 
.A(n_6381),
.Y(n_6740)
);

NAND2xp5_ASAP7_75t_L g6741 ( 
.A(n_6293),
.B(n_451),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6320),
.B(n_454),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_6353),
.Y(n_6743)
);

BUFx3_ASAP7_75t_L g6744 ( 
.A(n_6378),
.Y(n_6744)
);

INVx1_ASAP7_75t_L g6745 ( 
.A(n_6353),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6423),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_L g6747 ( 
.A(n_6293),
.B(n_455),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6423),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6425),
.B(n_456),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_6377),
.Y(n_6750)
);

NAND2xp5_ASAP7_75t_L g6751 ( 
.A(n_6455),
.B(n_457),
.Y(n_6751)
);

INVx3_ASAP7_75t_L g6752 ( 
.A(n_6381),
.Y(n_6752)
);

NAND4xp25_ASAP7_75t_L g6753 ( 
.A(n_6628),
.B(n_6461),
.C(n_6288),
.D(n_6479),
.Y(n_6753)
);

BUFx2_ASAP7_75t_L g6754 ( 
.A(n_6556),
.Y(n_6754)
);

AND2x2_ASAP7_75t_L g6755 ( 
.A(n_6575),
.B(n_6297),
.Y(n_6755)
);

NOR2xp33_ASAP7_75t_R g6756 ( 
.A(n_6700),
.B(n_6484),
.Y(n_6756)
);

BUFx3_ASAP7_75t_L g6757 ( 
.A(n_6541),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6566),
.Y(n_6758)
);

NOR2xp33_ASAP7_75t_R g6759 ( 
.A(n_6656),
.B(n_6484),
.Y(n_6759)
);

AND2x2_ASAP7_75t_L g6760 ( 
.A(n_6528),
.B(n_6297),
.Y(n_6760)
);

OAI22xp5_ASAP7_75t_L g6761 ( 
.A1(n_6534),
.A2(n_6400),
.B1(n_6449),
.B2(n_6334),
.Y(n_6761)
);

BUFx3_ASAP7_75t_L g6762 ( 
.A(n_6540),
.Y(n_6762)
);

OAI22xp5_ASAP7_75t_L g6763 ( 
.A1(n_6534),
.A2(n_6428),
.B1(n_6297),
.B2(n_6336),
.Y(n_6763)
);

OAI22xp5_ASAP7_75t_L g6764 ( 
.A1(n_6546),
.A2(n_6428),
.B1(n_6336),
.B2(n_6461),
.Y(n_6764)
);

AND2x2_ASAP7_75t_L g6765 ( 
.A(n_6532),
.B(n_6514),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6566),
.Y(n_6766)
);

AOI221xp5_ASAP7_75t_L g6767 ( 
.A1(n_6546),
.A2(n_6411),
.B1(n_6479),
.B2(n_6326),
.C(n_6464),
.Y(n_6767)
);

OA21x2_ASAP7_75t_L g6768 ( 
.A1(n_6740),
.A2(n_6665),
.B(n_6652),
.Y(n_6768)
);

OAI33xp33_ASAP7_75t_L g6769 ( 
.A1(n_6602),
.A2(n_6526),
.A3(n_6652),
.B1(n_6665),
.B2(n_6688),
.B3(n_6709),
.Y(n_6769)
);

AO221x2_ASAP7_75t_L g6770 ( 
.A1(n_6526),
.A2(n_6473),
.B1(n_6383),
.B2(n_6517),
.C(n_6493),
.Y(n_6770)
);

AOI33xp33_ASAP7_75t_L g6771 ( 
.A1(n_6725),
.A2(n_6511),
.A3(n_6415),
.B1(n_6507),
.B2(n_6360),
.B3(n_6308),
.Y(n_6771)
);

AND2x2_ASAP7_75t_L g6772 ( 
.A(n_6574),
.B(n_6514),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6608),
.Y(n_6773)
);

HB1xp67_ASAP7_75t_L g6774 ( 
.A(n_6608),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_6688),
.B(n_6345),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6587),
.Y(n_6776)
);

NAND2xp33_ASAP7_75t_R g6777 ( 
.A(n_6677),
.B(n_6420),
.Y(n_6777)
);

INVxp67_ASAP7_75t_L g6778 ( 
.A(n_6717),
.Y(n_6778)
);

INVx2_ASAP7_75t_L g6779 ( 
.A(n_6533),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6543),
.B(n_6514),
.Y(n_6780)
);

INVx2_ASAP7_75t_L g6781 ( 
.A(n_6537),
.Y(n_6781)
);

NAND3xp33_ASAP7_75t_L g6782 ( 
.A(n_6628),
.B(n_6511),
.C(n_6493),
.Y(n_6782)
);

AO21x2_ASAP7_75t_L g6783 ( 
.A1(n_6741),
.A2(n_6287),
.B(n_6465),
.Y(n_6783)
);

NAND4xp25_ASAP7_75t_L g6784 ( 
.A(n_6602),
.B(n_6384),
.C(n_6379),
.D(n_6383),
.Y(n_6784)
);

OAI31xp33_ASAP7_75t_L g6785 ( 
.A1(n_6709),
.A2(n_6491),
.A3(n_6473),
.B(n_6509),
.Y(n_6785)
);

BUFx2_ASAP7_75t_L g6786 ( 
.A(n_6656),
.Y(n_6786)
);

AND2x2_ASAP7_75t_L g6787 ( 
.A(n_6559),
.B(n_6345),
.Y(n_6787)
);

OR2x2_ASAP7_75t_L g6788 ( 
.A(n_6577),
.B(n_6287),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6560),
.Y(n_6789)
);

NOR4xp25_ASAP7_75t_SL g6790 ( 
.A(n_6549),
.B(n_6509),
.C(n_6451),
.D(n_6510),
.Y(n_6790)
);

BUFx6f_ASAP7_75t_L g6791 ( 
.A(n_6639),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_6561),
.Y(n_6792)
);

AND2x2_ASAP7_75t_L g6793 ( 
.A(n_6536),
.B(n_6485),
.Y(n_6793)
);

OAI21xp5_ASAP7_75t_L g6794 ( 
.A1(n_6725),
.A2(n_6403),
.B(n_6498),
.Y(n_6794)
);

NOR2xp33_ASAP7_75t_L g6795 ( 
.A(n_6673),
.B(n_6444),
.Y(n_6795)
);

OAI22xp5_ASAP7_75t_L g6796 ( 
.A1(n_6549),
.A2(n_6517),
.B1(n_6356),
.B2(n_6454),
.Y(n_6796)
);

INVx1_ASAP7_75t_SL g6797 ( 
.A(n_6617),
.Y(n_6797)
);

OAI211xp5_ASAP7_75t_SL g6798 ( 
.A1(n_6547),
.A2(n_6444),
.B(n_6491),
.C(n_6422),
.Y(n_6798)
);

OAI22xp5_ASAP7_75t_L g6799 ( 
.A1(n_6729),
.A2(n_6356),
.B1(n_6420),
.B2(n_6325),
.Y(n_6799)
);

OAI22xp5_ASAP7_75t_L g6800 ( 
.A1(n_6729),
.A2(n_6356),
.B1(n_6420),
.B2(n_6325),
.Y(n_6800)
);

AOI222xp33_ASAP7_75t_L g6801 ( 
.A1(n_6710),
.A2(n_6451),
.B1(n_6379),
.B2(n_6422),
.C1(n_6414),
.C2(n_6397),
.Y(n_6801)
);

AOI22xp33_ASAP7_75t_L g6802 ( 
.A1(n_6547),
.A2(n_6728),
.B1(n_6695),
.B2(n_6634),
.Y(n_6802)
);

INVx1_ASAP7_75t_SL g6803 ( 
.A(n_6617),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6690),
.Y(n_6804)
);

OAI211xp5_ASAP7_75t_L g6805 ( 
.A1(n_6648),
.A2(n_6715),
.B(n_6752),
.C(n_6721),
.Y(n_6805)
);

INVx2_ASAP7_75t_L g6806 ( 
.A(n_6690),
.Y(n_6806)
);

OAI332xp33_ASAP7_75t_L g6807 ( 
.A1(n_6721),
.A2(n_6414),
.A3(n_6385),
.B1(n_6398),
.B2(n_6328),
.B3(n_6434),
.C1(n_6424),
.C2(n_6406),
.Y(n_6807)
);

INVx1_ASAP7_75t_SL g6808 ( 
.A(n_6617),
.Y(n_6808)
);

AOI221xp5_ASAP7_75t_L g6809 ( 
.A1(n_6752),
.A2(n_6675),
.B1(n_6705),
.B2(n_6657),
.C(n_6710),
.Y(n_6809)
);

NAND2xp33_ASAP7_75t_R g6810 ( 
.A(n_6728),
.B(n_6417),
.Y(n_6810)
);

OAI22xp5_ASAP7_75t_L g6811 ( 
.A1(n_6577),
.A2(n_6325),
.B1(n_6417),
.B2(n_6284),
.Y(n_6811)
);

OR2x2_ASAP7_75t_L g6812 ( 
.A(n_6568),
.B(n_6412),
.Y(n_6812)
);

NAND3xp33_ASAP7_75t_L g6813 ( 
.A(n_6640),
.B(n_6417),
.C(n_6466),
.Y(n_6813)
);

AND2x2_ASAP7_75t_L g6814 ( 
.A(n_6539),
.B(n_6362),
.Y(n_6814)
);

AND2x2_ASAP7_75t_L g6815 ( 
.A(n_6555),
.B(n_6513),
.Y(n_6815)
);

NAND2xp5_ASAP7_75t_L g6816 ( 
.A(n_6600),
.B(n_6447),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6555),
.B(n_6516),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6563),
.Y(n_6818)
);

OA21x2_ASAP7_75t_L g6819 ( 
.A1(n_6670),
.A2(n_6486),
.B(n_6465),
.Y(n_6819)
);

CKINVDCx5p33_ASAP7_75t_R g6820 ( 
.A(n_6744),
.Y(n_6820)
);

BUFx2_ASAP7_75t_L g6821 ( 
.A(n_6656),
.Y(n_6821)
);

AOI22xp33_ASAP7_75t_L g6822 ( 
.A1(n_6695),
.A2(n_6284),
.B1(n_6332),
.B2(n_6510),
.Y(n_6822)
);

AND2x2_ASAP7_75t_L g6823 ( 
.A(n_6689),
.B(n_6474),
.Y(n_6823)
);

OAI22xp5_ASAP7_75t_L g6824 ( 
.A1(n_6724),
.A2(n_6284),
.B1(n_6445),
.B2(n_6466),
.Y(n_6824)
);

NAND4xp75_ASAP7_75t_L g6825 ( 
.A(n_6742),
.B(n_6445),
.C(n_6389),
.D(n_6466),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6565),
.Y(n_6826)
);

AOI222xp33_ASAP7_75t_L g6827 ( 
.A1(n_6719),
.A2(n_6681),
.B1(n_6657),
.B2(n_6675),
.C1(n_6668),
.C2(n_6640),
.Y(n_6827)
);

OAI211xp5_ASAP7_75t_L g6828 ( 
.A1(n_6668),
.A2(n_6486),
.B(n_6515),
.C(n_6389),
.Y(n_6828)
);

NAND2xp5_ASAP7_75t_L g6829 ( 
.A(n_6600),
.B(n_6447),
.Y(n_6829)
);

AOI33xp33_ASAP7_75t_L g6830 ( 
.A1(n_6595),
.A2(n_6472),
.A3(n_6363),
.B1(n_6346),
.B2(n_6340),
.B3(n_6459),
.Y(n_6830)
);

AOI22xp33_ASAP7_75t_L g6831 ( 
.A1(n_6632),
.A2(n_6332),
.B1(n_6338),
.B2(n_6506),
.Y(n_6831)
);

AND2x2_ASAP7_75t_L g6832 ( 
.A(n_6524),
.B(n_6501),
.Y(n_6832)
);

OAI211xp5_ASAP7_75t_L g6833 ( 
.A1(n_6617),
.A2(n_6515),
.B(n_6389),
.C(n_6338),
.Y(n_6833)
);

INVx1_ASAP7_75t_L g6834 ( 
.A(n_6523),
.Y(n_6834)
);

BUFx2_ASAP7_75t_L g6835 ( 
.A(n_6694),
.Y(n_6835)
);

INVx4_ASAP7_75t_L g6836 ( 
.A(n_6685),
.Y(n_6836)
);

OR2x2_ASAP7_75t_L g6837 ( 
.A(n_6568),
.B(n_6458),
.Y(n_6837)
);

HB1xp67_ASAP7_75t_L g6838 ( 
.A(n_6686),
.Y(n_6838)
);

OR2x2_ASAP7_75t_L g6839 ( 
.A(n_6569),
.B(n_6426),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6707),
.B(n_6518),
.Y(n_6840)
);

INVx1_ASAP7_75t_L g6841 ( 
.A(n_6527),
.Y(n_6841)
);

INVx2_ASAP7_75t_L g6842 ( 
.A(n_6696),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6654),
.B(n_6462),
.Y(n_6843)
);

HB1xp67_ASAP7_75t_L g6844 ( 
.A(n_6633),
.Y(n_6844)
);

AND2x2_ASAP7_75t_L g6845 ( 
.A(n_6676),
.B(n_6737),
.Y(n_6845)
);

OR2x2_ASAP7_75t_L g6846 ( 
.A(n_6573),
.B(n_6385),
.Y(n_6846)
);

NAND2xp5_ASAP7_75t_L g6847 ( 
.A(n_6633),
.B(n_6727),
.Y(n_6847)
);

NAND4xp25_ASAP7_75t_L g6848 ( 
.A(n_6719),
.B(n_6453),
.C(n_6506),
.D(n_6494),
.Y(n_6848)
);

OAI211xp5_ASAP7_75t_L g6849 ( 
.A1(n_6621),
.A2(n_6338),
.B(n_6445),
.C(n_6476),
.Y(n_6849)
);

INVx3_ASAP7_75t_L g6850 ( 
.A(n_6562),
.Y(n_6850)
);

NOR2xp33_ASAP7_75t_L g6851 ( 
.A(n_6726),
.B(n_6576),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6531),
.Y(n_6852)
);

AOI22xp33_ASAP7_75t_L g6853 ( 
.A1(n_6535),
.A2(n_6321),
.B1(n_6453),
.B2(n_6522),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6731),
.B(n_6522),
.Y(n_6854)
);

NAND2xp33_ASAP7_75t_R g6855 ( 
.A(n_6685),
.B(n_6476),
.Y(n_6855)
);

AND2x4_ASAP7_75t_SL g6856 ( 
.A(n_6599),
.B(n_6358),
.Y(n_6856)
);

OAI22xp33_ASAP7_75t_L g6857 ( 
.A1(n_6618),
.A2(n_6476),
.B1(n_6391),
.B2(n_6408),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6733),
.B(n_6390),
.Y(n_6858)
);

AND2x2_ASAP7_75t_L g6859 ( 
.A(n_6623),
.B(n_6390),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6538),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6630),
.B(n_6391),
.Y(n_6861)
);

AO21x2_ASAP7_75t_L g6862 ( 
.A1(n_6741),
.A2(n_6392),
.B(n_6352),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_6567),
.B(n_6391),
.Y(n_6863)
);

A2O1A1Ixp33_ASAP7_75t_L g6864 ( 
.A1(n_6535),
.A2(n_6408),
.B(n_6321),
.C(n_459),
.Y(n_6864)
);

OAI221xp5_ASAP7_75t_SL g6865 ( 
.A1(n_6722),
.A2(n_6530),
.B1(n_6705),
.B2(n_6635),
.C(n_6625),
.Y(n_6865)
);

AND2x2_ASAP7_75t_L g6866 ( 
.A(n_6732),
.B(n_6408),
.Y(n_6866)
);

OAI211xp5_ASAP7_75t_L g6867 ( 
.A1(n_6618),
.A2(n_6321),
.B(n_459),
.C(n_457),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6612),
.Y(n_6868)
);

HB1xp67_ASAP7_75t_L g6869 ( 
.A(n_6573),
.Y(n_6869)
);

INVx2_ASAP7_75t_L g6870 ( 
.A(n_6696),
.Y(n_6870)
);

OAI211xp5_ASAP7_75t_L g6871 ( 
.A1(n_6619),
.A2(n_461),
.B(n_458),
.C(n_460),
.Y(n_6871)
);

INVx2_ASAP7_75t_L g6872 ( 
.A(n_6696),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6562),
.Y(n_6873)
);

NAND3xp33_ASAP7_75t_L g6874 ( 
.A(n_6625),
.B(n_460),
.C(n_461),
.Y(n_6874)
);

AOI22xp33_ASAP7_75t_L g6875 ( 
.A1(n_6606),
.A2(n_465),
.B1(n_462),
.B2(n_464),
.Y(n_6875)
);

INVx2_ASAP7_75t_SL g6876 ( 
.A(n_6579),
.Y(n_6876)
);

NOR4xp25_ASAP7_75t_SL g6877 ( 
.A(n_6580),
.B(n_466),
.C(n_462),
.D(n_464),
.Y(n_6877)
);

AND2x4_ASAP7_75t_SL g6878 ( 
.A(n_6599),
.B(n_466),
.Y(n_6878)
);

OAI221xp5_ASAP7_75t_L g6879 ( 
.A1(n_6530),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.C(n_471),
.Y(n_6879)
);

OR2x2_ASAP7_75t_L g6880 ( 
.A(n_6609),
.B(n_468),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6743),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6745),
.Y(n_6882)
);

OA21x2_ASAP7_75t_L g6883 ( 
.A1(n_6670),
.A2(n_469),
.B(n_472),
.Y(n_6883)
);

CKINVDCx12_ASAP7_75t_R g6884 ( 
.A(n_6582),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6739),
.B(n_474),
.Y(n_6885)
);

BUFx2_ASAP7_75t_L g6886 ( 
.A(n_6723),
.Y(n_6886)
);

OA21x2_ASAP7_75t_L g6887 ( 
.A1(n_6712),
.A2(n_475),
.B(n_476),
.Y(n_6887)
);

AND2x2_ASAP7_75t_L g6888 ( 
.A(n_6604),
.B(n_6723),
.Y(n_6888)
);

INVx1_ASAP7_75t_L g6889 ( 
.A(n_6669),
.Y(n_6889)
);

AND2x2_ASAP7_75t_L g6890 ( 
.A(n_6711),
.B(n_477),
.Y(n_6890)
);

AOI22xp33_ASAP7_75t_L g6891 ( 
.A1(n_6564),
.A2(n_481),
.B1(n_478),
.B2(n_480),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6529),
.Y(n_6892)
);

INVxp67_ASAP7_75t_L g6893 ( 
.A(n_6557),
.Y(n_6893)
);

OAI211xp5_ASAP7_75t_L g6894 ( 
.A1(n_6619),
.A2(n_6650),
.B(n_6635),
.C(n_6747),
.Y(n_6894)
);

OAI21xp5_ASAP7_75t_L g6895 ( 
.A1(n_6747),
.A2(n_480),
.B(n_481),
.Y(n_6895)
);

BUFx3_ASAP7_75t_L g6896 ( 
.A(n_6615),
.Y(n_6896)
);

INVx2_ASAP7_75t_L g6897 ( 
.A(n_6548),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6672),
.Y(n_6898)
);

NAND2xp5_ASAP7_75t_L g6899 ( 
.A(n_6749),
.B(n_482),
.Y(n_6899)
);

AOI22xp33_ASAP7_75t_L g6900 ( 
.A1(n_6586),
.A2(n_486),
.B1(n_483),
.B2(n_485),
.Y(n_6900)
);

NOR2x1_ASAP7_75t_L g6901 ( 
.A(n_6584),
.B(n_486),
.Y(n_6901)
);

NAND4xp75_ASAP7_75t_L g6902 ( 
.A(n_6525),
.B(n_490),
.C(n_487),
.D(n_488),
.Y(n_6902)
);

INVx2_ASAP7_75t_L g6903 ( 
.A(n_6550),
.Y(n_6903)
);

NOR2xp33_ASAP7_75t_L g6904 ( 
.A(n_6578),
.B(n_488),
.Y(n_6904)
);

AND2x2_ASAP7_75t_L g6905 ( 
.A(n_6590),
.B(n_491),
.Y(n_6905)
);

OR2x2_ASAP7_75t_L g6906 ( 
.A(n_6542),
.B(n_491),
.Y(n_6906)
);

INVxp67_ASAP7_75t_SL g6907 ( 
.A(n_6650),
.Y(n_6907)
);

AOI33xp33_ASAP7_75t_L g6908 ( 
.A1(n_6735),
.A2(n_492),
.A3(n_493),
.B1(n_494),
.B2(n_496),
.B3(n_497),
.Y(n_6908)
);

NOR2xp33_ASAP7_75t_R g6909 ( 
.A(n_6591),
.B(n_492),
.Y(n_6909)
);

OAI221xp5_ASAP7_75t_SL g6910 ( 
.A1(n_6584),
.A2(n_6592),
.B1(n_6545),
.B2(n_6598),
.C(n_6751),
.Y(n_6910)
);

INVxp67_ASAP7_75t_L g6911 ( 
.A(n_6557),
.Y(n_6911)
);

OR2x2_ASAP7_75t_L g6912 ( 
.A(n_6692),
.B(n_493),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6680),
.Y(n_6913)
);

HB1xp67_ASAP7_75t_L g6914 ( 
.A(n_6698),
.Y(n_6914)
);

AOI22xp33_ASAP7_75t_L g6915 ( 
.A1(n_6738),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6683),
.Y(n_6916)
);

AOI22xp33_ASAP7_75t_L g6917 ( 
.A1(n_6746),
.A2(n_501),
.B1(n_498),
.B2(n_499),
.Y(n_6917)
);

BUFx3_ASAP7_75t_L g6918 ( 
.A(n_6594),
.Y(n_6918)
);

OAI22xp33_ASAP7_75t_L g6919 ( 
.A1(n_6592),
.A2(n_502),
.B1(n_498),
.B2(n_501),
.Y(n_6919)
);

AOI221x1_ASAP7_75t_L g6920 ( 
.A1(n_6653),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.C(n_507),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6572),
.Y(n_6921)
);

AOI22xp5_ASAP7_75t_L g6922 ( 
.A1(n_6751),
.A2(n_509),
.B1(n_505),
.B2(n_508),
.Y(n_6922)
);

AO21x2_ASAP7_75t_L g6923 ( 
.A1(n_6712),
.A2(n_510),
.B(n_513),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6684),
.Y(n_6924)
);

OR2x6_ASAP7_75t_L g6925 ( 
.A(n_6554),
.B(n_513),
.Y(n_6925)
);

INVx2_ASAP7_75t_SL g6926 ( 
.A(n_6659),
.Y(n_6926)
);

OAI31xp33_ASAP7_75t_L g6927 ( 
.A1(n_6653),
.A2(n_516),
.A3(n_514),
.B(n_515),
.Y(n_6927)
);

INVx1_ASAP7_75t_SL g6928 ( 
.A(n_6596),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6687),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6544),
.Y(n_6930)
);

INVx4_ASAP7_75t_L g6931 ( 
.A(n_6639),
.Y(n_6931)
);

OAI31xp33_ASAP7_75t_L g6932 ( 
.A1(n_6642),
.A2(n_517),
.A3(n_514),
.B(n_516),
.Y(n_6932)
);

INVx2_ASAP7_75t_SL g6933 ( 
.A(n_6659),
.Y(n_6933)
);

INVx2_ASAP7_75t_L g6934 ( 
.A(n_6551),
.Y(n_6934)
);

OAI22xp5_ASAP7_75t_L g6935 ( 
.A1(n_6545),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_6935)
);

AND2x2_ASAP7_75t_L g6936 ( 
.A(n_6754),
.B(n_6757),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6774),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6844),
.Y(n_6938)
);

INVx2_ASAP7_75t_L g6939 ( 
.A(n_6791),
.Y(n_6939)
);

HB1xp67_ASAP7_75t_L g6940 ( 
.A(n_6768),
.Y(n_6940)
);

AND2x2_ASAP7_75t_L g6941 ( 
.A(n_6755),
.B(n_6605),
.Y(n_6941)
);

AND2x4_ASAP7_75t_L g6942 ( 
.A(n_6886),
.B(n_6583),
.Y(n_6942)
);

INVxp67_ASAP7_75t_SL g6943 ( 
.A(n_6768),
.Y(n_6943)
);

HB1xp67_ASAP7_75t_L g6944 ( 
.A(n_6838),
.Y(n_6944)
);

CKINVDCx20_ASAP7_75t_R g6945 ( 
.A(n_6756),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6914),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_6840),
.B(n_6616),
.Y(n_6947)
);

OR2x2_ASAP7_75t_L g6948 ( 
.A(n_6835),
.B(n_6570),
.Y(n_6948)
);

NAND2xp5_ASAP7_75t_L g6949 ( 
.A(n_6767),
.B(n_6748),
.Y(n_6949)
);

NAND2xp5_ASAP7_75t_L g6950 ( 
.A(n_6827),
.B(n_6613),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6907),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6762),
.B(n_6585),
.Y(n_6952)
);

AND2x4_ASAP7_75t_SL g6953 ( 
.A(n_6931),
.B(n_6601),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6758),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6791),
.Y(n_6955)
);

OR2x2_ASAP7_75t_L g6956 ( 
.A(n_6847),
.B(n_6636),
.Y(n_6956)
);

OR2x2_ASAP7_75t_L g6957 ( 
.A(n_6928),
.B(n_6816),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6786),
.B(n_6671),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6821),
.B(n_6674),
.Y(n_6959)
);

BUFx2_ASAP7_75t_L g6960 ( 
.A(n_6759),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6766),
.Y(n_6961)
);

OR2x2_ASAP7_75t_L g6962 ( 
.A(n_6928),
.B(n_6829),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6773),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6760),
.B(n_6571),
.Y(n_6964)
);

OR2x2_ASAP7_75t_L g6965 ( 
.A(n_6839),
.B(n_6666),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6819),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6819),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6815),
.B(n_6647),
.Y(n_6968)
);

AND2x2_ASAP7_75t_L g6969 ( 
.A(n_6817),
.B(n_6793),
.Y(n_6969)
);

BUFx3_ASAP7_75t_L g6970 ( 
.A(n_6791),
.Y(n_6970)
);

INVx2_ASAP7_75t_L g6971 ( 
.A(n_6896),
.Y(n_6971)
);

NAND2x1_ASAP7_75t_L g6972 ( 
.A(n_6836),
.B(n_6697),
.Y(n_6972)
);

AND2x2_ASAP7_75t_L g6973 ( 
.A(n_6779),
.B(n_6651),
.Y(n_6973)
);

AND2x2_ASAP7_75t_L g6974 ( 
.A(n_6781),
.B(n_6704),
.Y(n_6974)
);

NAND2xp5_ASAP7_75t_SL g6975 ( 
.A(n_6785),
.B(n_6598),
.Y(n_6975)
);

INVx2_ASAP7_75t_L g6976 ( 
.A(n_6931),
.Y(n_6976)
);

AND2x4_ASAP7_75t_L g6977 ( 
.A(n_6836),
.B(n_6666),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6881),
.Y(n_6978)
);

OR2x2_ASAP7_75t_L g6979 ( 
.A(n_6854),
.B(n_6716),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6876),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_L g6981 ( 
.A(n_6827),
.B(n_6614),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6882),
.Y(n_6982)
);

BUFx2_ASAP7_75t_L g6983 ( 
.A(n_6925),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6923),
.Y(n_6984)
);

INVx3_ASAP7_75t_SL g6985 ( 
.A(n_6820),
.Y(n_6985)
);

NAND2xp5_ASAP7_75t_L g6986 ( 
.A(n_6809),
.B(n_6629),
.Y(n_6986)
);

OR2x2_ASAP7_75t_L g6987 ( 
.A(n_6812),
.B(n_6750),
.Y(n_6987)
);

NOR2x1_ASAP7_75t_SL g6988 ( 
.A(n_6925),
.B(n_6699),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6845),
.B(n_6736),
.Y(n_6989)
);

INVx2_ASAP7_75t_L g6990 ( 
.A(n_6850),
.Y(n_6990)
);

AND2x2_ASAP7_75t_L g6991 ( 
.A(n_6823),
.B(n_6706),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6923),
.Y(n_6992)
);

OR2x2_ASAP7_75t_L g6993 ( 
.A(n_6926),
.B(n_6611),
.Y(n_6993)
);

AND2x4_ASAP7_75t_L g6994 ( 
.A(n_6797),
.B(n_6631),
.Y(n_6994)
);

AND2x2_ASAP7_75t_L g6995 ( 
.A(n_6856),
.B(n_6708),
.Y(n_6995)
);

AND2x4_ASAP7_75t_L g6996 ( 
.A(n_6797),
.B(n_6803),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6850),
.Y(n_6997)
);

INVx2_ASAP7_75t_L g6998 ( 
.A(n_6918),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6888),
.B(n_6702),
.Y(n_6999)
);

OR2x2_ASAP7_75t_L g7000 ( 
.A(n_6933),
.B(n_6607),
.Y(n_7000)
);

INVx2_ASAP7_75t_L g7001 ( 
.A(n_6925),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6832),
.B(n_6658),
.Y(n_7002)
);

AND2x4_ASAP7_75t_L g7003 ( 
.A(n_6803),
.B(n_6638),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6776),
.Y(n_7004)
);

NAND2xp5_ASAP7_75t_L g7005 ( 
.A(n_6771),
.B(n_6643),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6843),
.B(n_6661),
.Y(n_7006)
);

NAND2xp5_ASAP7_75t_L g7007 ( 
.A(n_6764),
.B(n_6646),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6834),
.Y(n_7008)
);

NAND2x1p5_ASAP7_75t_L g7009 ( 
.A(n_6883),
.B(n_6655),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6841),
.Y(n_7010)
);

OR2x2_ASAP7_75t_L g7011 ( 
.A(n_6788),
.B(n_6593),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6852),
.Y(n_7012)
);

INVxp67_ASAP7_75t_SL g7013 ( 
.A(n_6883),
.Y(n_7013)
);

OAI221xp5_ASAP7_75t_L g7014 ( 
.A1(n_6753),
.A2(n_6642),
.B1(n_6597),
.B2(n_6603),
.C(n_6641),
.Y(n_7014)
);

OR2x2_ASAP7_75t_L g7015 ( 
.A(n_6837),
.B(n_6858),
.Y(n_7015)
);

BUFx2_ASAP7_75t_L g7016 ( 
.A(n_6909),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6842),
.B(n_6679),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6860),
.Y(n_7018)
);

AND2x2_ASAP7_75t_L g7019 ( 
.A(n_6870),
.B(n_6678),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6868),
.Y(n_7020)
);

INVx2_ASAP7_75t_SL g7021 ( 
.A(n_6878),
.Y(n_7021)
);

AND2x2_ASAP7_75t_L g7022 ( 
.A(n_6872),
.B(n_6682),
.Y(n_7022)
);

AND2x4_ASAP7_75t_L g7023 ( 
.A(n_6808),
.B(n_6649),
.Y(n_7023)
);

AND2x4_ASAP7_75t_L g7024 ( 
.A(n_6808),
.B(n_6804),
.Y(n_7024)
);

HB1xp67_ASAP7_75t_L g7025 ( 
.A(n_6884),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6930),
.Y(n_7026)
);

INVxp67_ASAP7_75t_L g7027 ( 
.A(n_6777),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6887),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6887),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6789),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6792),
.Y(n_7031)
);

AND2x4_ASAP7_75t_L g7032 ( 
.A(n_6806),
.B(n_6662),
.Y(n_7032)
);

OR2x2_ASAP7_75t_L g7033 ( 
.A(n_6848),
.B(n_6846),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6818),
.Y(n_7034)
);

HB1xp67_ASAP7_75t_L g7035 ( 
.A(n_6855),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_6826),
.Y(n_7036)
);

AND2x2_ASAP7_75t_L g7037 ( 
.A(n_6814),
.B(n_6624),
.Y(n_7037)
);

INVxp67_ASAP7_75t_SL g7038 ( 
.A(n_6799),
.Y(n_7038)
);

INVx2_ASAP7_75t_L g7039 ( 
.A(n_6873),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_L g7040 ( 
.A(n_6782),
.B(n_6663),
.Y(n_7040)
);

INVx2_ASAP7_75t_L g7041 ( 
.A(n_6905),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6934),
.Y(n_7042)
);

OR2x2_ASAP7_75t_L g7043 ( 
.A(n_6848),
.B(n_6588),
.Y(n_7043)
);

NOR2xp67_ASAP7_75t_L g7044 ( 
.A(n_6813),
.B(n_6703),
.Y(n_7044)
);

HB1xp67_ASAP7_75t_L g7045 ( 
.A(n_6810),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_6765),
.B(n_6626),
.Y(n_7046)
);

NOR3xp33_ASAP7_75t_L g7047 ( 
.A(n_6769),
.B(n_6597),
.C(n_6691),
.Y(n_7047)
);

AND2x4_ASAP7_75t_SL g7048 ( 
.A(n_6890),
.B(n_6610),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6889),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6898),
.Y(n_7050)
);

OR2x2_ASAP7_75t_L g7051 ( 
.A(n_6906),
.B(n_6589),
.Y(n_7051)
);

AND2x2_ASAP7_75t_L g7052 ( 
.A(n_6851),
.B(n_6620),
.Y(n_7052)
);

NAND3xp33_ASAP7_75t_L g7053 ( 
.A(n_6805),
.B(n_6894),
.C(n_6927),
.Y(n_7053)
);

AND2x2_ASAP7_75t_L g7054 ( 
.A(n_6795),
.B(n_6772),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_SL g7055 ( 
.A(n_6785),
.B(n_6622),
.Y(n_7055)
);

NOR2xp33_ASAP7_75t_L g7056 ( 
.A(n_6784),
.B(n_6581),
.Y(n_7056)
);

AND2x2_ASAP7_75t_L g7057 ( 
.A(n_6780),
.B(n_6660),
.Y(n_7057)
);

NAND2xp5_ASAP7_75t_L g7058 ( 
.A(n_6782),
.B(n_6664),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_6753),
.B(n_6693),
.Y(n_7059)
);

INVx2_ASAP7_75t_SL g7060 ( 
.A(n_6901),
.Y(n_7060)
);

NAND2xp5_ASAP7_75t_L g7061 ( 
.A(n_6770),
.B(n_6790),
.Y(n_7061)
);

OR2x2_ASAP7_75t_L g7062 ( 
.A(n_6775),
.B(n_6713),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6770),
.B(n_6667),
.Y(n_7063)
);

NAND2xp5_ASAP7_75t_L g7064 ( 
.A(n_6790),
.B(n_6552),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6913),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_6916),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6807),
.B(n_6553),
.Y(n_7067)
);

OR2x2_ASAP7_75t_L g7068 ( 
.A(n_6912),
.B(n_6714),
.Y(n_7068)
);

AND2x2_ASAP7_75t_L g7069 ( 
.A(n_6787),
.B(n_6627),
.Y(n_7069)
);

INVx2_ASAP7_75t_L g7070 ( 
.A(n_6892),
.Y(n_7070)
);

INVx2_ASAP7_75t_L g7071 ( 
.A(n_6897),
.Y(n_7071)
);

AND2x2_ASAP7_75t_L g7072 ( 
.A(n_6802),
.B(n_6637),
.Y(n_7072)
);

HB1xp67_ASAP7_75t_L g7073 ( 
.A(n_6783),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6924),
.Y(n_7074)
);

AND2x2_ASAP7_75t_L g7075 ( 
.A(n_6869),
.B(n_6644),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6929),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6880),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6885),
.Y(n_7078)
);

AND2x2_ASAP7_75t_L g7079 ( 
.A(n_6936),
.B(n_6893),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6940),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_7016),
.B(n_6801),
.Y(n_7081)
);

NOR2xp67_ASAP7_75t_L g7082 ( 
.A(n_7060),
.B(n_6813),
.Y(n_7082)
);

INVx2_ASAP7_75t_SL g7083 ( 
.A(n_6970),
.Y(n_7083)
);

AND2x2_ASAP7_75t_L g7084 ( 
.A(n_6960),
.B(n_6911),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6940),
.Y(n_7085)
);

OR2x2_ASAP7_75t_L g7086 ( 
.A(n_6948),
.B(n_6865),
.Y(n_7086)
);

OR2x2_ASAP7_75t_L g7087 ( 
.A(n_7045),
.B(n_6910),
.Y(n_7087)
);

NOR2xp67_ASAP7_75t_SL g7088 ( 
.A(n_7025),
.B(n_6874),
.Y(n_7088)
);

AND2x2_ASAP7_75t_L g7089 ( 
.A(n_6971),
.B(n_6985),
.Y(n_7089)
);

AND2x2_ASAP7_75t_L g7090 ( 
.A(n_6958),
.B(n_6903),
.Y(n_7090)
);

AND2x2_ASAP7_75t_L g7091 ( 
.A(n_6959),
.B(n_6921),
.Y(n_7091)
);

AND2x2_ASAP7_75t_L g7092 ( 
.A(n_6980),
.B(n_6859),
.Y(n_7092)
);

INVxp67_ASAP7_75t_SL g7093 ( 
.A(n_6988),
.Y(n_7093)
);

BUFx2_ASAP7_75t_L g7094 ( 
.A(n_6983),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6996),
.Y(n_7095)
);

OR2x2_ASAP7_75t_L g7096 ( 
.A(n_7035),
.B(n_6763),
.Y(n_7096)
);

AND2x4_ASAP7_75t_L g7097 ( 
.A(n_6996),
.B(n_6778),
.Y(n_7097)
);

OR2x2_ASAP7_75t_L g7098 ( 
.A(n_6938),
.B(n_6796),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_7027),
.B(n_6801),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_7027),
.B(n_6807),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_7024),
.B(n_6830),
.Y(n_7101)
);

NAND2xp67_ASAP7_75t_L g7102 ( 
.A(n_6939),
.B(n_6899),
.Y(n_7102)
);

INVx2_ASAP7_75t_L g7103 ( 
.A(n_6972),
.Y(n_7103)
);

NOR2xp33_ASAP7_75t_L g7104 ( 
.A(n_6945),
.B(n_6798),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6944),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6943),
.Y(n_7106)
);

AND2x2_ASAP7_75t_L g7107 ( 
.A(n_6969),
.B(n_6904),
.Y(n_7107)
);

INVx2_ASAP7_75t_L g7108 ( 
.A(n_7024),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6943),
.Y(n_7109)
);

AND2x4_ASAP7_75t_L g7110 ( 
.A(n_6942),
.B(n_6794),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_7073),
.Y(n_7111)
);

NAND2xp5_ASAP7_75t_L g7112 ( 
.A(n_6942),
.B(n_6761),
.Y(n_7112)
);

AND2x2_ASAP7_75t_L g7113 ( 
.A(n_7046),
.B(n_6953),
.Y(n_7113)
);

AND2x2_ASAP7_75t_L g7114 ( 
.A(n_6947),
.B(n_6863),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_7073),
.Y(n_7115)
);

INVx2_ASAP7_75t_L g7116 ( 
.A(n_7021),
.Y(n_7116)
);

AND2x2_ASAP7_75t_L g7117 ( 
.A(n_7057),
.B(n_6794),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6966),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6967),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_6951),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6937),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6946),
.Y(n_7122)
);

INVx2_ASAP7_75t_SL g7123 ( 
.A(n_6977),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_7013),
.Y(n_7124)
);

OR2x6_ASAP7_75t_L g7125 ( 
.A(n_7061),
.B(n_6874),
.Y(n_7125)
);

AND2x2_ASAP7_75t_L g7126 ( 
.A(n_6952),
.B(n_6866),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6994),
.Y(n_7127)
);

AND2x2_ASAP7_75t_L g7128 ( 
.A(n_6989),
.B(n_6861),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6994),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_6955),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_7013),
.Y(n_7131)
);

AND2x2_ASAP7_75t_L g7132 ( 
.A(n_7069),
.B(n_6862),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_L g7133 ( 
.A(n_7001),
.B(n_6932),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_7044),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_7044),
.Y(n_7135)
);

AND2x4_ASAP7_75t_L g7136 ( 
.A(n_7003),
.B(n_7023),
.Y(n_7136)
);

OR2x2_ASAP7_75t_L g7137 ( 
.A(n_7043),
.B(n_6864),
.Y(n_7137)
);

NOR2xp33_ASAP7_75t_L g7138 ( 
.A(n_7056),
.B(n_6784),
.Y(n_7138)
);

AND2x2_ASAP7_75t_SL g7139 ( 
.A(n_7061),
.B(n_6853),
.Y(n_7139)
);

OR2x6_ASAP7_75t_L g7140 ( 
.A(n_6976),
.B(n_6895),
.Y(n_7140)
);

NAND2xp5_ASAP7_75t_L g7141 ( 
.A(n_7038),
.B(n_6932),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6990),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6984),
.Y(n_7143)
);

OR2x2_ASAP7_75t_L g7144 ( 
.A(n_7063),
.B(n_7000),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_L g7145 ( 
.A(n_7038),
.B(n_6927),
.Y(n_7145)
);

INVx2_ASAP7_75t_L g7146 ( 
.A(n_6997),
.Y(n_7146)
);

OR2x2_ASAP7_75t_L g7147 ( 
.A(n_7063),
.B(n_6783),
.Y(n_7147)
);

INVx2_ASAP7_75t_SL g7148 ( 
.A(n_6977),
.Y(n_7148)
);

INVx1_ASAP7_75t_L g7149 ( 
.A(n_6992),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_7054),
.B(n_6922),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_7002),
.B(n_6862),
.Y(n_7151)
);

NOR2x1_ASAP7_75t_L g7152 ( 
.A(n_7053),
.B(n_6902),
.Y(n_7152)
);

INVx2_ASAP7_75t_L g7153 ( 
.A(n_7003),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_7028),
.Y(n_7154)
);

NOR2xp67_ASAP7_75t_L g7155 ( 
.A(n_7053),
.B(n_6833),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_6941),
.B(n_6645),
.Y(n_7156)
);

INVx1_ASAP7_75t_L g7157 ( 
.A(n_7029),
.Y(n_7157)
);

AND3x2_ASAP7_75t_L g7158 ( 
.A(n_7047),
.B(n_6877),
.C(n_6920),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_7072),
.B(n_6922),
.Y(n_7159)
);

NOR2x1_ASAP7_75t_L g7160 ( 
.A(n_6975),
.B(n_6867),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_6995),
.B(n_6720),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_6999),
.B(n_6730),
.Y(n_7162)
);

AND2x2_ASAP7_75t_L g7163 ( 
.A(n_6968),
.B(n_6734),
.Y(n_7163)
);

INVx2_ASAP7_75t_L g7164 ( 
.A(n_7023),
.Y(n_7164)
);

OR2x2_ASAP7_75t_L g7165 ( 
.A(n_6993),
.B(n_6825),
.Y(n_7165)
);

NAND2xp5_ASAP7_75t_L g7166 ( 
.A(n_7006),
.B(n_6919),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_7009),
.Y(n_7167)
);

AND2x2_ASAP7_75t_L g7168 ( 
.A(n_7037),
.B(n_6558),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_7068),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_6991),
.B(n_6935),
.Y(n_7170)
);

NAND2xp5_ASAP7_75t_L g7171 ( 
.A(n_6973),
.B(n_6800),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6964),
.B(n_6718),
.Y(n_7172)
);

AND2x2_ASAP7_75t_L g7173 ( 
.A(n_7052),
.B(n_6822),
.Y(n_7173)
);

AND2x2_ASAP7_75t_L g7174 ( 
.A(n_7048),
.B(n_6891),
.Y(n_7174)
);

AND2x2_ASAP7_75t_L g7175 ( 
.A(n_7075),
.B(n_6824),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_7017),
.B(n_6831),
.Y(n_7176)
);

NOR2xp33_ASAP7_75t_SL g7177 ( 
.A(n_7014),
.B(n_6879),
.Y(n_7177)
);

AND2x2_ASAP7_75t_L g7178 ( 
.A(n_7019),
.B(n_6811),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_7009),
.Y(n_7179)
);

NAND2xp5_ASAP7_75t_L g7180 ( 
.A(n_6998),
.B(n_6828),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_7040),
.Y(n_7181)
);

INVx1_ASAP7_75t_L g7182 ( 
.A(n_7040),
.Y(n_7182)
);

AND2x2_ASAP7_75t_L g7183 ( 
.A(n_7022),
.B(n_6701),
.Y(n_7183)
);

HB1xp67_ASAP7_75t_L g7184 ( 
.A(n_7011),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_7058),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_7058),
.Y(n_7186)
);

NAND2xp5_ASAP7_75t_L g7187 ( 
.A(n_7041),
.B(n_6871),
.Y(n_7187)
);

INVx1_ASAP7_75t_SL g7188 ( 
.A(n_6957),
.Y(n_7188)
);

INVx2_ASAP7_75t_L g7189 ( 
.A(n_6956),
.Y(n_7189)
);

INVx2_ASAP7_75t_SL g7190 ( 
.A(n_7032),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_7077),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6987),
.Y(n_7192)
);

INVxp67_ASAP7_75t_SL g7193 ( 
.A(n_6962),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_7078),
.Y(n_7194)
);

INVx2_ASAP7_75t_L g7195 ( 
.A(n_6974),
.Y(n_7195)
);

AND2x2_ASAP7_75t_L g7196 ( 
.A(n_7042),
.B(n_6877),
.Y(n_7196)
);

AND2x2_ASAP7_75t_L g7197 ( 
.A(n_7039),
.B(n_6849),
.Y(n_7197)
);

HB1xp67_ASAP7_75t_L g7198 ( 
.A(n_7051),
.Y(n_7198)
);

OR2x2_ASAP7_75t_L g7199 ( 
.A(n_7059),
.B(n_6857),
.Y(n_7199)
);

NAND2x1p5_ASAP7_75t_L g7200 ( 
.A(n_7070),
.B(n_6908),
.Y(n_7200)
);

OR2x6_ASAP7_75t_L g7201 ( 
.A(n_6950),
.B(n_6900),
.Y(n_7201)
);

INVx2_ASAP7_75t_L g7202 ( 
.A(n_7032),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_6986),
.Y(n_7203)
);

NAND2xp5_ASAP7_75t_L g7204 ( 
.A(n_7047),
.B(n_6875),
.Y(n_7204)
);

OR2x2_ASAP7_75t_L g7205 ( 
.A(n_7059),
.B(n_6915),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_7071),
.B(n_6917),
.Y(n_7206)
);

OAI21xp33_ASAP7_75t_L g7207 ( 
.A1(n_7067),
.A2(n_520),
.B(n_521),
.Y(n_7207)
);

HB1xp67_ASAP7_75t_L g7208 ( 
.A(n_6965),
.Y(n_7208)
);

OR2x2_ASAP7_75t_L g7209 ( 
.A(n_6950),
.B(n_521),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_7055),
.B(n_522),
.Y(n_7210)
);

INVx1_ASAP7_75t_SL g7211 ( 
.A(n_7015),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6986),
.Y(n_7212)
);

INVx3_ASAP7_75t_L g7213 ( 
.A(n_6954),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_6981),
.Y(n_7214)
);

AND2x2_ASAP7_75t_L g7215 ( 
.A(n_6961),
.B(n_524),
.Y(n_7215)
);

OR2x2_ASAP7_75t_L g7216 ( 
.A(n_6981),
.B(n_524),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_7136),
.B(n_7067),
.Y(n_7217)
);

CKINVDCx16_ASAP7_75t_R g7218 ( 
.A(n_7160),
.Y(n_7218)
);

NOR2xp33_ASAP7_75t_L g7219 ( 
.A(n_7207),
.B(n_7014),
.Y(n_7219)
);

AND2x2_ASAP7_75t_L g7220 ( 
.A(n_7126),
.B(n_6963),
.Y(n_7220)
);

AND2x2_ASAP7_75t_L g7221 ( 
.A(n_7089),
.B(n_7007),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_7080),
.Y(n_7222)
);

NAND2xp5_ASAP7_75t_L g7223 ( 
.A(n_7136),
.B(n_7158),
.Y(n_7223)
);

INVx2_ASAP7_75t_SL g7224 ( 
.A(n_7095),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_7080),
.Y(n_7225)
);

OAI21xp33_ASAP7_75t_SL g7226 ( 
.A1(n_7082),
.A2(n_7064),
.B(n_6949),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_7085),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_7108),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_7085),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_7094),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7198),
.Y(n_7231)
);

INVx3_ASAP7_75t_R g7232 ( 
.A(n_7097),
.Y(n_7232)
);

NOR2x1_ASAP7_75t_SL g7233 ( 
.A(n_7190),
.B(n_7064),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_7124),
.Y(n_7234)
);

AND2x2_ASAP7_75t_L g7235 ( 
.A(n_7113),
.B(n_7007),
.Y(n_7235)
);

AND2x2_ASAP7_75t_L g7236 ( 
.A(n_7116),
.B(n_7090),
.Y(n_7236)
);

INVxp33_ASAP7_75t_L g7237 ( 
.A(n_7104),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_7124),
.Y(n_7238)
);

NOR2x1p5_ASAP7_75t_L g7239 ( 
.A(n_7093),
.B(n_7005),
.Y(n_7239)
);

AND2x4_ASAP7_75t_L g7240 ( 
.A(n_7153),
.B(n_7004),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_7131),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_7110),
.B(n_7033),
.Y(n_7242)
);

INVx1_ASAP7_75t_SL g7243 ( 
.A(n_7110),
.Y(n_7243)
);

INVxp67_ASAP7_75t_L g7244 ( 
.A(n_7208),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_7131),
.Y(n_7245)
);

INVx2_ASAP7_75t_L g7246 ( 
.A(n_7164),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_7097),
.B(n_7005),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7127),
.B(n_6949),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7184),
.Y(n_7249)
);

INVx2_ASAP7_75t_L g7250 ( 
.A(n_7129),
.Y(n_7250)
);

OR2x2_ASAP7_75t_L g7251 ( 
.A(n_7096),
.B(n_6979),
.Y(n_7251)
);

INVx2_ASAP7_75t_SL g7252 ( 
.A(n_7123),
.Y(n_7252)
);

INVx2_ASAP7_75t_L g7253 ( 
.A(n_7148),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_L g7254 ( 
.A(n_7083),
.B(n_7008),
.Y(n_7254)
);

INVx3_ASAP7_75t_L g7255 ( 
.A(n_7202),
.Y(n_7255)
);

NOR2xp67_ASAP7_75t_SL g7256 ( 
.A(n_7105),
.B(n_7062),
.Y(n_7256)
);

OAI21xp33_ASAP7_75t_L g7257 ( 
.A1(n_7177),
.A2(n_7012),
.B(n_7010),
.Y(n_7257)
);

AND2x2_ASAP7_75t_L g7258 ( 
.A(n_7091),
.B(n_7018),
.Y(n_7258)
);

NOR2x1p5_ASAP7_75t_L g7259 ( 
.A(n_7193),
.B(n_7020),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_L g7260 ( 
.A(n_7178),
.B(n_7030),
.Y(n_7260)
);

INVx2_ASAP7_75t_L g7261 ( 
.A(n_7103),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7106),
.Y(n_7262)
);

OR2x6_ASAP7_75t_L g7263 ( 
.A(n_7210),
.B(n_7031),
.Y(n_7263)
);

AND2x2_ASAP7_75t_SL g7264 ( 
.A(n_7139),
.B(n_7034),
.Y(n_7264)
);

AND2x2_ASAP7_75t_SL g7265 ( 
.A(n_7145),
.B(n_7036),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7109),
.Y(n_7266)
);

NAND2xp5_ASAP7_75t_L g7267 ( 
.A(n_7175),
.B(n_7049),
.Y(n_7267)
);

INVx2_ASAP7_75t_L g7268 ( 
.A(n_7156),
.Y(n_7268)
);

OR2x2_ASAP7_75t_L g7269 ( 
.A(n_7144),
.B(n_7050),
.Y(n_7269)
);

NAND2xp5_ASAP7_75t_L g7270 ( 
.A(n_7117),
.B(n_7065),
.Y(n_7270)
);

INVx2_ASAP7_75t_SL g7271 ( 
.A(n_7079),
.Y(n_7271)
);

AND2x2_ASAP7_75t_L g7272 ( 
.A(n_7114),
.B(n_7066),
.Y(n_7272)
);

NOR2xp33_ASAP7_75t_L g7273 ( 
.A(n_7112),
.B(n_7074),
.Y(n_7273)
);

AND2x2_ASAP7_75t_L g7274 ( 
.A(n_7128),
.B(n_7084),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_7167),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_7167),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_7179),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_7179),
.Y(n_7278)
);

AND2x2_ASAP7_75t_L g7279 ( 
.A(n_7172),
.B(n_7076),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_7174),
.B(n_7026),
.Y(n_7280)
);

OAI31xp33_ASAP7_75t_SL g7281 ( 
.A1(n_7152),
.A2(n_6982),
.A3(n_6978),
.B(n_528),
.Y(n_7281)
);

NAND2xp5_ASAP7_75t_L g7282 ( 
.A(n_7155),
.B(n_526),
.Y(n_7282)
);

AND2x2_ASAP7_75t_L g7283 ( 
.A(n_7107),
.B(n_526),
.Y(n_7283)
);

NOR3xp33_ASAP7_75t_L g7284 ( 
.A(n_7138),
.B(n_527),
.C(n_528),
.Y(n_7284)
);

NOR2xp33_ASAP7_75t_L g7285 ( 
.A(n_7088),
.B(n_529),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_7154),
.Y(n_7286)
);

NAND4xp25_ASAP7_75t_SL g7287 ( 
.A(n_7204),
.B(n_7141),
.C(n_7100),
.D(n_7099),
.Y(n_7287)
);

INVx1_ASAP7_75t_L g7288 ( 
.A(n_7154),
.Y(n_7288)
);

INVx1_ASAP7_75t_SL g7289 ( 
.A(n_7134),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_L g7290 ( 
.A(n_7188),
.B(n_529),
.Y(n_7290)
);

INVx1_ASAP7_75t_L g7291 ( 
.A(n_7157),
.Y(n_7291)
);

OR2x2_ASAP7_75t_L g7292 ( 
.A(n_7086),
.B(n_530),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_7092),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7157),
.Y(n_7294)
);

NAND2xp5_ASAP7_75t_L g7295 ( 
.A(n_7196),
.B(n_530),
.Y(n_7295)
);

INVx2_ASAP7_75t_L g7296 ( 
.A(n_7195),
.Y(n_7296)
);

AND2x2_ASAP7_75t_L g7297 ( 
.A(n_7161),
.B(n_531),
.Y(n_7297)
);

INVxp67_ASAP7_75t_L g7298 ( 
.A(n_7098),
.Y(n_7298)
);

OR2x2_ASAP7_75t_L g7299 ( 
.A(n_7133),
.B(n_531),
.Y(n_7299)
);

NOR2x1_ASAP7_75t_L g7300 ( 
.A(n_7134),
.B(n_532),
.Y(n_7300)
);

OR2x6_ASAP7_75t_L g7301 ( 
.A(n_7209),
.B(n_533),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7143),
.Y(n_7302)
);

HB1xp67_ASAP7_75t_L g7303 ( 
.A(n_7135),
.Y(n_7303)
);

INVx2_ASAP7_75t_L g7304 ( 
.A(n_7130),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_7163),
.B(n_534),
.Y(n_7305)
);

BUFx2_ASAP7_75t_L g7306 ( 
.A(n_7135),
.Y(n_7306)
);

AOI322xp5_ASAP7_75t_L g7307 ( 
.A1(n_7081),
.A2(n_535),
.A3(n_537),
.B1(n_538),
.B2(n_539),
.C1(n_540),
.C2(n_542),
.Y(n_7307)
);

AOI22xp5_ASAP7_75t_L g7308 ( 
.A1(n_7201),
.A2(n_543),
.B1(n_537),
.B2(n_539),
.Y(n_7308)
);

OAI22xp5_ASAP7_75t_L g7309 ( 
.A1(n_7201),
.A2(n_7137),
.B1(n_7087),
.B2(n_7214),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_7173),
.B(n_543),
.Y(n_7310)
);

AND2x2_ASAP7_75t_L g7311 ( 
.A(n_7162),
.B(n_544),
.Y(n_7311)
);

OR2x2_ASAP7_75t_L g7312 ( 
.A(n_7165),
.B(n_544),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_7143),
.Y(n_7313)
);

AND2x2_ASAP7_75t_L g7314 ( 
.A(n_7211),
.B(n_545),
.Y(n_7314)
);

AND2x2_ASAP7_75t_L g7315 ( 
.A(n_7168),
.B(n_546),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_7149),
.Y(n_7316)
);

INVxp67_ASAP7_75t_SL g7317 ( 
.A(n_7213),
.Y(n_7317)
);

INVxp67_ASAP7_75t_SL g7318 ( 
.A(n_7213),
.Y(n_7318)
);

INVx2_ASAP7_75t_L g7319 ( 
.A(n_7183),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7197),
.B(n_547),
.Y(n_7320)
);

NOR2xp33_ASAP7_75t_L g7321 ( 
.A(n_7187),
.B(n_548),
.Y(n_7321)
);

OR2x2_ASAP7_75t_L g7322 ( 
.A(n_7171),
.B(n_7125),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_7149),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7111),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_7115),
.Y(n_7325)
);

AOI22xp33_ASAP7_75t_L g7326 ( 
.A1(n_7214),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_7326)
);

A2O1A1Ixp33_ASAP7_75t_L g7327 ( 
.A1(n_7203),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_7327)
);

AND2x2_ASAP7_75t_L g7328 ( 
.A(n_7192),
.B(n_7189),
.Y(n_7328)
);

AND2x2_ASAP7_75t_L g7329 ( 
.A(n_7176),
.B(n_553),
.Y(n_7329)
);

OR2x2_ASAP7_75t_L g7330 ( 
.A(n_7125),
.B(n_554),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_L g7331 ( 
.A(n_7151),
.B(n_555),
.Y(n_7331)
);

INVx2_ASAP7_75t_L g7332 ( 
.A(n_7142),
.Y(n_7332)
);

BUFx2_ASAP7_75t_L g7333 ( 
.A(n_7169),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_L g7334 ( 
.A(n_7102),
.B(n_556),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_L g7335 ( 
.A(n_7203),
.B(n_556),
.Y(n_7335)
);

AOI22xp5_ASAP7_75t_L g7336 ( 
.A1(n_7218),
.A2(n_7212),
.B1(n_7101),
.B2(n_7140),
.Y(n_7336)
);

NAND2xp5_ASAP7_75t_L g7337 ( 
.A(n_7243),
.B(n_7212),
.Y(n_7337)
);

OAI21xp33_ASAP7_75t_L g7338 ( 
.A1(n_7219),
.A2(n_7159),
.B(n_7180),
.Y(n_7338)
);

OAI21xp5_ASAP7_75t_L g7339 ( 
.A1(n_7226),
.A2(n_7199),
.B(n_7216),
.Y(n_7339)
);

AOI22xp33_ASAP7_75t_SL g7340 ( 
.A1(n_7264),
.A2(n_7182),
.B1(n_7185),
.B2(n_7181),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_7300),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7243),
.B(n_7146),
.Y(n_7342)
);

INVx2_ASAP7_75t_SL g7343 ( 
.A(n_7259),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_L g7344 ( 
.A(n_7274),
.B(n_7215),
.Y(n_7344)
);

INVx1_ASAP7_75t_L g7345 ( 
.A(n_7300),
.Y(n_7345)
);

O2A1O1Ixp33_ASAP7_75t_SL g7346 ( 
.A1(n_7307),
.A2(n_7147),
.B(n_7182),
.C(n_7181),
.Y(n_7346)
);

AOI22xp5_ASAP7_75t_L g7347 ( 
.A1(n_7287),
.A2(n_7140),
.B1(n_7186),
.B2(n_7185),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_7317),
.Y(n_7348)
);

NAND2x1p5_ASAP7_75t_L g7349 ( 
.A(n_7255),
.B(n_7120),
.Y(n_7349)
);

INVx2_ASAP7_75t_SL g7350 ( 
.A(n_7255),
.Y(n_7350)
);

AND2x2_ASAP7_75t_L g7351 ( 
.A(n_7236),
.B(n_7200),
.Y(n_7351)
);

HB1xp67_ASAP7_75t_L g7352 ( 
.A(n_7232),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7318),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_7303),
.Y(n_7354)
);

AOI21xp33_ASAP7_75t_L g7355 ( 
.A1(n_7226),
.A2(n_7205),
.B(n_7166),
.Y(n_7355)
);

AND2x4_ASAP7_75t_L g7356 ( 
.A(n_7252),
.B(n_7224),
.Y(n_7356)
);

AOI33xp33_ASAP7_75t_L g7357 ( 
.A1(n_7230),
.A2(n_7186),
.A3(n_7121),
.B1(n_7122),
.B2(n_7194),
.B3(n_7191),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_7306),
.Y(n_7358)
);

NAND2xp5_ASAP7_75t_L g7359 ( 
.A(n_7281),
.B(n_7132),
.Y(n_7359)
);

NAND2xp33_ASAP7_75t_SL g7360 ( 
.A(n_7256),
.B(n_7251),
.Y(n_7360)
);

AND2x2_ASAP7_75t_L g7361 ( 
.A(n_7235),
.B(n_7170),
.Y(n_7361)
);

AND2x2_ASAP7_75t_L g7362 ( 
.A(n_7221),
.B(n_7150),
.Y(n_7362)
);

AOI22xp5_ASAP7_75t_L g7363 ( 
.A1(n_7309),
.A2(n_7206),
.B1(n_7119),
.B2(n_7118),
.Y(n_7363)
);

INVxp67_ASAP7_75t_SL g7364 ( 
.A(n_7233),
.Y(n_7364)
);

INVx1_ASAP7_75t_SL g7365 ( 
.A(n_7265),
.Y(n_7365)
);

AND2x2_ASAP7_75t_L g7366 ( 
.A(n_7253),
.B(n_557),
.Y(n_7366)
);

INVx1_ASAP7_75t_SL g7367 ( 
.A(n_7333),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_7222),
.Y(n_7368)
);

AOI22xp5_ASAP7_75t_L g7369 ( 
.A1(n_7309),
.A2(n_558),
.B1(n_559),
.B2(n_560),
.Y(n_7369)
);

NAND2xp5_ASAP7_75t_L g7370 ( 
.A(n_7281),
.B(n_561),
.Y(n_7370)
);

OR2x2_ASAP7_75t_L g7371 ( 
.A(n_7242),
.B(n_561),
.Y(n_7371)
);

XNOR2xp5_ASAP7_75t_L g7372 ( 
.A(n_7239),
.B(n_562),
.Y(n_7372)
);

INVx1_ASAP7_75t_L g7373 ( 
.A(n_7225),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_L g7374 ( 
.A(n_7271),
.B(n_563),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_7227),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_7229),
.Y(n_7376)
);

AND2x2_ASAP7_75t_L g7377 ( 
.A(n_7279),
.B(n_563),
.Y(n_7377)
);

OR2x2_ASAP7_75t_L g7378 ( 
.A(n_7247),
.B(n_568),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_7231),
.B(n_569),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_7234),
.Y(n_7380)
);

AOI32xp33_ASAP7_75t_L g7381 ( 
.A1(n_7285),
.A2(n_569),
.A3(n_570),
.B1(n_571),
.B2(n_572),
.Y(n_7381)
);

INVx1_ASAP7_75t_L g7382 ( 
.A(n_7249),
.Y(n_7382)
);

OR2x2_ASAP7_75t_L g7383 ( 
.A(n_7223),
.B(n_570),
.Y(n_7383)
);

INVx2_ASAP7_75t_L g7384 ( 
.A(n_7228),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_7238),
.Y(n_7385)
);

INVx2_ASAP7_75t_SL g7386 ( 
.A(n_7240),
.Y(n_7386)
);

AND2x4_ASAP7_75t_L g7387 ( 
.A(n_7240),
.B(n_571),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_7241),
.Y(n_7388)
);

AND2x2_ASAP7_75t_L g7389 ( 
.A(n_7220),
.B(n_572),
.Y(n_7389)
);

OR2x2_ASAP7_75t_L g7390 ( 
.A(n_7322),
.B(n_573),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_7245),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_7246),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_7283),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7305),
.Y(n_7394)
);

INVx1_ASAP7_75t_SL g7395 ( 
.A(n_7330),
.Y(n_7395)
);

NOR2xp67_ASAP7_75t_L g7396 ( 
.A(n_7244),
.B(n_573),
.Y(n_7396)
);

NAND2xp5_ASAP7_75t_L g7397 ( 
.A(n_7329),
.B(n_574),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_7311),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_7315),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_7314),
.Y(n_7400)
);

AND2x4_ASAP7_75t_L g7401 ( 
.A(n_7261),
.B(n_575),
.Y(n_7401)
);

INVx2_ASAP7_75t_L g7402 ( 
.A(n_7250),
.Y(n_7402)
);

AOI32xp33_ASAP7_75t_L g7403 ( 
.A1(n_7282),
.A2(n_575),
.A3(n_576),
.B1(n_577),
.B2(n_579),
.Y(n_7403)
);

AOI31xp33_ASAP7_75t_L g7404 ( 
.A1(n_7237),
.A2(n_576),
.A3(n_580),
.B(n_581),
.Y(n_7404)
);

OAI21xp33_ASAP7_75t_L g7405 ( 
.A1(n_7217),
.A2(n_580),
.B(n_582),
.Y(n_7405)
);

AND2x2_ASAP7_75t_L g7406 ( 
.A(n_7280),
.B(n_582),
.Y(n_7406)
);

HB1xp67_ASAP7_75t_L g7407 ( 
.A(n_7301),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_7297),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_7258),
.Y(n_7409)
);

NAND2xp5_ASAP7_75t_L g7410 ( 
.A(n_7298),
.B(n_583),
.Y(n_7410)
);

AND2x4_ASAP7_75t_L g7411 ( 
.A(n_7268),
.B(n_583),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_7286),
.Y(n_7412)
);

INVx2_ASAP7_75t_L g7413 ( 
.A(n_7319),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_7288),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7289),
.Y(n_7415)
);

NAND2xp67_ASAP7_75t_SL g7416 ( 
.A(n_7272),
.B(n_7328),
.Y(n_7416)
);

AOI22xp5_ASAP7_75t_L g7417 ( 
.A1(n_7257),
.A2(n_584),
.B1(n_585),
.B2(n_586),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_7293),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_L g7419 ( 
.A(n_7308),
.B(n_584),
.Y(n_7419)
);

NAND3xp33_ASAP7_75t_L g7420 ( 
.A(n_7257),
.B(n_587),
.C(n_588),
.Y(n_7420)
);

NAND2x1_ASAP7_75t_L g7421 ( 
.A(n_7301),
.B(n_588),
.Y(n_7421)
);

NOR2xp33_ASAP7_75t_L g7422 ( 
.A(n_7292),
.B(n_589),
.Y(n_7422)
);

OAI22xp5_ASAP7_75t_L g7423 ( 
.A1(n_7308),
.A2(n_589),
.B1(n_590),
.B2(n_591),
.Y(n_7423)
);

AOI22xp33_ASAP7_75t_L g7424 ( 
.A1(n_7355),
.A2(n_7263),
.B1(n_7273),
.B2(n_7248),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_7341),
.Y(n_7425)
);

AND2x2_ASAP7_75t_L g7426 ( 
.A(n_7352),
.B(n_7296),
.Y(n_7426)
);

NOR2xp33_ASAP7_75t_L g7427 ( 
.A(n_7359),
.B(n_7312),
.Y(n_7427)
);

HB1xp67_ASAP7_75t_L g7428 ( 
.A(n_7345),
.Y(n_7428)
);

HB1xp67_ASAP7_75t_L g7429 ( 
.A(n_7396),
.Y(n_7429)
);

NAND2xp5_ASAP7_75t_L g7430 ( 
.A(n_7364),
.B(n_7289),
.Y(n_7430)
);

AOI22x1_ASAP7_75t_L g7431 ( 
.A1(n_7367),
.A2(n_7269),
.B1(n_7304),
.B2(n_7332),
.Y(n_7431)
);

NAND2xp33_ASAP7_75t_L g7432 ( 
.A(n_7365),
.B(n_7284),
.Y(n_7432)
);

NAND2xp5_ASAP7_75t_L g7433 ( 
.A(n_7386),
.B(n_7307),
.Y(n_7433)
);

NOR2xp33_ASAP7_75t_L g7434 ( 
.A(n_7407),
.B(n_7295),
.Y(n_7434)
);

NOR2xp33_ASAP7_75t_L g7435 ( 
.A(n_7370),
.B(n_7299),
.Y(n_7435)
);

NAND2x1_ASAP7_75t_L g7436 ( 
.A(n_7356),
.B(n_7262),
.Y(n_7436)
);

INVx2_ASAP7_75t_L g7437 ( 
.A(n_7349),
.Y(n_7437)
);

NAND2xp5_ASAP7_75t_L g7438 ( 
.A(n_7356),
.B(n_7321),
.Y(n_7438)
);

NAND2xp5_ASAP7_75t_L g7439 ( 
.A(n_7350),
.B(n_7275),
.Y(n_7439)
);

AND2x4_ASAP7_75t_L g7440 ( 
.A(n_7358),
.B(n_7276),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_7421),
.Y(n_7441)
);

NAND2xp33_ASAP7_75t_L g7442 ( 
.A(n_7343),
.B(n_7267),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_7415),
.Y(n_7443)
);

OR2x2_ASAP7_75t_L g7444 ( 
.A(n_7342),
.B(n_7260),
.Y(n_7444)
);

INVx1_ASAP7_75t_SL g7445 ( 
.A(n_7360),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_7415),
.Y(n_7446)
);

AND2x2_ASAP7_75t_L g7447 ( 
.A(n_7351),
.B(n_7263),
.Y(n_7447)
);

AND2x2_ASAP7_75t_L g7448 ( 
.A(n_7362),
.B(n_7263),
.Y(n_7448)
);

NAND2xp5_ASAP7_75t_L g7449 ( 
.A(n_7361),
.B(n_7277),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_7406),
.Y(n_7450)
);

NAND3xp33_ASAP7_75t_SL g7451 ( 
.A(n_7339),
.B(n_7270),
.C(n_7320),
.Y(n_7451)
);

INVx1_ASAP7_75t_SL g7452 ( 
.A(n_7337),
.Y(n_7452)
);

INVx1_ASAP7_75t_SL g7453 ( 
.A(n_7387),
.Y(n_7453)
);

AND2x4_ASAP7_75t_L g7454 ( 
.A(n_7354),
.B(n_7278),
.Y(n_7454)
);

INVx2_ASAP7_75t_L g7455 ( 
.A(n_7387),
.Y(n_7455)
);

INVx3_ASAP7_75t_L g7456 ( 
.A(n_7401),
.Y(n_7456)
);

AND4x1_ASAP7_75t_L g7457 ( 
.A(n_7336),
.B(n_7310),
.C(n_7290),
.D(n_7326),
.Y(n_7457)
);

INVxp67_ASAP7_75t_L g7458 ( 
.A(n_7344),
.Y(n_7458)
);

OAI22xp33_ASAP7_75t_L g7459 ( 
.A1(n_7347),
.A2(n_7334),
.B1(n_7301),
.B2(n_7254),
.Y(n_7459)
);

AOI22xp33_ASAP7_75t_L g7460 ( 
.A1(n_7338),
.A2(n_7266),
.B1(n_7325),
.B2(n_7324),
.Y(n_7460)
);

HB1xp67_ASAP7_75t_L g7461 ( 
.A(n_7372),
.Y(n_7461)
);

CKINVDCx16_ASAP7_75t_R g7462 ( 
.A(n_7363),
.Y(n_7462)
);

INVx2_ASAP7_75t_SL g7463 ( 
.A(n_7411),
.Y(n_7463)
);

NAND2xp5_ASAP7_75t_L g7464 ( 
.A(n_7348),
.B(n_7327),
.Y(n_7464)
);

INVx1_ASAP7_75t_SL g7465 ( 
.A(n_7377),
.Y(n_7465)
);

NOR2x1_ASAP7_75t_L g7466 ( 
.A(n_7416),
.B(n_7291),
.Y(n_7466)
);

INVx1_ASAP7_75t_SL g7467 ( 
.A(n_7389),
.Y(n_7467)
);

INVxp67_ASAP7_75t_L g7468 ( 
.A(n_7422),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7353),
.Y(n_7469)
);

NAND2xp5_ASAP7_75t_L g7470 ( 
.A(n_7409),
.B(n_7331),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_7366),
.Y(n_7471)
);

NAND2xp5_ASAP7_75t_L g7472 ( 
.A(n_7340),
.B(n_7294),
.Y(n_7472)
);

INVx1_ASAP7_75t_L g7473 ( 
.A(n_7411),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7395),
.B(n_7335),
.Y(n_7474)
);

INVx1_ASAP7_75t_SL g7475 ( 
.A(n_7401),
.Y(n_7475)
);

OR2x2_ASAP7_75t_L g7476 ( 
.A(n_7383),
.B(n_7335),
.Y(n_7476)
);

NOR2x1_ASAP7_75t_L g7477 ( 
.A(n_7420),
.B(n_7302),
.Y(n_7477)
);

NOR2xp33_ASAP7_75t_L g7478 ( 
.A(n_7405),
.B(n_7313),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_7390),
.Y(n_7479)
);

INVx1_ASAP7_75t_SL g7480 ( 
.A(n_7371),
.Y(n_7480)
);

BUFx2_ASAP7_75t_L g7481 ( 
.A(n_7393),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7357),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_7418),
.Y(n_7483)
);

BUFx3_ASAP7_75t_L g7484 ( 
.A(n_7394),
.Y(n_7484)
);

NAND2xp5_ASAP7_75t_L g7485 ( 
.A(n_7400),
.B(n_7316),
.Y(n_7485)
);

AND2x2_ASAP7_75t_L g7486 ( 
.A(n_7398),
.B(n_7323),
.Y(n_7486)
);

OR2x2_ASAP7_75t_L g7487 ( 
.A(n_7378),
.B(n_590),
.Y(n_7487)
);

AND2x2_ASAP7_75t_L g7488 ( 
.A(n_7399),
.B(n_591),
.Y(n_7488)
);

NAND2xp5_ASAP7_75t_L g7489 ( 
.A(n_7408),
.B(n_592),
.Y(n_7489)
);

BUFx3_ASAP7_75t_L g7490 ( 
.A(n_7384),
.Y(n_7490)
);

AND2x2_ASAP7_75t_L g7491 ( 
.A(n_7413),
.B(n_597),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_7369),
.B(n_597),
.Y(n_7492)
);

INVx1_ASAP7_75t_SL g7493 ( 
.A(n_7374),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7397),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7410),
.Y(n_7495)
);

AOI21xp5_ASAP7_75t_L g7496 ( 
.A1(n_7346),
.A2(n_598),
.B(n_599),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7379),
.Y(n_7497)
);

AND2x2_ASAP7_75t_L g7498 ( 
.A(n_7392),
.B(n_598),
.Y(n_7498)
);

OAI22xp5_ASAP7_75t_L g7499 ( 
.A1(n_7417),
.A2(n_599),
.B1(n_600),
.B2(n_601),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7402),
.B(n_600),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7429),
.Y(n_7501)
);

INVx2_ASAP7_75t_SL g7502 ( 
.A(n_7436),
.Y(n_7502)
);

AOI22xp5_ASAP7_75t_L g7503 ( 
.A1(n_7462),
.A2(n_7382),
.B1(n_7373),
.B2(n_7375),
.Y(n_7503)
);

AOI21xp5_ASAP7_75t_L g7504 ( 
.A1(n_7496),
.A2(n_7419),
.B(n_7404),
.Y(n_7504)
);

NAND2xp5_ASAP7_75t_L g7505 ( 
.A(n_7445),
.B(n_7403),
.Y(n_7505)
);

AOI22xp33_ASAP7_75t_SL g7506 ( 
.A1(n_7445),
.A2(n_7368),
.B1(n_7376),
.B2(n_7385),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_7456),
.Y(n_7507)
);

AOI22xp5_ASAP7_75t_L g7508 ( 
.A1(n_7427),
.A2(n_7391),
.B1(n_7388),
.B2(n_7423),
.Y(n_7508)
);

AOI222xp33_ASAP7_75t_L g7509 ( 
.A1(n_7472),
.A2(n_7380),
.B1(n_7414),
.B2(n_7412),
.C1(n_7381),
.C2(n_607),
.Y(n_7509)
);

AOI21xp5_ASAP7_75t_L g7510 ( 
.A1(n_7442),
.A2(n_7380),
.B(n_602),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7430),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7456),
.Y(n_7512)
);

CKINVDCx14_ASAP7_75t_R g7513 ( 
.A(n_7447),
.Y(n_7513)
);

NAND2x1_ASAP7_75t_L g7514 ( 
.A(n_7441),
.B(n_603),
.Y(n_7514)
);

NAND2xp5_ASAP7_75t_L g7515 ( 
.A(n_7453),
.B(n_603),
.Y(n_7515)
);

OAI21xp5_ASAP7_75t_L g7516 ( 
.A1(n_7466),
.A2(n_7424),
.B(n_7433),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7428),
.Y(n_7517)
);

OAI22xp5_ASAP7_75t_L g7518 ( 
.A1(n_7482),
.A2(n_604),
.B1(n_605),
.B2(n_607),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7426),
.Y(n_7519)
);

OAI22xp5_ASAP7_75t_L g7520 ( 
.A1(n_7460),
.A2(n_604),
.B1(n_605),
.B2(n_608),
.Y(n_7520)
);

INVx1_ASAP7_75t_SL g7521 ( 
.A(n_7453),
.Y(n_7521)
);

OAI22xp5_ASAP7_75t_SL g7522 ( 
.A1(n_7465),
.A2(n_608),
.B1(n_609),
.B2(n_610),
.Y(n_7522)
);

AOI21xp33_ASAP7_75t_SL g7523 ( 
.A1(n_7463),
.A2(n_7431),
.B(n_7473),
.Y(n_7523)
);

INVx2_ASAP7_75t_L g7524 ( 
.A(n_7455),
.Y(n_7524)
);

NOR2xp33_ASAP7_75t_L g7525 ( 
.A(n_7475),
.B(n_611),
.Y(n_7525)
);

AND2x4_ASAP7_75t_L g7526 ( 
.A(n_7475),
.B(n_611),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7481),
.Y(n_7527)
);

INVx3_ASAP7_75t_L g7528 ( 
.A(n_7440),
.Y(n_7528)
);

INVx1_ASAP7_75t_SL g7529 ( 
.A(n_7448),
.Y(n_7529)
);

OAI21xp33_ASAP7_75t_L g7530 ( 
.A1(n_7434),
.A2(n_612),
.B(n_613),
.Y(n_7530)
);

OR2x2_ASAP7_75t_L g7531 ( 
.A(n_7452),
.B(n_613),
.Y(n_7531)
);

AND2x2_ASAP7_75t_L g7532 ( 
.A(n_7465),
.B(n_614),
.Y(n_7532)
);

NOR2x1_ASAP7_75t_L g7533 ( 
.A(n_7452),
.B(n_614),
.Y(n_7533)
);

INVx1_ASAP7_75t_L g7534 ( 
.A(n_7440),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_7461),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_7467),
.B(n_615),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7449),
.Y(n_7537)
);

INVx1_ASAP7_75t_SL g7538 ( 
.A(n_7467),
.Y(n_7538)
);

AOI221xp5_ASAP7_75t_L g7539 ( 
.A1(n_7459),
.A2(n_7451),
.B1(n_7432),
.B2(n_7478),
.C(n_7446),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_7488),
.Y(n_7540)
);

INVxp67_ASAP7_75t_L g7541 ( 
.A(n_7435),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7484),
.Y(n_7542)
);

AOI22xp5_ASAP7_75t_L g7543 ( 
.A1(n_7458),
.A2(n_616),
.B1(n_617),
.B2(n_618),
.Y(n_7543)
);

NOR2x1_ASAP7_75t_L g7544 ( 
.A(n_7490),
.B(n_617),
.Y(n_7544)
);

NAND3xp33_ASAP7_75t_L g7545 ( 
.A(n_7457),
.B(n_7437),
.C(n_7443),
.Y(n_7545)
);

AOI222xp33_ASAP7_75t_L g7546 ( 
.A1(n_7425),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.C1(n_622),
.C2(n_624),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_7454),
.Y(n_7547)
);

OAI22xp5_ASAP7_75t_L g7548 ( 
.A1(n_7444),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7439),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7454),
.Y(n_7550)
);

NAND2xp5_ASAP7_75t_L g7551 ( 
.A(n_7450),
.B(n_622),
.Y(n_7551)
);

AND2x2_ASAP7_75t_L g7552 ( 
.A(n_7479),
.B(n_625),
.Y(n_7552)
);

AND2x2_ASAP7_75t_L g7553 ( 
.A(n_7471),
.B(n_625),
.Y(n_7553)
);

AND2x2_ASAP7_75t_L g7554 ( 
.A(n_7480),
.B(n_626),
.Y(n_7554)
);

OAI221xp5_ASAP7_75t_L g7555 ( 
.A1(n_7464),
.A2(n_627),
.B1(n_629),
.B2(n_632),
.C(n_633),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7486),
.Y(n_7556)
);

AOI22xp33_ASAP7_75t_L g7557 ( 
.A1(n_7477),
.A2(n_7494),
.B1(n_7483),
.B2(n_7495),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7491),
.Y(n_7558)
);

AOI22xp33_ASAP7_75t_SL g7559 ( 
.A1(n_7480),
.A2(n_632),
.B1(n_633),
.B2(n_634),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7487),
.Y(n_7560)
);

NAND2x1p5_ASAP7_75t_L g7561 ( 
.A(n_7498),
.B(n_634),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_7474),
.Y(n_7562)
);

NAND2xp5_ASAP7_75t_L g7563 ( 
.A(n_7500),
.B(n_7469),
.Y(n_7563)
);

AND2x2_ASAP7_75t_L g7564 ( 
.A(n_7493),
.B(n_7438),
.Y(n_7564)
);

NAND2xp5_ASAP7_75t_L g7565 ( 
.A(n_7502),
.B(n_7499),
.Y(n_7565)
);

OAI22xp5_ASAP7_75t_L g7566 ( 
.A1(n_7513),
.A2(n_7476),
.B1(n_7468),
.B2(n_7492),
.Y(n_7566)
);

NAND2xp5_ASAP7_75t_L g7567 ( 
.A(n_7528),
.B(n_7497),
.Y(n_7567)
);

AND2x2_ASAP7_75t_L g7568 ( 
.A(n_7521),
.B(n_7470),
.Y(n_7568)
);

NOR2xp33_ASAP7_75t_L g7569 ( 
.A(n_7529),
.B(n_7489),
.Y(n_7569)
);

NAND2xp5_ASAP7_75t_L g7570 ( 
.A(n_7528),
.B(n_7485),
.Y(n_7570)
);

AOI22xp5_ASAP7_75t_L g7571 ( 
.A1(n_7538),
.A2(n_635),
.B1(n_636),
.B2(n_637),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7533),
.Y(n_7572)
);

NAND2xp5_ASAP7_75t_L g7573 ( 
.A(n_7526),
.B(n_635),
.Y(n_7573)
);

AOI22xp5_ASAP7_75t_L g7574 ( 
.A1(n_7542),
.A2(n_638),
.B1(n_639),
.B2(n_640),
.Y(n_7574)
);

HB1xp67_ASAP7_75t_L g7575 ( 
.A(n_7533),
.Y(n_7575)
);

OAI22xp33_ASAP7_75t_L g7576 ( 
.A1(n_7527),
.A2(n_638),
.B1(n_639),
.B2(n_641),
.Y(n_7576)
);

AOI221xp5_ASAP7_75t_L g7577 ( 
.A1(n_7516),
.A2(n_641),
.B1(n_642),
.B2(n_644),
.C(n_646),
.Y(n_7577)
);

HB1xp67_ASAP7_75t_L g7578 ( 
.A(n_7544),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7544),
.Y(n_7579)
);

NOR2xp33_ASAP7_75t_L g7580 ( 
.A(n_7547),
.B(n_644),
.Y(n_7580)
);

NAND2xp33_ASAP7_75t_SL g7581 ( 
.A(n_7514),
.B(n_646),
.Y(n_7581)
);

AND2x2_ASAP7_75t_L g7582 ( 
.A(n_7524),
.B(n_647),
.Y(n_7582)
);

NAND2xp5_ASAP7_75t_L g7583 ( 
.A(n_7526),
.B(n_648),
.Y(n_7583)
);

NAND2xp5_ASAP7_75t_L g7584 ( 
.A(n_7550),
.B(n_648),
.Y(n_7584)
);

INVx1_ASAP7_75t_SL g7585 ( 
.A(n_7532),
.Y(n_7585)
);

AOI31xp33_ASAP7_75t_L g7586 ( 
.A1(n_7523),
.A2(n_7534),
.A3(n_7539),
.B(n_7506),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_7536),
.Y(n_7587)
);

NAND3xp33_ASAP7_75t_SL g7588 ( 
.A(n_7523),
.B(n_7509),
.C(n_7503),
.Y(n_7588)
);

OAI22xp5_ASAP7_75t_L g7589 ( 
.A1(n_7545),
.A2(n_649),
.B1(n_650),
.B2(n_651),
.Y(n_7589)
);

OAI21xp5_ASAP7_75t_L g7590 ( 
.A1(n_7504),
.A2(n_649),
.B(n_651),
.Y(n_7590)
);

AOI21xp5_ASAP7_75t_SL g7591 ( 
.A1(n_7531),
.A2(n_652),
.B(n_653),
.Y(n_7591)
);

NAND3xp33_ASAP7_75t_L g7592 ( 
.A(n_7546),
.B(n_653),
.C(n_654),
.Y(n_7592)
);

AOI21xp33_ASAP7_75t_L g7593 ( 
.A1(n_7512),
.A2(n_654),
.B(n_655),
.Y(n_7593)
);

NOR2xp33_ASAP7_75t_L g7594 ( 
.A(n_7507),
.B(n_656),
.Y(n_7594)
);

XOR2x2_ASAP7_75t_L g7595 ( 
.A(n_7505),
.B(n_657),
.Y(n_7595)
);

NAND2xp5_ASAP7_75t_L g7596 ( 
.A(n_7519),
.B(n_657),
.Y(n_7596)
);

AOI31xp33_ASAP7_75t_L g7597 ( 
.A1(n_7561),
.A2(n_658),
.A3(n_659),
.B(n_660),
.Y(n_7597)
);

OA21x2_ASAP7_75t_L g7598 ( 
.A1(n_7510),
.A2(n_7515),
.B(n_7501),
.Y(n_7598)
);

INVx1_ASAP7_75t_L g7599 ( 
.A(n_7522),
.Y(n_7599)
);

INVx2_ASAP7_75t_SL g7600 ( 
.A(n_7554),
.Y(n_7600)
);

AOI32xp33_ASAP7_75t_L g7601 ( 
.A1(n_7535),
.A2(n_658),
.A3(n_659),
.B1(n_660),
.B2(n_661),
.Y(n_7601)
);

AOI21xp5_ASAP7_75t_L g7602 ( 
.A1(n_7525),
.A2(n_662),
.B(n_663),
.Y(n_7602)
);

AND2x2_ASAP7_75t_L g7603 ( 
.A(n_7564),
.B(n_7540),
.Y(n_7603)
);

NAND2xp5_ASAP7_75t_L g7604 ( 
.A(n_7559),
.B(n_663),
.Y(n_7604)
);

AND2x2_ASAP7_75t_L g7605 ( 
.A(n_7556),
.B(n_664),
.Y(n_7605)
);

AOI21xp5_ASAP7_75t_L g7606 ( 
.A1(n_7563),
.A2(n_664),
.B(n_665),
.Y(n_7606)
);

OAI22xp5_ASAP7_75t_L g7607 ( 
.A1(n_7557),
.A2(n_666),
.B1(n_667),
.B2(n_668),
.Y(n_7607)
);

NAND2xp5_ASAP7_75t_L g7608 ( 
.A(n_7552),
.B(n_666),
.Y(n_7608)
);

OAI22xp5_ASAP7_75t_L g7609 ( 
.A1(n_7508),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.Y(n_7609)
);

OAI221xp5_ASAP7_75t_L g7610 ( 
.A1(n_7517),
.A2(n_669),
.B1(n_670),
.B2(n_671),
.C(n_673),
.Y(n_7610)
);

AOI221xp5_ASAP7_75t_L g7611 ( 
.A1(n_7518),
.A2(n_671),
.B1(n_673),
.B2(n_674),
.C(n_675),
.Y(n_7611)
);

AOI21xp33_ASAP7_75t_L g7612 ( 
.A1(n_7511),
.A2(n_675),
.B(n_677),
.Y(n_7612)
);

NOR2xp33_ASAP7_75t_L g7613 ( 
.A(n_7597),
.B(n_7530),
.Y(n_7613)
);

AND2x2_ASAP7_75t_L g7614 ( 
.A(n_7603),
.B(n_7553),
.Y(n_7614)
);

OR2x6_ASAP7_75t_L g7615 ( 
.A(n_7591),
.B(n_7541),
.Y(n_7615)
);

AND2x2_ASAP7_75t_L g7616 ( 
.A(n_7568),
.B(n_7560),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_7575),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_7572),
.Y(n_7618)
);

AND2x2_ASAP7_75t_L g7619 ( 
.A(n_7585),
.B(n_7558),
.Y(n_7619)
);

AOI22xp5_ASAP7_75t_L g7620 ( 
.A1(n_7588),
.A2(n_7520),
.B1(n_7562),
.B2(n_7537),
.Y(n_7620)
);

AND2x2_ASAP7_75t_L g7621 ( 
.A(n_7600),
.B(n_7549),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7578),
.Y(n_7622)
);

AND2x2_ASAP7_75t_L g7623 ( 
.A(n_7599),
.B(n_7587),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_7579),
.Y(n_7624)
);

AOI21xp5_ASAP7_75t_L g7625 ( 
.A1(n_7581),
.A2(n_7551),
.B(n_7555),
.Y(n_7625)
);

NAND2xp5_ASAP7_75t_L g7626 ( 
.A(n_7582),
.B(n_7548),
.Y(n_7626)
);

OAI22xp5_ASAP7_75t_L g7627 ( 
.A1(n_7586),
.A2(n_7543),
.B1(n_678),
.B2(n_680),
.Y(n_7627)
);

NOR2xp67_ASAP7_75t_SL g7628 ( 
.A(n_7570),
.B(n_677),
.Y(n_7628)
);

NOR2xp33_ASAP7_75t_L g7629 ( 
.A(n_7592),
.B(n_681),
.Y(n_7629)
);

OR2x2_ASAP7_75t_L g7630 ( 
.A(n_7584),
.B(n_682),
.Y(n_7630)
);

NAND2xp5_ASAP7_75t_L g7631 ( 
.A(n_7605),
.B(n_682),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_7573),
.Y(n_7632)
);

NAND2xp5_ASAP7_75t_L g7633 ( 
.A(n_7580),
.B(n_683),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_L g7634 ( 
.A(n_7601),
.B(n_683),
.Y(n_7634)
);

NAND2x1p5_ASAP7_75t_L g7635 ( 
.A(n_7598),
.B(n_684),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7583),
.Y(n_7636)
);

NOR2xp33_ASAP7_75t_L g7637 ( 
.A(n_7592),
.B(n_684),
.Y(n_7637)
);

AND2x2_ASAP7_75t_L g7638 ( 
.A(n_7598),
.B(n_685),
.Y(n_7638)
);

NAND2xp5_ASAP7_75t_L g7639 ( 
.A(n_7594),
.B(n_685),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7608),
.Y(n_7640)
);

AND2x2_ASAP7_75t_L g7641 ( 
.A(n_7590),
.B(n_686),
.Y(n_7641)
);

NAND2xp33_ASAP7_75t_L g7642 ( 
.A(n_7567),
.B(n_687),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7569),
.B(n_687),
.Y(n_7643)
);

INVx1_ASAP7_75t_L g7644 ( 
.A(n_7635),
.Y(n_7644)
);

NAND4xp75_ASAP7_75t_L g7645 ( 
.A(n_7638),
.B(n_7616),
.C(n_7617),
.D(n_7623),
.Y(n_7645)
);

AOI221xp5_ASAP7_75t_SL g7646 ( 
.A1(n_7627),
.A2(n_7566),
.B1(n_7589),
.B2(n_7565),
.C(n_7607),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_7615),
.Y(n_7647)
);

NAND3xp33_ASAP7_75t_L g7648 ( 
.A(n_7628),
.B(n_7577),
.C(n_7606),
.Y(n_7648)
);

NOR2xp33_ASAP7_75t_L g7649 ( 
.A(n_7615),
.B(n_7604),
.Y(n_7649)
);

OAI221xp5_ASAP7_75t_L g7650 ( 
.A1(n_7620),
.A2(n_7596),
.B1(n_7609),
.B2(n_7611),
.C(n_7595),
.Y(n_7650)
);

NAND3xp33_ASAP7_75t_L g7651 ( 
.A(n_7642),
.B(n_7620),
.C(n_7637),
.Y(n_7651)
);

OAI21xp33_ASAP7_75t_L g7652 ( 
.A1(n_7613),
.A2(n_7571),
.B(n_7602),
.Y(n_7652)
);

AOI21xp5_ASAP7_75t_L g7653 ( 
.A1(n_7615),
.A2(n_7625),
.B(n_7622),
.Y(n_7653)
);

AOI21xp5_ASAP7_75t_L g7654 ( 
.A1(n_7627),
.A2(n_7612),
.B(n_7593),
.Y(n_7654)
);

NOR2xp33_ASAP7_75t_SL g7655 ( 
.A(n_7614),
.B(n_7621),
.Y(n_7655)
);

NAND4xp25_ASAP7_75t_L g7656 ( 
.A(n_7619),
.B(n_7610),
.C(n_7574),
.D(n_7576),
.Y(n_7656)
);

NOR3xp33_ASAP7_75t_L g7657 ( 
.A(n_7634),
.B(n_688),
.C(n_689),
.Y(n_7657)
);

INVx2_ASAP7_75t_L g7658 ( 
.A(n_7618),
.Y(n_7658)
);

NAND2xp5_ASAP7_75t_SL g7659 ( 
.A(n_7624),
.B(n_688),
.Y(n_7659)
);

NAND2xp5_ASAP7_75t_L g7660 ( 
.A(n_7643),
.B(n_689),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_7631),
.B(n_691),
.Y(n_7661)
);

INVxp67_ASAP7_75t_SL g7662 ( 
.A(n_7629),
.Y(n_7662)
);

NOR2xp67_ASAP7_75t_L g7663 ( 
.A(n_7626),
.B(n_691),
.Y(n_7663)
);

OAI21xp33_ASAP7_75t_SL g7664 ( 
.A1(n_7641),
.A2(n_692),
.B(n_693),
.Y(n_7664)
);

NAND4xp25_ASAP7_75t_L g7665 ( 
.A(n_7640),
.B(n_7636),
.C(n_7632),
.D(n_7633),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7630),
.Y(n_7666)
);

NAND3xp33_ASAP7_75t_L g7667 ( 
.A(n_7639),
.B(n_692),
.C(n_693),
.Y(n_7667)
);

AOI322xp5_ASAP7_75t_L g7668 ( 
.A1(n_7613),
.A2(n_694),
.A3(n_695),
.B1(n_696),
.B2(n_698),
.C1(n_699),
.C2(n_702),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_7635),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_7635),
.Y(n_7670)
);

AOI21xp5_ASAP7_75t_L g7671 ( 
.A1(n_7642),
.A2(n_695),
.B(n_696),
.Y(n_7671)
);

NAND3xp33_ASAP7_75t_L g7672 ( 
.A(n_7655),
.B(n_698),
.C(n_699),
.Y(n_7672)
);

NAND2xp5_ASAP7_75t_L g7673 ( 
.A(n_7663),
.B(n_703),
.Y(n_7673)
);

AND4x1_ASAP7_75t_L g7674 ( 
.A(n_7653),
.B(n_703),
.C(n_704),
.D(n_705),
.Y(n_7674)
);

INVx1_ASAP7_75t_L g7675 ( 
.A(n_7660),
.Y(n_7675)
);

OAI21xp33_ASAP7_75t_L g7676 ( 
.A1(n_7652),
.A2(n_706),
.B(n_1713),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7645),
.Y(n_7677)
);

O2A1O1Ixp33_ASAP7_75t_L g7678 ( 
.A1(n_7664),
.A2(n_2144),
.B(n_2184),
.C(n_2226),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7644),
.B(n_7669),
.Y(n_7679)
);

AOI21xp5_ASAP7_75t_L g7680 ( 
.A1(n_7647),
.A2(n_2012),
.B(n_2031),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7670),
.Y(n_7681)
);

NAND2xp5_ASAP7_75t_L g7682 ( 
.A(n_7649),
.B(n_1995),
.Y(n_7682)
);

NAND2xp5_ASAP7_75t_SL g7683 ( 
.A(n_7658),
.B(n_2012),
.Y(n_7683)
);

XNOR2x2_ASAP7_75t_L g7684 ( 
.A(n_7651),
.B(n_2012),
.Y(n_7684)
);

NAND4xp25_ASAP7_75t_L g7685 ( 
.A(n_7646),
.B(n_2144),
.C(n_2184),
.D(n_2226),
.Y(n_7685)
);

OR2x2_ASAP7_75t_L g7686 ( 
.A(n_7656),
.B(n_2184),
.Y(n_7686)
);

AND2x2_ASAP7_75t_L g7687 ( 
.A(n_7662),
.B(n_2031),
.Y(n_7687)
);

NOR3xp33_ASAP7_75t_L g7688 ( 
.A(n_7650),
.B(n_2226),
.C(n_2391),
.Y(n_7688)
);

NAND2xp33_ASAP7_75t_SL g7689 ( 
.A(n_7659),
.B(n_2481),
.Y(n_7689)
);

INVx1_ASAP7_75t_SL g7690 ( 
.A(n_7671),
.Y(n_7690)
);

NOR3xp33_ASAP7_75t_L g7691 ( 
.A(n_7665),
.B(n_2226),
.C(n_2391),
.Y(n_7691)
);

INVx2_ASAP7_75t_SL g7692 ( 
.A(n_7666),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_7667),
.Y(n_7693)
);

NAND5xp2_ASAP7_75t_L g7694 ( 
.A(n_7654),
.B(n_1882),
.C(n_1933),
.D(n_2017),
.E(n_2012),
.Y(n_7694)
);

NAND2xp5_ASAP7_75t_SL g7695 ( 
.A(n_7648),
.B(n_2022),
.Y(n_7695)
);

NAND2xp5_ASAP7_75t_L g7696 ( 
.A(n_7661),
.B(n_2022),
.Y(n_7696)
);

NAND2xp5_ASAP7_75t_L g7697 ( 
.A(n_7668),
.B(n_2022),
.Y(n_7697)
);

AND2x2_ASAP7_75t_L g7698 ( 
.A(n_7657),
.B(n_2022),
.Y(n_7698)
);

AOI211xp5_ASAP7_75t_L g7699 ( 
.A1(n_7650),
.A2(n_2481),
.B(n_2480),
.C(n_2479),
.Y(n_7699)
);

NAND3xp33_ASAP7_75t_L g7700 ( 
.A(n_7655),
.B(n_2022),
.C(n_2031),
.Y(n_7700)
);

INVx2_ASAP7_75t_L g7701 ( 
.A(n_7645),
.Y(n_7701)
);

AND2x2_ASAP7_75t_L g7702 ( 
.A(n_7658),
.B(n_2031),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7660),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7674),
.Y(n_7704)
);

NOR2xp33_ASAP7_75t_L g7705 ( 
.A(n_7674),
.B(n_2031),
.Y(n_7705)
);

AOI32xp33_ASAP7_75t_L g7706 ( 
.A1(n_7677),
.A2(n_2017),
.A3(n_1995),
.B1(n_2004),
.B2(n_2012),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7673),
.Y(n_7707)
);

AOI21xp5_ASAP7_75t_L g7708 ( 
.A1(n_7679),
.A2(n_2017),
.B(n_2004),
.Y(n_7708)
);

AND2x4_ASAP7_75t_L g7709 ( 
.A(n_7681),
.B(n_7692),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_7701),
.B(n_2017),
.Y(n_7710)
);

NAND3xp33_ASAP7_75t_SL g7711 ( 
.A(n_7690),
.B(n_1882),
.C(n_1933),
.Y(n_7711)
);

NOR4xp25_ASAP7_75t_L g7712 ( 
.A(n_7676),
.B(n_7693),
.C(n_7703),
.D(n_7675),
.Y(n_7712)
);

NAND2xp5_ASAP7_75t_SL g7713 ( 
.A(n_7672),
.B(n_1995),
.Y(n_7713)
);

NAND4xp75_ASAP7_75t_L g7714 ( 
.A(n_7697),
.B(n_2004),
.C(n_2017),
.D(n_1882),
.Y(n_7714)
);

OAI21xp5_ASAP7_75t_SL g7715 ( 
.A1(n_7686),
.A2(n_2481),
.B(n_2480),
.Y(n_7715)
);

INVx1_ASAP7_75t_L g7716 ( 
.A(n_7687),
.Y(n_7716)
);

NOR2xp33_ASAP7_75t_L g7717 ( 
.A(n_7685),
.B(n_2004),
.Y(n_7717)
);

NAND3xp33_ASAP7_75t_L g7718 ( 
.A(n_7699),
.B(n_2004),
.C(n_1882),
.Y(n_7718)
);

OAI21xp5_ASAP7_75t_L g7719 ( 
.A1(n_7678),
.A2(n_1882),
.B(n_1933),
.Y(n_7719)
);

NOR3x1_ASAP7_75t_L g7720 ( 
.A(n_7700),
.B(n_1933),
.C(n_1943),
.Y(n_7720)
);

A2O1A1Ixp33_ASAP7_75t_L g7721 ( 
.A1(n_7689),
.A2(n_1933),
.B(n_2480),
.C(n_2479),
.Y(n_7721)
);

NOR2xp33_ASAP7_75t_L g7722 ( 
.A(n_7696),
.B(n_1992),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_7698),
.Y(n_7723)
);

OAI322xp33_ASAP7_75t_L g7724 ( 
.A1(n_7695),
.A2(n_2481),
.A3(n_2480),
.B1(n_2479),
.B2(n_2470),
.C1(n_2469),
.C2(n_2460),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_7702),
.Y(n_7725)
);

NAND2xp5_ASAP7_75t_SL g7726 ( 
.A(n_7688),
.B(n_2481),
.Y(n_7726)
);

NAND2xp5_ASAP7_75t_L g7727 ( 
.A(n_7691),
.B(n_1992),
.Y(n_7727)
);

NOR2x1_ASAP7_75t_L g7728 ( 
.A(n_7694),
.B(n_2481),
.Y(n_7728)
);

NAND2xp5_ASAP7_75t_L g7729 ( 
.A(n_7682),
.B(n_1988),
.Y(n_7729)
);

NOR2xp33_ASAP7_75t_L g7730 ( 
.A(n_7683),
.B(n_7684),
.Y(n_7730)
);

NOR2x1_ASAP7_75t_L g7731 ( 
.A(n_7680),
.B(n_2480),
.Y(n_7731)
);

NOR2xp33_ASAP7_75t_SL g7732 ( 
.A(n_7672),
.B(n_1935),
.Y(n_7732)
);

NOR2xp33_ASAP7_75t_SL g7733 ( 
.A(n_7672),
.B(n_1935),
.Y(n_7733)
);

NAND2xp5_ASAP7_75t_SL g7734 ( 
.A(n_7674),
.B(n_2480),
.Y(n_7734)
);

NAND2xp5_ASAP7_75t_L g7735 ( 
.A(n_7674),
.B(n_1956),
.Y(n_7735)
);

XNOR2x1_ASAP7_75t_L g7736 ( 
.A(n_7709),
.B(n_2479),
.Y(n_7736)
);

NAND4xp25_ASAP7_75t_SL g7737 ( 
.A(n_7704),
.B(n_2470),
.C(n_2469),
.D(n_2460),
.Y(n_7737)
);

OAI211xp5_ASAP7_75t_L g7738 ( 
.A1(n_7712),
.A2(n_7728),
.B(n_7715),
.C(n_7734),
.Y(n_7738)
);

OAI211xp5_ASAP7_75t_SL g7739 ( 
.A1(n_7707),
.A2(n_7723),
.B(n_7713),
.C(n_7725),
.Y(n_7739)
);

NAND2xp5_ASAP7_75t_L g7740 ( 
.A(n_7709),
.B(n_1956),
.Y(n_7740)
);

AOI321xp33_ASAP7_75t_L g7741 ( 
.A1(n_7716),
.A2(n_2479),
.A3(n_2470),
.B1(n_2469),
.B2(n_2460),
.C(n_2435),
.Y(n_7741)
);

OR3x1_ASAP7_75t_L g7742 ( 
.A(n_7711),
.B(n_2479),
.C(n_2470),
.Y(n_7742)
);

OAI211xp5_ASAP7_75t_SL g7743 ( 
.A1(n_7710),
.A2(n_1800),
.B(n_1782),
.C(n_1777),
.Y(n_7743)
);

AOI21xp5_ASAP7_75t_L g7744 ( 
.A1(n_7735),
.A2(n_1800),
.B(n_1782),
.Y(n_7744)
);

AND2x2_ASAP7_75t_L g7745 ( 
.A(n_7705),
.B(n_1992),
.Y(n_7745)
);

NAND4xp25_ASAP7_75t_L g7746 ( 
.A(n_7732),
.B(n_2391),
.C(n_2228),
.D(n_2354),
.Y(n_7746)
);

NAND2xp5_ASAP7_75t_L g7747 ( 
.A(n_7733),
.B(n_1950),
.Y(n_7747)
);

NOR3xp33_ASAP7_75t_L g7748 ( 
.A(n_7714),
.B(n_2206),
.C(n_2228),
.Y(n_7748)
);

OAI221xp5_ASAP7_75t_L g7749 ( 
.A1(n_7721),
.A2(n_7719),
.B1(n_7730),
.B2(n_7706),
.C(n_7718),
.Y(n_7749)
);

NOR3xp33_ASAP7_75t_L g7750 ( 
.A(n_7722),
.B(n_2206),
.C(n_2228),
.Y(n_7750)
);

AOI211x1_ASAP7_75t_L g7751 ( 
.A1(n_7726),
.A2(n_1992),
.B(n_1943),
.C(n_1950),
.Y(n_7751)
);

NAND4xp25_ASAP7_75t_SL g7752 ( 
.A(n_7731),
.B(n_2469),
.C(n_2460),
.D(n_2435),
.Y(n_7752)
);

NAND3xp33_ASAP7_75t_L g7753 ( 
.A(n_7717),
.B(n_2470),
.C(n_2469),
.Y(n_7753)
);

AOI211xp5_ASAP7_75t_L g7754 ( 
.A1(n_7724),
.A2(n_2470),
.B(n_2469),
.C(n_2460),
.Y(n_7754)
);

OAI21xp5_ASAP7_75t_L g7755 ( 
.A1(n_7708),
.A2(n_1800),
.B(n_1782),
.Y(n_7755)
);

NAND4xp25_ASAP7_75t_L g7756 ( 
.A(n_7720),
.B(n_2354),
.C(n_2391),
.D(n_2206),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7727),
.B(n_1988),
.Y(n_7757)
);

NAND4xp25_ASAP7_75t_SL g7758 ( 
.A(n_7729),
.B(n_2435),
.C(n_2432),
.D(n_2428),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7709),
.Y(n_7759)
);

NOR2xp33_ASAP7_75t_R g7760 ( 
.A(n_7704),
.B(n_2460),
.Y(n_7760)
);

NOR4xp75_ASAP7_75t_L g7761 ( 
.A(n_7713),
.B(n_2435),
.C(n_2432),
.D(n_2428),
.Y(n_7761)
);

NAND5xp2_ASAP7_75t_L g7762 ( 
.A(n_7704),
.B(n_1777),
.C(n_1782),
.D(n_1800),
.E(n_2432),
.Y(n_7762)
);

NAND2xp5_ASAP7_75t_L g7763 ( 
.A(n_7709),
.B(n_1956),
.Y(n_7763)
);

NOR3xp33_ASAP7_75t_L g7764 ( 
.A(n_7704),
.B(n_2354),
.C(n_1800),
.Y(n_7764)
);

NOR2xp33_ASAP7_75t_L g7765 ( 
.A(n_7759),
.B(n_1956),
.Y(n_7765)
);

NOR2xp33_ASAP7_75t_R g7766 ( 
.A(n_7752),
.B(n_2435),
.Y(n_7766)
);

AOI221xp5_ASAP7_75t_L g7767 ( 
.A1(n_7749),
.A2(n_2432),
.B1(n_2435),
.B2(n_2213),
.C(n_2208),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7736),
.Y(n_7768)
);

OAI211xp5_ASAP7_75t_SL g7769 ( 
.A1(n_7738),
.A2(n_1782),
.B(n_1777),
.C(n_1740),
.Y(n_7769)
);

NAND2x1_ASAP7_75t_SL g7770 ( 
.A(n_7745),
.B(n_2432),
.Y(n_7770)
);

INVxp67_ASAP7_75t_L g7771 ( 
.A(n_7762),
.Y(n_7771)
);

BUFx6f_ASAP7_75t_L g7772 ( 
.A(n_7740),
.Y(n_7772)
);

NOR2x1p5_ASAP7_75t_L g7773 ( 
.A(n_7756),
.B(n_2213),
.Y(n_7773)
);

CKINVDCx20_ASAP7_75t_R g7774 ( 
.A(n_7760),
.Y(n_7774)
);

NOR2xp33_ASAP7_75t_R g7775 ( 
.A(n_7758),
.B(n_1777),
.Y(n_7775)
);

NOR2xp33_ASAP7_75t_R g7776 ( 
.A(n_7737),
.B(n_1777),
.Y(n_7776)
);

NAND2x1p5_ASAP7_75t_L g7777 ( 
.A(n_7763),
.B(n_7747),
.Y(n_7777)
);

CKINVDCx16_ASAP7_75t_R g7778 ( 
.A(n_7755),
.Y(n_7778)
);

AOI22xp5_ASAP7_75t_L g7779 ( 
.A1(n_7739),
.A2(n_2213),
.B1(n_2208),
.B2(n_2203),
.Y(n_7779)
);

NOR2x1p5_ASAP7_75t_L g7780 ( 
.A(n_7746),
.B(n_2213),
.Y(n_7780)
);

NAND4xp75_ASAP7_75t_L g7781 ( 
.A(n_7751),
.B(n_2213),
.C(n_2208),
.D(n_2203),
.Y(n_7781)
);

NAND2xp5_ASAP7_75t_L g7782 ( 
.A(n_7750),
.B(n_1956),
.Y(n_7782)
);

OAI221xp5_ASAP7_75t_L g7783 ( 
.A1(n_7741),
.A2(n_2213),
.B1(n_2208),
.B2(n_2203),
.C(n_2179),
.Y(n_7783)
);

NOR2x1_ASAP7_75t_L g7784 ( 
.A(n_7769),
.B(n_7742),
.Y(n_7784)
);

INVxp67_ASAP7_75t_L g7785 ( 
.A(n_7765),
.Y(n_7785)
);

XNOR2xp5_ASAP7_75t_L g7786 ( 
.A(n_7774),
.B(n_7761),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_7770),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7768),
.Y(n_7788)
);

XNOR2xp5_ASAP7_75t_L g7789 ( 
.A(n_7773),
.B(n_7753),
.Y(n_7789)
);

AOI22xp5_ASAP7_75t_L g7790 ( 
.A1(n_7771),
.A2(n_7764),
.B1(n_7743),
.B2(n_7754),
.Y(n_7790)
);

NOR2xp33_ASAP7_75t_SL g7791 ( 
.A(n_7783),
.B(n_7744),
.Y(n_7791)
);

NOR2x1_ASAP7_75t_L g7792 ( 
.A(n_7781),
.B(n_7757),
.Y(n_7792)
);

NOR2x1_ASAP7_75t_L g7793 ( 
.A(n_7780),
.B(n_7782),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7777),
.Y(n_7794)
);

NAND4xp75_ASAP7_75t_L g7795 ( 
.A(n_7779),
.B(n_7748),
.C(n_2208),
.D(n_2203),
.Y(n_7795)
);

AND2x4_ASAP7_75t_L g7796 ( 
.A(n_7772),
.B(n_7778),
.Y(n_7796)
);

AND2x4_ASAP7_75t_L g7797 ( 
.A(n_7772),
.B(n_7766),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7772),
.Y(n_7798)
);

NOR2x1_ASAP7_75t_L g7799 ( 
.A(n_7776),
.B(n_2208),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_7775),
.Y(n_7800)
);

INVx1_ASAP7_75t_L g7801 ( 
.A(n_7786),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_7798),
.Y(n_7802)
);

NOR2x1_ASAP7_75t_L g7803 ( 
.A(n_7787),
.B(n_7767),
.Y(n_7803)
);

AND4x1_ASAP7_75t_L g7804 ( 
.A(n_7788),
.B(n_1950),
.C(n_1992),
.D(n_1988),
.Y(n_7804)
);

OR3x2_ASAP7_75t_L g7805 ( 
.A(n_7794),
.B(n_1943),
.C(n_1988),
.Y(n_7805)
);

OAI211xp5_ASAP7_75t_SL g7806 ( 
.A1(n_7790),
.A2(n_1721),
.B(n_1740),
.C(n_1742),
.Y(n_7806)
);

AO211x2_ASAP7_75t_L g7807 ( 
.A1(n_7800),
.A2(n_2203),
.B(n_2179),
.C(n_2169),
.Y(n_7807)
);

AND4x1_ASAP7_75t_L g7808 ( 
.A(n_7793),
.B(n_1943),
.C(n_1988),
.D(n_1950),
.Y(n_7808)
);

NAND3xp33_ASAP7_75t_L g7809 ( 
.A(n_7791),
.B(n_2203),
.C(n_2179),
.Y(n_7809)
);

NAND2xp5_ASAP7_75t_L g7810 ( 
.A(n_7796),
.B(n_1935),
.Y(n_7810)
);

NOR3xp33_ASAP7_75t_L g7811 ( 
.A(n_7785),
.B(n_1742),
.C(n_1721),
.Y(n_7811)
);

NAND2xp5_ASAP7_75t_L g7812 ( 
.A(n_7797),
.B(n_1935),
.Y(n_7812)
);

INVxp67_ASAP7_75t_L g7813 ( 
.A(n_7784),
.Y(n_7813)
);

NOR3xp33_ASAP7_75t_SL g7814 ( 
.A(n_7789),
.B(n_1935),
.C(n_1950),
.Y(n_7814)
);

NAND2xp5_ASAP7_75t_SL g7815 ( 
.A(n_7792),
.B(n_7799),
.Y(n_7815)
);

NOR2x1_ASAP7_75t_L g7816 ( 
.A(n_7795),
.B(n_2179),
.Y(n_7816)
);

NAND5xp2_ASAP7_75t_L g7817 ( 
.A(n_7788),
.B(n_1742),
.C(n_1740),
.D(n_1721),
.E(n_1943),
.Y(n_7817)
);

OA22x2_ASAP7_75t_L g7818 ( 
.A1(n_7790),
.A2(n_2179),
.B1(n_2169),
.B2(n_2133),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_7786),
.Y(n_7819)
);

CKINVDCx5p33_ASAP7_75t_R g7820 ( 
.A(n_7802),
.Y(n_7820)
);

HB1xp67_ASAP7_75t_L g7821 ( 
.A(n_7813),
.Y(n_7821)
);

HB1xp67_ASAP7_75t_L g7822 ( 
.A(n_7801),
.Y(n_7822)
);

BUFx12f_ASAP7_75t_L g7823 ( 
.A(n_7819),
.Y(n_7823)
);

INVx1_ASAP7_75t_SL g7824 ( 
.A(n_7803),
.Y(n_7824)
);

CKINVDCx5p33_ASAP7_75t_R g7825 ( 
.A(n_7815),
.Y(n_7825)
);

OR2x2_ASAP7_75t_L g7826 ( 
.A(n_7817),
.B(n_2179),
.Y(n_7826)
);

NAND2xp33_ASAP7_75t_R g7827 ( 
.A(n_7814),
.B(n_2169),
.Y(n_7827)
);

BUFx2_ASAP7_75t_L g7828 ( 
.A(n_7816),
.Y(n_7828)
);

AND2x2_ASAP7_75t_L g7829 ( 
.A(n_7810),
.B(n_7812),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7818),
.Y(n_7830)
);

AOI21xp5_ASAP7_75t_L g7831 ( 
.A1(n_7806),
.A2(n_1742),
.B(n_1740),
.Y(n_7831)
);

AND2x4_ASAP7_75t_L g7832 ( 
.A(n_7809),
.B(n_2169),
.Y(n_7832)
);

INVx2_ASAP7_75t_L g7833 ( 
.A(n_7805),
.Y(n_7833)
);

CKINVDCx5p33_ASAP7_75t_R g7834 ( 
.A(n_7804),
.Y(n_7834)
);

CKINVDCx5p33_ASAP7_75t_R g7835 ( 
.A(n_7808),
.Y(n_7835)
);

INVx2_ASAP7_75t_L g7836 ( 
.A(n_7807),
.Y(n_7836)
);

CKINVDCx5p33_ASAP7_75t_R g7837 ( 
.A(n_7811),
.Y(n_7837)
);

AOI322xp5_ASAP7_75t_L g7838 ( 
.A1(n_7824),
.A2(n_2169),
.A3(n_2133),
.B1(n_2121),
.B2(n_2112),
.C1(n_2093),
.C2(n_2097),
.Y(n_7838)
);

INVx1_ASAP7_75t_SL g7839 ( 
.A(n_7821),
.Y(n_7839)
);

AOI221xp5_ASAP7_75t_L g7840 ( 
.A1(n_7822),
.A2(n_2056),
.B1(n_2133),
.B2(n_2121),
.C(n_2112),
.Y(n_7840)
);

OAI221xp5_ASAP7_75t_L g7841 ( 
.A1(n_7820),
.A2(n_2169),
.B1(n_2133),
.B2(n_2121),
.C(n_2112),
.Y(n_7841)
);

AOI322xp5_ASAP7_75t_L g7842 ( 
.A1(n_7823),
.A2(n_2133),
.A3(n_2121),
.B1(n_2112),
.B2(n_2104),
.C1(n_2093),
.C2(n_2056),
.Y(n_7842)
);

XOR2x2_ASAP7_75t_L g7843 ( 
.A(n_7826),
.B(n_1740),
.Y(n_7843)
);

OAI221xp5_ASAP7_75t_L g7844 ( 
.A1(n_7825),
.A2(n_2133),
.B1(n_2121),
.B2(n_2112),
.C(n_2104),
.Y(n_7844)
);

BUFx2_ASAP7_75t_L g7845 ( 
.A(n_7836),
.Y(n_7845)
);

NAND2xp5_ASAP7_75t_L g7846 ( 
.A(n_7835),
.B(n_1721),
.Y(n_7846)
);

AND2x4_ASAP7_75t_L g7847 ( 
.A(n_7830),
.B(n_2121),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7832),
.Y(n_7848)
);

HB1xp67_ASAP7_75t_L g7849 ( 
.A(n_7827),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_7845),
.Y(n_7850)
);

AOI22xp5_ASAP7_75t_L g7851 ( 
.A1(n_7839),
.A2(n_7834),
.B1(n_7837),
.B2(n_7833),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7847),
.Y(n_7852)
);

AOI22xp5_ASAP7_75t_L g7853 ( 
.A1(n_7847),
.A2(n_7829),
.B1(n_7828),
.B2(n_7832),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_7843),
.Y(n_7854)
);

OAI22xp33_ASAP7_75t_L g7855 ( 
.A1(n_7849),
.A2(n_7831),
.B1(n_2112),
.B2(n_2104),
.Y(n_7855)
);

AOI22xp5_ASAP7_75t_L g7856 ( 
.A1(n_7848),
.A2(n_2104),
.B1(n_2103),
.B2(n_2097),
.Y(n_7856)
);

OR3x1_ASAP7_75t_L g7857 ( 
.A(n_7850),
.B(n_7844),
.C(n_7841),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_SL g7858 ( 
.A(n_7851),
.B(n_7840),
.Y(n_7858)
);

NOR3xp33_ASAP7_75t_L g7859 ( 
.A(n_7852),
.B(n_7846),
.C(n_7838),
.Y(n_7859)
);

AOI22xp5_ASAP7_75t_L g7860 ( 
.A1(n_7854),
.A2(n_7853),
.B1(n_7855),
.B2(n_7856),
.Y(n_7860)
);

AOI21xp5_ASAP7_75t_L g7861 ( 
.A1(n_7858),
.A2(n_7842),
.B(n_1721),
.Y(n_7861)
);

OAI22xp5_ASAP7_75t_L g7862 ( 
.A1(n_7860),
.A2(n_2104),
.B1(n_2103),
.B2(n_2097),
.Y(n_7862)
);

AND2x2_ASAP7_75t_L g7863 ( 
.A(n_7859),
.B(n_7857),
.Y(n_7863)
);

AOI22xp5_ASAP7_75t_L g7864 ( 
.A1(n_7863),
.A2(n_2103),
.B1(n_2097),
.B2(n_2093),
.Y(n_7864)
);

HB1xp67_ASAP7_75t_L g7865 ( 
.A(n_7862),
.Y(n_7865)
);

OAI21xp5_ASAP7_75t_L g7866 ( 
.A1(n_7865),
.A2(n_7861),
.B(n_1742),
.Y(n_7866)
);

OAI22xp5_ASAP7_75t_L g7867 ( 
.A1(n_7864),
.A2(n_2104),
.B1(n_2103),
.B2(n_2097),
.Y(n_7867)
);

AND2x2_ASAP7_75t_L g7868 ( 
.A(n_7866),
.B(n_2103),
.Y(n_7868)
);

OAI22xp33_ASAP7_75t_L g7869 ( 
.A1(n_7868),
.A2(n_7867),
.B1(n_2103),
.B2(n_2097),
.Y(n_7869)
);

AOI22xp5_ASAP7_75t_L g7870 ( 
.A1(n_7868),
.A2(n_2093),
.B1(n_2056),
.B2(n_1717),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7869),
.Y(n_7871)
);

NAND2xp5_ASAP7_75t_L g7872 ( 
.A(n_7870),
.B(n_2093),
.Y(n_7872)
);

OAI22xp33_ASAP7_75t_L g7873 ( 
.A1(n_7872),
.A2(n_2093),
.B1(n_2056),
.B2(n_1717),
.Y(n_7873)
);

AOI21xp5_ASAP7_75t_L g7874 ( 
.A1(n_7871),
.A2(n_1698),
.B(n_1707),
.Y(n_7874)
);

AOI221xp5_ASAP7_75t_L g7875 ( 
.A1(n_7873),
.A2(n_7874),
.B1(n_2056),
.B2(n_1717),
.C(n_1720),
.Y(n_7875)
);

AOI221xp5_ASAP7_75t_L g7876 ( 
.A1(n_7875),
.A2(n_2056),
.B1(n_1707),
.B2(n_1717),
.C(n_1720),
.Y(n_7876)
);

AOI211xp5_ASAP7_75t_L g7877 ( 
.A1(n_7876),
.A2(n_1698),
.B(n_1707),
.C(n_1717),
.Y(n_7877)
);


endmodule