module fake_netlist_6_547_n_890 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_890);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_890;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_683;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_796;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_811;
wire n_630;
wire n_394;
wire n_312;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_110),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_67),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_172),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_78),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_69),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_83),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_74),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_124),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_111),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_148),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_9),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_131),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_86),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_102),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_89),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_52),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_80),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_38),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_140),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_153),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_4),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_154),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_123),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_90),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_35),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_211),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_184),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_239),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_212),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_185),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_0),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_0),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_176),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_179),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_194),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_186),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_217),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_235),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_248),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_177),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_182),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_187),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_178),
.B(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_188),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_190),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_206),
.B(n_236),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_191),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_178),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_208),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_178),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_195),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_196),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

AND3x1_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_226),
.C(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_226),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_2),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_262),
.A2(n_198),
.B(n_197),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_199),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_289),
.B(n_257),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_289),
.B(n_200),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_201),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_275),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_254),
.B(n_246),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_265),
.B(n_204),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_263),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_245),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_209),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

NOR2x1p5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_210),
.Y(n_359)
);

BUFx6f_ASAP7_75t_SL g360 ( 
.A(n_344),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_326),
.Y(n_362)
);

OR2x6_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_214),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_281),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_337),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_215),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_219),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_283),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_319),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_220),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_222),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_225),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_283),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

NAND3x1_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_3),
.C(n_5),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_303),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_228),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_231),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_232),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_284),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_340),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_233),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_234),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_237),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_330),
.B(n_238),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_230),
.B1(n_221),
.B2(n_224),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_325),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_307),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_307),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_307),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_284),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_340),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_349),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_313),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_325),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_361),
.A2(n_317),
.B1(n_352),
.B2(n_351),
.Y(n_430)
);

OAI221xp5_ASAP7_75t_L g431 ( 
.A1(n_398),
.A2(n_424),
.B1(n_371),
.B2(n_425),
.C(n_414),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_352),
.B1(n_351),
.B2(n_355),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_388),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_328),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_332),
.B1(n_349),
.B2(n_346),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

NAND2x1p5_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_346),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_308),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_387),
.A2(n_309),
.B1(n_331),
.B2(n_349),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g447 ( 
.A1(n_383),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_409),
.A2(n_331),
.B1(n_349),
.B2(n_329),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_318),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_360),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_371),
.B(n_328),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

AO22x2_ASAP7_75t_L g455 ( 
.A1(n_383),
.A2(n_356),
.B1(n_323),
.B2(n_350),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_386),
.A2(n_331),
.B1(n_336),
.B2(n_339),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_360),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_358),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_378),
.A2(n_356),
.B1(n_380),
.B2(n_366),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_327),
.Y(n_471)
);

AO22x2_ASAP7_75t_L g472 ( 
.A1(n_378),
.A2(n_356),
.B1(n_323),
.B2(n_6),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_363),
.B(n_337),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

AO22x2_ASAP7_75t_L g477 ( 
.A1(n_380),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_477)
);

AO22x2_ASAP7_75t_L g478 ( 
.A1(n_366),
.A2(n_386),
.B1(n_391),
.B2(n_392),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_363),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_415),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_391),
.A2(n_404),
.B1(n_8),
.B2(n_9),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_404),
.B(n_327),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_367),
.B(n_241),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_376),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_488)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_377),
.A2(n_305),
.B(n_304),
.Y(n_489)
);

OAI221xp5_ASAP7_75t_L g490 ( 
.A1(n_363),
.A2(n_329),
.B1(n_327),
.B2(n_311),
.C(n_310),
.Y(n_490)
);

NAND2x1p5_ASAP7_75t_L g491 ( 
.A(n_419),
.B(n_304),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_401),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_359),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_384),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

OAI221xp5_ASAP7_75t_L g496 ( 
.A1(n_407),
.A2(n_310),
.B1(n_242),
.B2(n_335),
.C(n_307),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_335),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_285),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_442),
.B(n_426),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_443),
.B(n_426),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_457),
.B(n_467),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_429),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_476),
.B(n_417),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_452),
.B(n_357),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_370),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_433),
.B(n_370),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_437),
.B(n_417),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_453),
.B(n_417),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_436),
.B(n_369),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_484),
.B(n_369),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_462),
.B(n_373),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_459),
.B(n_369),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_441),
.B(n_369),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_479),
.B(n_373),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_471),
.B(n_393),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_428),
.B(n_418),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_427),
.B(n_393),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_482),
.B(n_483),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_434),
.B(n_420),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_435),
.B(n_420),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_438),
.B(n_421),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_440),
.B(n_396),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_389),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_444),
.B(n_397),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_486),
.B(n_406),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_446),
.B(n_399),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_465),
.B(n_411),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_451),
.B(n_416),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_448),
.B(n_374),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_491),
.B(n_374),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_466),
.B(n_379),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_489),
.B(n_379),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_469),
.B(n_379),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_312),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_474),
.B(n_312),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_487),
.B(n_475),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_480),
.B(n_312),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_481),
.B(n_221),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_449),
.B(n_221),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_464),
.B(n_221),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_430),
.B(n_312),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_454),
.B(n_224),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_456),
.B(n_224),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_375),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_468),
.B(n_12),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_458),
.B(n_460),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_461),
.B(n_224),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_463),
.B(n_494),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_12),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_478),
.B(n_431),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_505),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_430),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_516),
.A2(n_498),
.B(n_497),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_499),
.B(n_455),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_R g556 ( 
.A(n_515),
.B(n_495),
.Y(n_556)
);

AO31x2_ASAP7_75t_L g557 ( 
.A1(n_551),
.A2(n_447),
.A3(n_496),
.B(n_490),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_528),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_447),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_473),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_517),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_501),
.B(n_432),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_503),
.B(n_432),
.Y(n_563)
);

AOI21xp33_ASAP7_75t_L g564 ( 
.A1(n_545),
.A2(n_485),
.B(n_455),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_508),
.A2(n_375),
.B(n_485),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_513),
.A2(n_473),
.B(n_375),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_528),
.B(n_537),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_549),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_375),
.B(n_224),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_503),
.B(n_477),
.Y(n_571)
);

NOR4xp25_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_477),
.C(n_488),
.D(n_492),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_550),
.Y(n_574)
);

AOI211x1_ASAP7_75t_L g575 ( 
.A1(n_519),
.A2(n_492),
.B(n_472),
.C(n_15),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_538),
.A2(n_230),
.B(n_93),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_518),
.B(n_29),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

OAI21x1_ASAP7_75t_SL g579 ( 
.A1(n_534),
.A2(n_94),
.B(n_150),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_504),
.B(n_533),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_510),
.A2(n_472),
.B1(n_14),
.B2(n_16),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_520),
.A2(n_92),
.B(n_171),
.Y(n_583)
);

AO31x2_ASAP7_75t_L g584 ( 
.A1(n_527),
.A2(n_13),
.A3(n_14),
.B(n_16),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_500),
.B(n_33),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_509),
.A2(n_95),
.B(n_170),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_507),
.B(n_34),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_521),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_522),
.A2(n_97),
.B(n_169),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_529),
.Y(n_590)
);

AO31x2_ASAP7_75t_L g591 ( 
.A1(n_542),
.A2(n_13),
.A3(n_17),
.B(n_18),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_511),
.A2(n_88),
.B(n_167),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_532),
.A2(n_87),
.B(n_159),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_514),
.B(n_17),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_592),
.B(n_531),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_552),
.B(n_523),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_568),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_554),
.A2(n_576),
.B(n_559),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_570),
.A2(n_541),
.B(n_540),
.Y(n_600)
);

AOI221xp5_ASAP7_75t_L g601 ( 
.A1(n_582),
.A2(n_512),
.B1(n_539),
.B2(n_525),
.C(n_541),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_SL g602 ( 
.A1(n_585),
.A2(n_548),
.B(n_544),
.C(n_543),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_563),
.Y(n_603)
);

AO21x2_ASAP7_75t_L g604 ( 
.A1(n_565),
.A2(n_536),
.B(n_98),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_583),
.A2(n_82),
.B(n_157),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_589),
.A2(n_81),
.B(n_152),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_582),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_574),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_593),
.A2(n_100),
.B(n_149),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_567),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_36),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_580),
.A2(n_79),
.B(n_147),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_569),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_558),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_580),
.A2(n_77),
.B(n_146),
.Y(n_617)
);

OAI211xp5_ASAP7_75t_L g618 ( 
.A1(n_575),
.A2(n_20),
.B(n_23),
.C(n_24),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_588),
.Y(n_619)
);

NAND2x1p5_ASAP7_75t_L g620 ( 
.A(n_578),
.B(n_76),
.Y(n_620)
);

OAI221xp5_ASAP7_75t_L g621 ( 
.A1(n_590),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_566),
.A2(n_103),
.B(n_144),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_571),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_566),
.A2(n_101),
.B(n_143),
.Y(n_624)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_559),
.A2(n_25),
.B(n_26),
.Y(n_625)
);

AO31x2_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_27),
.A3(n_28),
.B(n_37),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_579),
.A2(n_105),
.B(n_39),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_585),
.A2(n_107),
.B(n_41),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_586),
.A2(n_108),
.B(n_44),
.Y(n_629)
);

OAI22x1_ASAP7_75t_L g630 ( 
.A1(n_555),
.A2(n_27),
.B1(n_45),
.B2(n_46),
.Y(n_630)
);

AO21x2_ASAP7_75t_L g631 ( 
.A1(n_564),
.A2(n_48),
.B(n_49),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_560),
.B(n_50),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_53),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_577),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_587),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_587),
.A2(n_59),
.B(n_60),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

CKINVDCx8_ASAP7_75t_R g638 ( 
.A(n_577),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_581),
.Y(n_639)
);

CKINVDCx6p67_ASAP7_75t_R g640 ( 
.A(n_616),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_619),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_619),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_612),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_609),
.B(n_572),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_611),
.B(n_572),
.Y(n_645)
);

NOR2x1_ASAP7_75t_L g646 ( 
.A(n_597),
.B(n_578),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_634),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_608),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_634),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_616),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_596),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_634),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_623),
.B(n_564),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_598),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_615),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_615),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_612),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_613),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_599),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_599),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_603),
.B(n_562),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_612),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_633),
.B(n_584),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_608),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_599),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_633),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_SL g670 ( 
.A1(n_614),
.A2(n_556),
.B(n_557),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_557),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_625),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

BUFx2_ASAP7_75t_SL g674 ( 
.A(n_638),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_630),
.Y(n_675)
);

AO21x1_ASAP7_75t_L g676 ( 
.A1(n_636),
.A2(n_584),
.B(n_591),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_625),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_620),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_625),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_638),
.B(n_607),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_600),
.A2(n_557),
.B(n_584),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_621),
.A2(n_591),
.B1(n_62),
.B2(n_63),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_620),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_630),
.B(n_591),
.Y(n_684)
);

CKINVDCx11_ASAP7_75t_R g685 ( 
.A(n_618),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_620),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_632),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_626),
.B(n_61),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_635),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_626),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_631),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_654),
.B(n_628),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_653),
.B(n_626),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_R g695 ( 
.A(n_647),
.B(n_70),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_674),
.B(n_610),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_648),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_R g698 ( 
.A(n_654),
.B(n_628),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_647),
.B(n_622),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_647),
.B(n_72),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_653),
.B(n_626),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_650),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_644),
.B(n_631),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_641),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_645),
.B(n_631),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_647),
.B(n_624),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_647),
.B(n_624),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_660),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_R g709 ( 
.A(n_649),
.B(n_652),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_687),
.B(n_617),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_642),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_649),
.B(n_627),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_649),
.B(n_652),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_649),
.B(n_627),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_649),
.B(n_610),
.Y(n_715)
);

XNOR2xp5_ASAP7_75t_L g716 ( 
.A(n_680),
.B(n_601),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_651),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_R g718 ( 
.A(n_659),
.B(n_606),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_R g719 ( 
.A(n_659),
.B(n_606),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_663),
.B(n_604),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_655),
.Y(n_721)
);

CKINVDCx12_ASAP7_75t_R g722 ( 
.A(n_663),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_646),
.B(n_604),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_R g724 ( 
.A(n_652),
.B(n_75),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_669),
.B(n_604),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_668),
.B(n_629),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_R g729 ( 
.A(n_659),
.B(n_605),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_650),
.Y(n_730)
);

OR2x4_ASAP7_75t_L g731 ( 
.A(n_652),
.B(n_602),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_656),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_640),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_668),
.B(n_629),
.Y(n_734)
);

XOR2x2_ASAP7_75t_SL g735 ( 
.A(n_689),
.B(n_595),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_657),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_736),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_717),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_699),
.B(n_672),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_711),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_694),
.B(n_692),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_701),
.B(n_690),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_716),
.A2(n_685),
.B1(n_675),
.B2(n_682),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_732),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_715),
.B(n_670),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_703),
.B(n_684),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_722),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_705),
.B(n_684),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_704),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_737),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_721),
.Y(n_752)
);

NOR2x1_ASAP7_75t_SL g753 ( 
.A(n_696),
.B(n_677),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_727),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_720),
.B(n_679),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_708),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_728),
.Y(n_757)
);

OAI221xp5_ASAP7_75t_SL g758 ( 
.A1(n_710),
.A2(n_688),
.B1(n_670),
.B2(n_691),
.C(n_665),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_697),
.B(n_671),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_731),
.A2(n_652),
.B1(n_640),
.B2(n_643),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_723),
.B(n_685),
.C(n_688),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_725),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_726),
.B(n_665),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_734),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_712),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_699),
.B(n_673),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_681),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_730),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_755),
.B(n_662),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_755),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_739),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_739),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_750),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_740),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_741),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_761),
.B(n_693),
.C(n_698),
.Y(n_777)
);

INVx5_ASAP7_75t_SL g778 ( 
.A(n_746),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_747),
.B(n_749),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_747),
.B(n_661),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_754),
.B(n_733),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_750),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_741),
.Y(n_783)
);

AO21x2_ASAP7_75t_L g784 ( 
.A1(n_753),
.A2(n_661),
.B(n_667),
.Y(n_784)
);

AO21x2_ASAP7_75t_L g785 ( 
.A1(n_753),
.A2(n_662),
.B(n_667),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_749),
.B(n_681),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_752),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_776),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_779),
.B(n_738),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_771),
.B(n_754),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_786),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_779),
.B(n_757),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_776),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_780),
.B(n_757),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_775),
.B(n_768),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_775),
.B(n_768),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_786),
.B(n_764),
.Y(n_797)
);

NOR2xp67_ASAP7_75t_L g798 ( 
.A(n_777),
.B(n_764),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_778),
.B(n_780),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_772),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_781),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_792),
.B(n_790),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_798),
.A2(n_746),
.B1(n_801),
.B2(n_789),
.Y(n_803)
);

AO221x2_ASAP7_75t_L g804 ( 
.A1(n_797),
.A2(n_760),
.B1(n_783),
.B2(n_759),
.C(n_765),
.Y(n_804)
);

AO221x2_ASAP7_75t_L g805 ( 
.A1(n_788),
.A2(n_765),
.B1(n_766),
.B2(n_773),
.C(n_756),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_789),
.B(n_738),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_791),
.B(n_795),
.Y(n_807)
);

AO221x2_ASAP7_75t_L g808 ( 
.A1(n_793),
.A2(n_766),
.B1(n_756),
.B2(n_772),
.C(n_782),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_794),
.B(n_770),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_799),
.B(n_748),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_R g811 ( 
.A(n_799),
.B(n_702),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_795),
.B(n_769),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_805),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_806),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_804),
.B(n_762),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_812),
.B(n_807),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_807),
.B(n_796),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_808),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_802),
.B(n_770),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_810),
.B(n_796),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_813),
.A2(n_803),
.B(n_758),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_816),
.B(n_702),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_814),
.B(n_809),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_818),
.A2(n_744),
.B(n_746),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_SL g825 ( 
.A1(n_815),
.A2(n_746),
.B(n_696),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_821),
.B(n_817),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_823),
.B(n_820),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_822),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_828),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_826),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_827),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_829),
.B(n_824),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_829),
.B(n_817),
.Y(n_834)
);

NOR4xp25_ASAP7_75t_L g835 ( 
.A(n_831),
.B(n_819),
.C(n_825),
.D(n_800),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_830),
.B(n_686),
.C(n_643),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_832),
.A2(n_811),
.B1(n_800),
.B2(n_751),
.C(n_745),
.Y(n_837)
);

AOI211xp5_ASAP7_75t_L g838 ( 
.A1(n_831),
.A2(n_700),
.B(n_724),
.C(n_695),
.Y(n_838)
);

NAND4xp25_ASAP7_75t_L g839 ( 
.A(n_831),
.B(n_713),
.C(n_686),
.D(n_763),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_835),
.A2(n_745),
.B1(n_751),
.B2(n_702),
.C(n_782),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_834),
.Y(n_841)
);

AOI221x1_ASAP7_75t_L g842 ( 
.A1(n_836),
.A2(n_713),
.B1(n_787),
.B2(n_774),
.C(n_658),
.Y(n_842)
);

OAI211xp5_ASAP7_75t_SL g843 ( 
.A1(n_833),
.A2(n_787),
.B(n_774),
.C(n_683),
.Y(n_843)
);

AO22x2_ASAP7_75t_SL g844 ( 
.A1(n_838),
.A2(n_709),
.B1(n_778),
.B2(n_763),
.Y(n_844)
);

OAI211xp5_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_837),
.B(n_686),
.C(n_643),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_833),
.A2(n_715),
.B(n_676),
.C(n_678),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_841),
.B(n_778),
.Y(n_847)
);

AOI31xp33_ASAP7_75t_L g848 ( 
.A1(n_840),
.A2(n_678),
.A3(n_714),
.B(n_676),
.Y(n_848)
);

NAND4xp75_ASAP7_75t_L g849 ( 
.A(n_842),
.B(n_844),
.C(n_845),
.D(n_846),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_843),
.A2(n_778),
.B1(n_740),
.B2(n_767),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_841),
.B(n_742),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_841),
.B(n_752),
.Y(n_852)
);

NOR2x1_ASAP7_75t_L g853 ( 
.A(n_841),
.B(n_785),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_849),
.B(n_740),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_R g855 ( 
.A(n_847),
.B(n_852),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_R g856 ( 
.A(n_851),
.B(n_104),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_SL g857 ( 
.A(n_848),
.B(n_718),
.C(n_719),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_850),
.B(n_112),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_R g859 ( 
.A(n_853),
.B(n_113),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_847),
.B(n_735),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_R g861 ( 
.A(n_847),
.B(n_114),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_847),
.B(n_714),
.Y(n_862)
);

OR5x1_ASAP7_75t_L g863 ( 
.A(n_854),
.B(n_785),
.C(n_784),
.D(n_122),
.E(n_125),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_860),
.A2(n_862),
.B(n_855),
.Y(n_864)
);

XOR2xp5_ASAP7_75t_L g865 ( 
.A(n_861),
.B(n_117),
.Y(n_865)
);

OAI311xp33_ASAP7_75t_L g866 ( 
.A1(n_858),
.A2(n_664),
.A3(n_673),
.B1(n_742),
.C1(n_743),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_856),
.B(n_743),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_859),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_857),
.Y(n_869)
);

XNOR2xp5_ASAP7_75t_L g870 ( 
.A(n_860),
.B(n_118),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_861),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_868),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_867),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_865),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_767),
.Y(n_875)
);

NOR2x1_ASAP7_75t_L g876 ( 
.A(n_871),
.B(n_785),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_872),
.A2(n_864),
.B(n_870),
.Y(n_877)
);

OAI211xp5_ASAP7_75t_L g878 ( 
.A1(n_873),
.A2(n_869),
.B(n_863),
.C(n_866),
.Y(n_878)
);

AOI31xp33_ASAP7_75t_SL g879 ( 
.A1(n_874),
.A2(n_126),
.A3(n_127),
.B(n_128),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_875),
.A2(n_767),
.B(n_707),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_877),
.A2(n_876),
.B1(n_707),
.B2(n_706),
.Y(n_881)
);

AOI31xp33_ASAP7_75t_L g882 ( 
.A1(n_878),
.A2(n_879),
.A3(n_880),
.B(n_729),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_882),
.Y(n_883)
);

XOR2xp5_ASAP7_75t_L g884 ( 
.A(n_881),
.B(n_130),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_883),
.A2(n_884),
.B1(n_784),
.B2(n_767),
.Y(n_885)
);

AOI21xp33_ASAP7_75t_SL g886 ( 
.A1(n_884),
.A2(n_132),
.B(n_133),
.Y(n_886)
);

XOR2xp5_ASAP7_75t_L g887 ( 
.A(n_885),
.B(n_134),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_886),
.Y(n_888)
);

OAI221xp5_ASAP7_75t_R g889 ( 
.A1(n_887),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_889)
);

AOI211xp5_ASAP7_75t_L g890 ( 
.A1(n_889),
.A2(n_888),
.B(n_139),
.C(n_141),
.Y(n_890)
);


endmodule