module fake_netlist_6_2922_n_1751 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1751);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1751;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_73),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_21),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_23),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_17),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_66),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_184),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_81),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_35),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_78),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_64),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_95),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_65),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_70),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_76),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_123),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_93),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_103),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_67),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_171),
.Y(n_239)
);

CKINVDCx11_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_136),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_106),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_58),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_28),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_37),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_30),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_114),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_79),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_46),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_14),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_82),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_131),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_122),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_154),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_28),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_145),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_182),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_118),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_80),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_92),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_41),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_129),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_49),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_111),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_48),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_126),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_61),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_94),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_74),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_110),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_117),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_20),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_29),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_52),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_88),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_54),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_24),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_77),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_97),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_86),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_180),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_19),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_1),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_22),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_32),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_89),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_155),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_61),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_37),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_175),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_75),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_7),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_57),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_9),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_83),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_90),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_159),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_91),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_139),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_33),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_185),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_38),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_51),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_32),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_153),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_156),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_59),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_160),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_25),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_172),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_10),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_144),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_72),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_26),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_113),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_98),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_62),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_165),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_31),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_178),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_45),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_16),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_31),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_161),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_39),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_24),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_55),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_104),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_140),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_143),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_58),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_205),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_274),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_274),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_246),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_1),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_2),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_301),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_240),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_250),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_346),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_232),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_235),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_236),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_265),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_238),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_309),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_200),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_331),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_208),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_237),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_244),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_241),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_242),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_258),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_248),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_281),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_298),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_279),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_259),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_261),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_262),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_267),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_280),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_200),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_188),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_268),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_359),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_188),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_283),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_286),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_332),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_328),
.B(n_3),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_269),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_270),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_314),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_197),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_288),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_200),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_272),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_294),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_275),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_277),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_190),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_289),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_292),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_196),
.B(n_4),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_200),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_302),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_212),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_291),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_295),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_296),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_231),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_297),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_196),
.B(n_4),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_300),
.B(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_234),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_187),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_187),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_212),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_193),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_212),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_206),
.B(n_6),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_291),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_305),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_382),
.B(n_276),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_421),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_384),
.B(n_206),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_211),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_364),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_386),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_389),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_363),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_364),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_401),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_402),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_404),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_409),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_410),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_211),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_264),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_199),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_366),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_368),
.B(n_304),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_366),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_416),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_367),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_375),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_369),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_369),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_383),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_371),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_390),
.B(n_293),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_371),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_433),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_423),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_435),
.B(n_436),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_430),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_440),
.B(n_293),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_293),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_377),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_378),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_449),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_432),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_418),
.B(n_271),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_441),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_455),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_395),
.B(n_306),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_391),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_439),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_379),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_378),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_450),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_380),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_381),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_264),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_387),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_381),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_407),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_323),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_370),
.B(n_452),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_417),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_397),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_440),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_398),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_392),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_451),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_457),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_529),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_527),
.A2(n_373),
.B1(n_453),
.B2(n_451),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_453),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_391),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_459),
.B(n_426),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_471),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_323),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_460),
.B(n_376),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_479),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_522),
.A2(n_446),
.B1(n_422),
.B2(n_447),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_526),
.A2(n_447),
.B1(n_454),
.B2(n_437),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_476),
.A2(n_418),
.B1(n_434),
.B2(n_429),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_501),
.B(n_376),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_530),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_230),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_530),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_512),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_532),
.A2(n_374),
.B1(n_316),
.B2(n_321),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_519),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_474),
.B(n_376),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_479),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_532),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_398),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_497),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_475),
.B(n_376),
.Y(n_570)
);

AND3x2_ASAP7_75t_L g571 ( 
.A(n_483),
.B(n_257),
.C(n_311),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_495),
.B(n_239),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_494),
.B(n_456),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_507),
.A2(n_278),
.B1(n_194),
.B2(n_198),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_500),
.B(n_399),
.Y(n_576)
);

NOR2x1p5_ASAP7_75t_L g577 ( 
.A(n_463),
.B(n_193),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_399),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_466),
.B(n_467),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_468),
.B(n_320),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_467),
.B(n_256),
.Y(n_582)
);

BUFx4f_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_477),
.B(n_273),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_469),
.B(n_306),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

AND3x4_ASAP7_75t_L g587 ( 
.A(n_458),
.B(n_374),
.C(n_243),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_464),
.B(n_400),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_471),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_478),
.B(n_326),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_470),
.B(n_400),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_472),
.B(n_403),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_471),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_480),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_480),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_473),
.B(n_291),
.Y(n_597)
);

INVxp33_ASAP7_75t_L g598 ( 
.A(n_483),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_485),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_485),
.A2(n_344),
.B1(n_350),
.B2(n_352),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_497),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_482),
.B(n_291),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_488),
.B(n_338),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_488),
.B(n_201),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_534),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_490),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_515),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_492),
.B(n_203),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_493),
.B(n_207),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_493),
.B(n_209),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_403),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_503),
.B(n_210),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_471),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_516),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_504),
.B(n_216),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_516),
.B(n_456),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_518),
.A2(n_330),
.B1(n_354),
.B2(n_356),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_518),
.B(n_217),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_520),
.A2(n_358),
.B1(n_443),
.B2(n_442),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_471),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_505),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_520),
.B(n_220),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_481),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_221),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_521),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_524),
.B(n_406),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_524),
.B(n_191),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_487),
.A2(n_347),
.B1(n_224),
.B2(n_227),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_229),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_509),
.B(n_233),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_481),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_514),
.B(n_445),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_481),
.B(n_249),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_465),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_481),
.B(n_255),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_481),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_481),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_508),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_508),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_508),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_508),
.B(n_263),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_505),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_517),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_508),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_458),
.B(n_408),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_486),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_511),
.A2(n_427),
.B1(n_443),
.B2(n_442),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_SL g656 ( 
.A(n_523),
.B(n_198),
.C(n_194),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_525),
.A2(n_202),
.B1(n_357),
.B2(n_353),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_528),
.B(n_408),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_511),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_511),
.B(n_282),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_511),
.B(n_287),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_511),
.Y(n_662)
);

BUFx8_ASAP7_75t_SL g663 ( 
.A(n_489),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_511),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_499),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_506),
.B(n_413),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_491),
.B(n_290),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_476),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_471),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_529),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_459),
.B(n_307),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_471),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_529),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_553),
.B(n_200),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_579),
.A2(n_355),
.B(n_361),
.C(n_336),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_579),
.A2(n_228),
.B1(n_360),
.B2(n_351),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_578),
.B(n_413),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_540),
.B(n_318),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_576),
.B(n_200),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_568),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_576),
.B(n_591),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_656),
.B(n_420),
.C(n_419),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_574),
.B(n_306),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_550),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_667),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_566),
.B(n_200),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_656),
.B(n_535),
.C(n_578),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_566),
.B(n_319),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_538),
.B(n_192),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_668),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_543),
.B(n_192),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_549),
.A2(n_226),
.B1(n_215),
.B2(n_213),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_549),
.A2(n_225),
.B1(n_215),
.B2(n_213),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_562),
.B(n_572),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_562),
.B(n_195),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_547),
.A2(n_202),
.B1(n_339),
.B2(n_218),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_543),
.B(n_195),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_591),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_668),
.B(n_204),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_574),
.B(n_204),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_609),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_592),
.B(n_219),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_588),
.B(n_223),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_588),
.B(n_223),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_539),
.B(n_419),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_539),
.B(n_556),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_585),
.A2(n_313),
.B1(n_218),
.B2(n_310),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_644),
.A2(n_392),
.B(n_438),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_545),
.B(n_225),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_SL g718 ( 
.A(n_587),
.B(n_310),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_570),
.B(n_669),
.Y(n_719)
);

AND2x6_ASAP7_75t_SL g720 ( 
.A(n_653),
.B(n_420),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

O2A1O1Ixp5_ASAP7_75t_L g722 ( 
.A1(n_672),
.A2(n_414),
.B(n_438),
.C(n_428),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_653),
.B(n_664),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_628),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_551),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_611),
.A2(n_623),
.B(n_602),
.C(n_597),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_564),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_542),
.B(n_324),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_663),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_640),
.B(n_324),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_SL g731 ( 
.A(n_589),
.B(n_327),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_669),
.B(n_327),
.Y(n_732)
);

AOI22x1_ASAP7_75t_L g733 ( 
.A1(n_635),
.A2(n_561),
.B1(n_555),
.B2(n_567),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_573),
.B(n_189),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_313),
.B1(n_312),
.B2(n_317),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_658),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_633),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_SL g739 ( 
.A(n_589),
.B(n_335),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_546),
.B(n_427),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_552),
.B(n_335),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_583),
.B(n_596),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_671),
.B(n_340),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_537),
.A2(n_340),
.B1(n_343),
.B2(n_342),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_583),
.B(n_343),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_445),
.C(n_431),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_674),
.B(n_349),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_675),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_597),
.B(n_245),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_565),
.B(n_428),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_602),
.B(n_247),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_596),
.B(n_251),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_569),
.B(n_252),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_589),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_632),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_586),
.B(n_253),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_594),
.B(n_266),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_626),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_637),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_555),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_607),
.Y(n_761)
);

CKINVDCx11_ASAP7_75t_R g762 ( 
.A(n_608),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_284),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_561),
.B(n_285),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_632),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_563),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_612),
.B(n_299),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_605),
.B(n_71),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_631),
.B(n_303),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_580),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_599),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_548),
.B(n_308),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_635),
.A2(n_334),
.B1(n_312),
.B2(n_317),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_618),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_615),
.Y(n_776)
);

XNOR2xp5_ASAP7_75t_L g777 ( 
.A(n_642),
.B(n_325),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_558),
.B(n_325),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_652),
.B(n_388),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_577),
.B(n_388),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_582),
.B(n_100),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_653),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_559),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_584),
.B(n_396),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_337),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_611),
.B(n_623),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_634),
.A2(n_339),
.B1(n_333),
.B2(n_357),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_603),
.B(n_189),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_598),
.B(n_189),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_598),
.B(n_341),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_541),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_SL g793 ( 
.A(n_589),
.B(n_353),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_627),
.B(n_348),
.Y(n_794)
);

INVx8_ASAP7_75t_L g795 ( 
.A(n_654),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_541),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_646),
.B(n_645),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_657),
.B(n_348),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_560),
.B(n_334),
.C(n_333),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_587),
.A2(n_396),
.B1(n_394),
.B2(n_341),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_627),
.B(n_394),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_646),
.B(n_147),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_647),
.B(n_141),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_657),
.B(n_341),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_604),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_627),
.B(n_132),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_608),
.B(n_329),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_613),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_648),
.B(n_659),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_651),
.B(n_329),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_571),
.B(n_181),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_666),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_655),
.B(n_329),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_571),
.B(n_243),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_662),
.B(n_130),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_665),
.B(n_128),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_595),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_614),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_650),
.B(n_243),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_655),
.B(n_173),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_700),
.B(n_616),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_687),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_755),
.B(n_600),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_762),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_678),
.A2(n_636),
.B(n_641),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_795),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_SL g827 ( 
.A(n_758),
.B(n_595),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_685),
.A2(n_627),
.B1(n_630),
.B2(n_619),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_704),
.B(n_650),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_792),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_678),
.A2(n_641),
.B(n_649),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_681),
.A2(n_575),
.B(n_638),
.C(n_649),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_734),
.B(n_560),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_771),
.B(n_627),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_761),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_772),
.A2(n_630),
.B1(n_638),
.B2(n_575),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_775),
.A2(n_600),
.B1(n_621),
.B2(n_624),
.Y(n_837)
);

BUFx4f_ASAP7_75t_L g838 ( 
.A(n_795),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_719),
.B(n_673),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_797),
.A2(n_624),
.B(n_621),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_719),
.B(n_673),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_754),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_676),
.A2(n_630),
.B(n_661),
.C(n_660),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_740),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_805),
.B(n_630),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_706),
.B(n_639),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_808),
.B(n_818),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_801),
.A2(n_670),
.B(n_617),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_776),
.B(n_630),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_720),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_710),
.B(n_711),
.Y(n_851)
);

OAI21xp33_ASAP7_75t_L g852 ( 
.A1(n_711),
.A2(n_639),
.B(n_629),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_809),
.A2(n_629),
.B(n_617),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_661),
.B(n_660),
.Y(n_854)
);

AO22x1_ASAP7_75t_L g855 ( 
.A1(n_798),
.A2(n_741),
.B1(n_693),
.B2(n_811),
.Y(n_855)
);

CKINVDCx10_ASAP7_75t_R g856 ( 
.A(n_723),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_778),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_765),
.B(n_712),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_754),
.A2(n_629),
.B(n_622),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_736),
.B(n_625),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_787),
.A2(n_661),
.B1(n_660),
.B2(n_643),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_726),
.A2(n_751),
.B(n_749),
.C(n_786),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_787),
.A2(n_661),
.B1(n_660),
.B2(n_643),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_712),
.B(n_593),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_691),
.Y(n_865)
);

BUFx4f_ASAP7_75t_L g866 ( 
.A(n_795),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_692),
.A2(n_625),
.B(n_622),
.Y(n_867)
);

OA22x2_ASAP7_75t_L g868 ( 
.A1(n_800),
.A2(n_12),
.B1(n_13),
.B2(n_19),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_716),
.A2(n_661),
.B1(n_660),
.B2(n_643),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_690),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_786),
.B(n_593),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_701),
.B(n_643),
.Y(n_872)
);

NAND2x2_ASAP7_75t_L g873 ( 
.A(n_721),
.B(n_13),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_688),
.B(n_125),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_759),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_708),
.B(n_717),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_810),
.B(n_25),
.Y(n_877)
);

BUFx4f_ASAP7_75t_L g878 ( 
.A(n_817),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_738),
.B(n_149),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_682),
.A2(n_643),
.B(n_166),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_767),
.B(n_163),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_682),
.A2(n_162),
.B(n_151),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_780),
.A2(n_742),
.B(n_806),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_749),
.B(n_150),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_742),
.A2(n_121),
.B(n_116),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_715),
.A2(n_102),
.B(n_101),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_766),
.Y(n_887)
);

NOR2xp67_ASAP7_75t_SL g888 ( 
.A(n_754),
.B(n_34),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_754),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_727),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_697),
.B(n_34),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_713),
.A2(n_85),
.B(n_84),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_697),
.B(n_819),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_728),
.A2(n_44),
.B(n_47),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_764),
.A2(n_50),
.B(n_52),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_696),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

OAI22x1_ASAP7_75t_L g898 ( 
.A1(n_798),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_785),
.B(n_56),
.Y(n_899)
);

AO32x1_ASAP7_75t_L g900 ( 
.A1(n_698),
.A2(n_59),
.A3(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_741),
.B(n_60),
.C(n_63),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_722),
.A2(n_733),
.B(n_705),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_753),
.B(n_756),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_696),
.A2(n_792),
.B(n_796),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_753),
.B(n_756),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_723),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_709),
.B(n_812),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_732),
.B(n_730),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_783),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_784),
.Y(n_910)
);

INVx6_ASAP7_75t_L g911 ( 
.A(n_783),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_702),
.B(n_735),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_781),
.B(n_811),
.Y(n_913)
);

NOR2x1_ASAP7_75t_L g914 ( 
.A(n_807),
.B(n_769),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_802),
.A2(n_803),
.B(n_816),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_702),
.A2(n_679),
.B(n_788),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_820),
.A2(n_694),
.B(n_773),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_729),
.B(n_783),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_768),
.B(n_757),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_683),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_750),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_763),
.B(n_770),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_744),
.A2(n_695),
.B1(n_680),
.B2(n_747),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_752),
.A2(n_745),
.B1(n_773),
.B2(n_695),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_684),
.A2(n_707),
.B(n_724),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_689),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_737),
.A2(n_743),
.B(n_779),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_779),
.A2(n_815),
.B(n_752),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_750),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_782),
.A2(n_794),
.B1(n_750),
.B2(n_703),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_813),
.A2(n_677),
.B(n_789),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_813),
.A2(n_791),
.B(n_790),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_699),
.B(n_750),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_777),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_746),
.A2(n_804),
.B(n_686),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_723),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_750),
.A2(n_774),
.B1(n_718),
.B2(n_799),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_814),
.A2(n_714),
.B(n_731),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_793),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_814),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_739),
.B(n_714),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_700),
.B(n_771),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_704),
.B(n_700),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_704),
.B(n_700),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_700),
.A2(n_685),
.B1(n_775),
.B2(n_772),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_761),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_700),
.A2(n_676),
.B(n_722),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_700),
.B(n_704),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_700),
.B(n_771),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_710),
.A2(n_711),
.B(n_741),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_704),
.B(n_700),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_700),
.A2(n_676),
.B(n_722),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_700),
.B(n_704),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_700),
.B(n_771),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

NOR2x1_ASAP7_75t_L g957 ( 
.A(n_685),
.B(n_574),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_685),
.A2(n_681),
.B(n_543),
.C(n_700),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_704),
.B(n_578),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_761),
.Y(n_960)
);

AO21x1_ASAP7_75t_L g961 ( 
.A1(n_700),
.A2(n_681),
.B(n_726),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_700),
.B(n_771),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_710),
.A2(n_711),
.B(n_700),
.C(n_726),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_755),
.B(n_765),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_700),
.B(n_771),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_678),
.A2(n_760),
.B(n_725),
.Y(n_966)
);

BUFx8_ASAP7_75t_SL g967 ( 
.A(n_729),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_758),
.B(n_574),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_700),
.B(n_771),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_678),
.A2(n_760),
.B(n_725),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_691),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_700),
.B(n_771),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_754),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_700),
.B(n_704),
.Y(n_974)
);

AND3x2_ASAP7_75t_L g975 ( 
.A(n_851),
.B(n_827),
.C(n_887),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_959),
.B(n_944),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_850),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_961),
.A2(n_862),
.A3(n_963),
.B(n_883),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_844),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_951),
.A2(n_953),
.B(n_948),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_912),
.B(n_838),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_822),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_943),
.A2(n_965),
.B1(n_955),
.B2(n_972),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_826),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_973),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_950),
.B(n_962),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_SL g987 ( 
.A1(n_896),
.A2(n_970),
.B(n_966),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_867),
.A2(n_904),
.B(n_902),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_973),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_969),
.B(n_945),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_952),
.B(n_821),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_893),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_870),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_946),
.B(n_919),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_968),
.B(n_957),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_897),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_890),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_896),
.B(n_842),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_837),
.A2(n_916),
.B1(n_938),
.B2(n_836),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_949),
.B(n_954),
.Y(n_1000)
);

NAND2x1_ASAP7_75t_L g1001 ( 
.A(n_842),
.B(n_830),
.Y(n_1001)
);

INVx5_ASAP7_75t_L g1002 ( 
.A(n_973),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_917),
.A2(n_934),
.B(n_883),
.Y(n_1003)
);

INVx8_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_974),
.B(n_829),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_907),
.B(n_923),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_911),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_865),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_922),
.B(n_958),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_847),
.B(n_833),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_855),
.B(n_908),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_924),
.B(n_936),
.C(n_901),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_830),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_917),
.A2(n_843),
.B(n_840),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_913),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_832),
.A2(n_929),
.B(n_849),
.Y(n_1016)
);

NAND2x1_ASAP7_75t_L g1017 ( 
.A(n_921),
.B(n_911),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_936),
.B(n_941),
.Y(n_1018)
);

AND3x4_ASAP7_75t_L g1019 ( 
.A(n_914),
.B(n_858),
.C(n_964),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_909),
.B(n_858),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_825),
.A2(n_853),
.B(n_848),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_823),
.B(n_927),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_971),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_911),
.Y(n_1024)
);

AND3x4_ASAP7_75t_L g1025 ( 
.A(n_964),
.B(n_823),
.C(n_856),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_891),
.A2(n_942),
.B1(n_931),
.B2(n_876),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_910),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_939),
.A2(n_932),
.B(n_933),
.C(n_929),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_831),
.A2(n_859),
.B(n_927),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_932),
.A2(n_834),
.B(n_831),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_967),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_877),
.B(n_941),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_915),
.A2(n_854),
.B(n_925),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_835),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_909),
.B(n_928),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_872),
.A2(n_845),
.B(n_930),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_880),
.A2(n_885),
.B(n_882),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_871),
.A2(n_852),
.B(n_841),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_899),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_838),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_839),
.B(n_960),
.Y(n_1041)
);

OAI22x1_ASAP7_75t_L g1042 ( 
.A1(n_906),
.A2(n_937),
.B1(n_935),
.B2(n_940),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_828),
.A2(n_884),
.B(n_880),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_889),
.A2(n_846),
.B(n_864),
.Y(n_1044)
);

CKINVDCx16_ASAP7_75t_R g1045 ( 
.A(n_918),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_881),
.A2(n_879),
.B(n_874),
.C(n_885),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_933),
.B(n_956),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_866),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_947),
.B(n_860),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_861),
.A2(n_863),
.B(n_895),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_882),
.A2(n_886),
.B(n_892),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_920),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_875),
.A2(n_926),
.B(n_869),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_888),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_824),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_894),
.B(n_868),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_866),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_868),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_857),
.A2(n_900),
.B(n_873),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_900),
.A2(n_851),
.B1(n_912),
.B2(n_943),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_900),
.A2(n_898),
.B(n_878),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_851),
.A2(n_912),
.B1(n_950),
.B2(n_943),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_851),
.B(n_943),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_822),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_L g1065 ( 
.A(n_968),
.B(n_574),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_959),
.B(n_944),
.Y(n_1066)
);

INVx3_ASAP7_75t_SL g1067 ( 
.A(n_826),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_959),
.B(n_944),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_844),
.Y(n_1069)
);

NAND2x1_ASAP7_75t_L g1070 ( 
.A(n_896),
.B(n_678),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_887),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_961),
.A2(n_862),
.A3(n_963),
.B(n_851),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_851),
.A2(n_951),
.B(n_905),
.C(n_903),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_951),
.B(n_851),
.C(n_903),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_961),
.A2(n_862),
.A3(n_963),
.B(n_851),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_851),
.A2(n_951),
.B(n_903),
.C(n_905),
.Y(n_1076)
);

INVx3_ASAP7_75t_SL g1077 ( 
.A(n_826),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_973),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_967),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_L g1080 ( 
.A(n_862),
.B(n_903),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_973),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_SL g1082 ( 
.A(n_896),
.B(n_973),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_890),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_896),
.B(n_842),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_851),
.B(n_943),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_851),
.B(n_944),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_851),
.B(n_944),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_890),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_973),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_851),
.A2(n_951),
.B(n_905),
.C(n_903),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_851),
.B(n_951),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_959),
.B(n_944),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_902),
.A2(n_953),
.B(n_948),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_967),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_851),
.B(n_943),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_851),
.A2(n_963),
.B(n_951),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_851),
.B(n_943),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1080),
.A2(n_1038),
.B(n_1009),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1071),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1086),
.A2(n_1087),
.B1(n_1085),
.B2(n_1095),
.Y(n_1100)
);

INVx3_ASAP7_75t_SL g1101 ( 
.A(n_1067),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_976),
.B(n_1066),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1068),
.B(n_1092),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_1004),
.B(n_1040),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_1091),
.A2(n_1096),
.B(n_1011),
.C(n_1016),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_1024),
.B(n_1002),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_993),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_979),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1055),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_985),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_994),
.A2(n_1043),
.B(n_1030),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_991),
.A2(n_990),
.B(n_1063),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1063),
.B(n_1085),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_992),
.B(n_1032),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_979),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_996),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1020),
.B(n_1035),
.Y(n_1117)
);

AO32x1_ASAP7_75t_L g1118 ( 
.A1(n_1060),
.A2(n_999),
.A3(n_1026),
.B1(n_1062),
.B2(n_983),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_SL g1119 ( 
.A1(n_1006),
.A2(n_1096),
.B(n_1060),
.C(n_1018),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1020),
.B(n_1035),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1024),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_1004),
.B(n_1040),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1024),
.B(n_1002),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_1039),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_1012),
.B(n_986),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1064),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1069),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_994),
.A2(n_1043),
.B(n_1030),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_L g1130 ( 
.A(n_1065),
.B(n_1048),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1069),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1024),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_990),
.B(n_983),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1023),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1008),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1017),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1003),
.A2(n_1028),
.B(n_987),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1015),
.B(n_1007),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_1002),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1039),
.B(n_1005),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1073),
.A2(n_1090),
.B1(n_1074),
.B2(n_1062),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_1002),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1007),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1014),
.A2(n_1003),
.B(n_980),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1000),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1083),
.Y(n_1148)
);

BUFx12f_ASAP7_75t_L g1149 ( 
.A(n_1057),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1007),
.B(n_1088),
.Y(n_1150)
);

BUFx4_ASAP7_75t_SL g1151 ( 
.A(n_1031),
.Y(n_1151)
);

BUFx4_ASAP7_75t_SL g1152 ( 
.A(n_1079),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1034),
.B(n_1027),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1010),
.B(n_1000),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1045),
.B(n_981),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_998),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1061),
.A2(n_980),
.B(n_1047),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_1049),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1052),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1004),
.B(n_984),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1058),
.B(n_1034),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1025),
.A2(n_1019),
.B1(n_1022),
.B2(n_1056),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_975),
.B(n_1082),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_985),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_1014),
.A2(n_1033),
.B(n_988),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

OAI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1041),
.A2(n_1054),
.B(n_1042),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1041),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_995),
.B(n_1013),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1050),
.B(n_1053),
.C(n_1046),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_985),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1050),
.A2(n_1037),
.B(n_1044),
.C(n_1051),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_978),
.B(n_989),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1093),
.A2(n_1084),
.B1(n_1078),
.B2(n_1081),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1077),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1078),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1093),
.B(n_1089),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1078),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1081),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1081),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1089),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1094),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1089),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1001),
.Y(n_1187)
);

NAND2x1_ASAP7_75t_L g1188 ( 
.A(n_1084),
.B(n_1070),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1036),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1059),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1029),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1021),
.B(n_977),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1091),
.A2(n_951),
.B1(n_851),
.B2(n_912),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1091),
.A2(n_851),
.B(n_951),
.C(n_1076),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1024),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_979),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1024),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_976),
.B(n_1066),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_982),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1071),
.Y(n_1200)
);

BUFx8_ASAP7_75t_L g1201 ( 
.A(n_977),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1020),
.B(n_1035),
.Y(n_1202)
);

OR2x2_ASAP7_75t_SL g1203 ( 
.A(n_1045),
.B(n_458),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1091),
.B(n_951),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1091),
.A2(n_951),
.B1(n_851),
.B2(n_912),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1091),
.A2(n_951),
.B(n_851),
.C(n_1073),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1071),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1004),
.B(n_795),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_976),
.B(n_1066),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1063),
.B(n_1085),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_979),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_976),
.B(n_1066),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1063),
.B(n_1085),
.Y(n_1213)
);

BUFx2_ASAP7_75t_SL g1214 ( 
.A(n_1024),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1024),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_1012),
.B(n_946),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1024),
.B(n_1002),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_851),
.B1(n_1087),
.B2(n_1085),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1219)
);

OAI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1091),
.A2(n_851),
.B(n_1086),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1024),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1020),
.B(n_1035),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1004),
.B(n_795),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_979),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1024),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1020),
.B(n_1035),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1055),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1071),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1169),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1218),
.A2(n_1100),
.B1(n_1158),
.B2(n_1141),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1170),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1172),
.Y(n_1234)
);

INVx6_ASAP7_75t_L g1235 ( 
.A(n_1215),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1218),
.B(n_1219),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1108),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1141),
.A2(n_1206),
.B(n_1098),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1132),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_SL g1240 ( 
.A(n_1149),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1215),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1100),
.A2(n_1140),
.B1(n_1225),
.B2(n_1223),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1180),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1193),
.A2(n_1205),
.B1(n_1204),
.B2(n_1220),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1132),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1115),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1220),
.A2(n_1126),
.B1(n_1216),
.B2(n_1162),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1199),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1105),
.B(n_1133),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1126),
.A2(n_1216),
.B1(n_1162),
.B2(n_1167),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1180),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1131),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1123),
.A2(n_1210),
.B1(n_1113),
.B2(n_1213),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1196),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1137),
.B(n_1192),
.Y(n_1256)
);

CKINVDCx8_ASAP7_75t_R g1257 ( 
.A(n_1214),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1147),
.B(n_1142),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1190),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1190),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1167),
.A2(n_1212),
.B1(n_1209),
.B2(n_1102),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1154),
.B(n_1168),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1229),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1155),
.A2(n_1198),
.B1(n_1103),
.B2(n_1112),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1157),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1112),
.A2(n_1178),
.B1(n_1114),
.B2(n_1163),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1173),
.A2(n_1163),
.B1(n_1125),
.B2(n_1178),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1107),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1151),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1116),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1175),
.A2(n_1129),
.B(n_1111),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1152),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1131),
.Y(n_1273)
);

INVx3_ASAP7_75t_SL g1274 ( 
.A(n_1195),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1127),
.Y(n_1275)
);

AO21x1_ASAP7_75t_SL g1276 ( 
.A1(n_1187),
.A2(n_1118),
.B(n_1119),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1121),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1211),
.A2(n_1226),
.B1(n_1135),
.B2(n_1128),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1211),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1161),
.B1(n_1101),
.B2(n_1153),
.Y(n_1280)
);

AND2x4_ASAP7_75t_SL g1281 ( 
.A(n_1227),
.B(n_1122),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1146),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1106),
.Y(n_1283)
);

OAI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1208),
.A2(n_1224),
.B1(n_1160),
.B2(n_1122),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1134),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1189),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1159),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1188),
.B(n_1165),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1124),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1117),
.B(n_1202),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1177),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1160),
.A2(n_1153),
.B1(n_1148),
.B2(n_1144),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1191),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

BUFx8_ASAP7_75t_SL g1295 ( 
.A(n_1109),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1145),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1164),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1118),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1136),
.Y(n_1299)
);

BUFx8_ASAP7_75t_SL g1300 ( 
.A(n_1207),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1118),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1201),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1117),
.B(n_1222),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1156),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1171),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1208),
.A2(n_1224),
.B1(n_1104),
.B2(n_1122),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1156),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1179),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1197),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1181),
.A2(n_1186),
.B(n_1184),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1201),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1182),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1166),
.A2(n_1228),
.B1(n_1202),
.B2(n_1222),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1138),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1183),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1150),
.A2(n_1228),
.B(n_1120),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1221),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1203),
.A2(n_1120),
.B1(n_1104),
.B2(n_1224),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1138),
.A2(n_1230),
.B1(n_1150),
.B2(n_1104),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1110),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1145),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1110),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1185),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1110),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1217),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1208),
.A2(n_1099),
.B1(n_1200),
.B2(n_1130),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1145),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1139),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1143),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1143),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1174),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1174),
.Y(n_1332)
);

BUFx2_ASAP7_75t_R g1333 ( 
.A(n_1207),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1132),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1218),
.A2(n_851),
.B1(n_912),
.B2(n_1091),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1108),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1147),
.B(n_1193),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1176),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1115),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1229),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1108),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1147),
.B(n_1193),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1132),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1108),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1194),
.A2(n_851),
.B(n_951),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1176),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1282),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1297),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1283),
.Y(n_1350)
);

INVx4_ASAP7_75t_SL g1351 ( 
.A(n_1256),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1259),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1288),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1256),
.B(n_1238),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1256),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1273),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1256),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1246),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1288),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1297),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1293),
.B(n_1286),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1310),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1259),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1295),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1258),
.B(n_1338),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1255),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1346),
.B(n_1250),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1288),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1335),
.A2(n_1244),
.B1(n_1345),
.B2(n_1232),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1231),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1260),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1337),
.B(n_1342),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1254),
.A2(n_1236),
.B(n_1284),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1242),
.A2(n_1247),
.B(n_1251),
.Y(n_1376)
);

NAND2x1_ASAP7_75t_L g1377 ( 
.A(n_1286),
.B(n_1293),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1233),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1233),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1340),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1234),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1234),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1260),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1268),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1316),
.B(n_1299),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1291),
.B(n_1294),
.Y(n_1387)
);

OAI21xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1262),
.A2(n_1266),
.B(n_1270),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1291),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1287),
.B(n_1298),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1339),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1253),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1287),
.B(n_1298),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1237),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1257),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1310),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1301),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1279),
.B(n_1264),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1261),
.A2(n_1318),
.B(n_1292),
.C(n_1305),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1301),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1294),
.A2(n_1305),
.B(n_1275),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_SL g1403 ( 
.A(n_1333),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1344),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1271),
.B(n_1344),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1249),
.Y(n_1406)
);

NOR2x1_ASAP7_75t_L g1407 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1267),
.A2(n_1285),
.B(n_1280),
.Y(n_1408)
);

AOI21xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1323),
.A2(n_1278),
.B(n_1326),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1328),
.A2(n_1330),
.B(n_1317),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1290),
.B(n_1303),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1317),
.A2(n_1330),
.B(n_1328),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1283),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1336),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1283),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1348),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1390),
.B(n_1276),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1405),
.B(n_1341),
.Y(n_1419)
);

AOI33xp33_ASAP7_75t_L g1420 ( 
.A1(n_1370),
.A2(n_1312),
.A3(n_1319),
.B1(n_1315),
.B2(n_1313),
.B3(n_1327),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.B(n_1308),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1351),
.B(n_1304),
.Y(n_1422)
);

NAND2xp33_ASAP7_75t_R g1423 ( 
.A(n_1380),
.B(n_1272),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1393),
.B(n_1308),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1329),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1405),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1351),
.B(n_1355),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1314),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1385),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1360),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1355),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1374),
.B(n_1356),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1381),
.B(n_1316),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1376),
.A2(n_1303),
.B1(n_1311),
.B2(n_1240),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1381),
.B(n_1368),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1408),
.A2(n_1309),
.B1(n_1248),
.B2(n_1277),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1358),
.B(n_1309),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1349),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1415),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1375),
.B(n_1412),
.Y(n_1440)
);

NOR2x1p5_ASAP7_75t_L g1441 ( 
.A(n_1355),
.B(n_1241),
.Y(n_1441)
);

NAND2x1_ASAP7_75t_L g1442 ( 
.A(n_1354),
.B(n_1235),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1388),
.A2(n_1325),
.B1(n_1331),
.B2(n_1321),
.C(n_1323),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1387),
.B(n_1332),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1392),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1397),
.Y(n_1446)
);

AND2x2_ASAP7_75t_SL g1447 ( 
.A(n_1402),
.B(n_1281),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1387),
.B(n_1398),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1401),
.B(n_1296),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1366),
.B(n_1325),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1384),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1389),
.B(n_1402),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1407),
.A2(n_1289),
.B1(n_1283),
.B2(n_1235),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1391),
.B(n_1245),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1365),
.B(n_1245),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1389),
.B(n_1296),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1386),
.B(n_1239),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1434),
.A2(n_1409),
.B(n_1400),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1433),
.B(n_1402),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1394),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1409),
.C(n_1407),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1443),
.C(n_1436),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1445),
.B(n_1414),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1420),
.B(n_1388),
.C(n_1399),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1425),
.B(n_1447),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_L g1466 ( 
.A(n_1425),
.B(n_1413),
.C(n_1350),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1433),
.B(n_1402),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1435),
.B(n_1354),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1428),
.B(n_1404),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1457),
.B(n_1354),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1437),
.B(n_1394),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1453),
.A2(n_1395),
.B1(n_1403),
.B2(n_1354),
.Y(n_1472)
);

NOR3xp33_ASAP7_75t_L g1473 ( 
.A(n_1450),
.B(n_1350),
.C(n_1413),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1447),
.A2(n_1386),
.B(n_1411),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1441),
.B(n_1355),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1447),
.B(n_1355),
.Y(n_1476)
);

OAI21xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1441),
.A2(n_1349),
.B(n_1383),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1442),
.B(n_1355),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1419),
.A2(n_1357),
.B1(n_1442),
.B2(n_1454),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1427),
.A2(n_1357),
.B(n_1281),
.Y(n_1480)
);

NOR3xp33_ASAP7_75t_L g1481 ( 
.A(n_1418),
.B(n_1350),
.C(n_1413),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1417),
.B(n_1362),
.Y(n_1482)
);

OAI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1426),
.A2(n_1367),
.B1(n_1357),
.B2(n_1350),
.C(n_1413),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1449),
.B(n_1377),
.C(n_1383),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1449),
.B(n_1377),
.C(n_1372),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1444),
.B(n_1347),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1438),
.B(n_1382),
.C(n_1379),
.Y(n_1487)
);

NAND4xp25_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1352),
.C(n_1363),
.D(n_1373),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1452),
.A2(n_1357),
.B(n_1406),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1372),
.C(n_1371),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1451),
.A2(n_1361),
.B1(n_1382),
.B2(n_1371),
.C(n_1379),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1427),
.A2(n_1324),
.B(n_1320),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1421),
.B(n_1396),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1427),
.A2(n_1415),
.B1(n_1369),
.B2(n_1359),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1451),
.A2(n_1361),
.B1(n_1378),
.B2(n_1373),
.C(n_1352),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_L g1496 ( 
.A(n_1418),
.B(n_1343),
.C(n_1410),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1455),
.B(n_1364),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1421),
.B(n_1396),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1424),
.B(n_1353),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1429),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1422),
.B(n_1351),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1500),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1459),
.B(n_1446),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1467),
.B(n_1448),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1468),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1493),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1478),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1498),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1470),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1501),
.B(n_1427),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1470),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1490),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1501),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1484),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1477),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1489),
.B(n_1416),
.Y(n_1520)
);

NOR2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1461),
.B(n_1439),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1488),
.B(n_1448),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1475),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1471),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1496),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1502),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1460),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1511),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1504),
.B(n_1465),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1513),
.B(n_1491),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1518),
.B(n_1476),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1511),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1511),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1525),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1508),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1507),
.B(n_1509),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1517),
.B(n_1430),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1518),
.B(n_1473),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1514),
.B(n_1458),
.C(n_1464),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1508),
.Y(n_1545)
);

INVx3_ASAP7_75t_SL g1546 ( 
.A(n_1516),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1507),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1512),
.B(n_1494),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1520),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1508),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1502),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1481),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1469),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1431),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1506),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1506),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1517),
.B(n_1495),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1520),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1525),
.B(n_1429),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1507),
.B(n_1466),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1506),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1554),
.B(n_1527),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1562),
.B(n_1509),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_SL g1569 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1554),
.B(n_1527),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1564),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1544),
.A2(n_1462),
.B1(n_1524),
.B2(n_1523),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1559),
.A2(n_1521),
.B1(n_1523),
.B2(n_1524),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1521),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1563),
.B(n_1526),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1528),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1562),
.B(n_1523),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1539),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1562),
.B(n_1524),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1538),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1531),
.A2(n_1474),
.B(n_1522),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1529),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1564),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1526),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1531),
.B(n_1503),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1552),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1534),
.B(n_1550),
.Y(n_1590)
);

INVxp33_ASAP7_75t_L g1591 ( 
.A(n_1543),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1534),
.B(n_1522),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.B(n_1503),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1535),
.A2(n_1521),
.B(n_1516),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1547),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1558),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1564),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1543),
.B(n_1522),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_SL g1601 ( 
.A(n_1547),
.B(n_1483),
.C(n_1492),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1535),
.B(n_1510),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1548),
.B(n_1516),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1548),
.B(n_1510),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1558),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1541),
.B(n_1505),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1541),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1540),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1566),
.B(n_1561),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1546),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1578),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1567),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1567),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1569),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1579),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1579),
.B(n_1546),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1571),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1570),
.B(n_1533),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1576),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1568),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1533),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1580),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1607),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1580),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1608),
.B(n_1532),
.Y(n_1632)
);

AND3x1_ASAP7_75t_L g1633 ( 
.A(n_1573),
.B(n_1553),
.C(n_1555),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1588),
.B(n_1582),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1572),
.A2(n_1511),
.B1(n_1536),
.B2(n_1532),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1584),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1571),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1588),
.B(n_1530),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1569),
.B(n_1555),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1585),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1604),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1584),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1587),
.B(n_1530),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1586),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1574),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1592),
.B(n_1515),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1574),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1619),
.B(n_1591),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1637),
.Y(n_1650)
);

O2A1O1Ixp33_ASAP7_75t_SL g1651 ( 
.A1(n_1618),
.A2(n_1601),
.B(n_1610),
.C(n_1302),
.Y(n_1651)
);

OAI32xp33_ASAP7_75t_L g1652 ( 
.A1(n_1642),
.A2(n_1594),
.A3(n_1600),
.B1(n_1583),
.B2(n_1575),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1633),
.A2(n_1578),
.B1(n_1574),
.B2(n_1608),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1640),
.A2(n_1578),
.B1(n_1537),
.B2(n_1536),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1633),
.A2(n_1605),
.B1(n_1607),
.B2(n_1602),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1619),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1613),
.A2(n_1605),
.B1(n_1602),
.B2(n_1581),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1614),
.B(n_1581),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1616),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1617),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1625),
.A2(n_1609),
.B(n_1603),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1617),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1635),
.A2(n_1648),
.B(n_1646),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1615),
.B(n_1269),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1624),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1629),
.B(n_1593),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1615),
.B(n_1272),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1629),
.B(n_1593),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

OAI32xp33_ASAP7_75t_L g1675 ( 
.A1(n_1634),
.A2(n_1586),
.A3(n_1589),
.B1(n_1537),
.B2(n_1595),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1626),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1613),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1653),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1655),
.B(n_1615),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1652),
.A2(n_1615),
.B1(n_1613),
.B2(n_1612),
.C(n_1630),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1654),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1653),
.Y(n_1683)
);

NOR2xp67_ASAP7_75t_SL g1684 ( 
.A(n_1663),
.B(n_1627),
.Y(n_1684)
);

INVx8_ASAP7_75t_L g1685 ( 
.A(n_1672),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1649),
.B(n_1671),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1651),
.A2(n_1630),
.B1(n_1623),
.B2(n_1472),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1674),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1665),
.B(n_1634),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1674),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1667),
.B(n_1659),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1654),
.Y(n_1693)
);

OAI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1657),
.A2(n_1660),
.B1(n_1662),
.B2(n_1661),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1660),
.B(n_1644),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1621),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1666),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1652),
.B1(n_1651),
.B2(n_1675),
.C(n_1656),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1692),
.A2(n_1675),
.B(n_1664),
.C(n_1668),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1682),
.B(n_1676),
.C(n_1670),
.D(n_1621),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1687),
.B(n_1679),
.C(n_1678),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1694),
.A2(n_1670),
.B(n_1647),
.Y(n_1703)
);

OAI322xp33_ASAP7_75t_L g1704 ( 
.A1(n_1687),
.A2(n_1645),
.A3(n_1643),
.B1(n_1626),
.B2(n_1628),
.C1(n_1631),
.C2(n_1636),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1683),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1677),
.B(n_1690),
.C(n_1686),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1684),
.A2(n_1632),
.B1(n_1628),
.B2(n_1631),
.Y(n_1707)
);

AOI322xp5_ASAP7_75t_L g1708 ( 
.A1(n_1695),
.A2(n_1645),
.A3(n_1643),
.B1(n_1636),
.B2(n_1553),
.C1(n_1589),
.C2(n_1606),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1696),
.A2(n_1639),
.B(n_1480),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1699),
.B(n_1689),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1711)
);

AOI211x1_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1702),
.B(n_1703),
.C(n_1706),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1707),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1701),
.Y(n_1714)
);

NAND4xp25_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1691),
.C(n_1689),
.D(n_1697),
.Y(n_1715)
);

NAND4xp25_ASAP7_75t_L g1716 ( 
.A(n_1709),
.B(n_1693),
.C(n_1681),
.D(n_1685),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1708),
.Y(n_1717)
);

NAND5xp2_ASAP7_75t_L g1718 ( 
.A(n_1704),
.B(n_1685),
.C(n_1497),
.D(n_1300),
.E(n_1463),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1705),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1712),
.A2(n_1685),
.B(n_1638),
.C(n_1622),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1716),
.B(n_1715),
.C(n_1711),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_SL g1722 ( 
.A(n_1719),
.B(n_1639),
.C(n_1638),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1714),
.B(n_1638),
.C(n_1622),
.Y(n_1723)
);

NAND5xp2_ASAP7_75t_L g1724 ( 
.A(n_1718),
.B(n_1713),
.C(n_1717),
.D(n_1710),
.E(n_1423),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1712),
.B(n_1641),
.C(n_1622),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1722),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_L g1727 ( 
.A(n_1725),
.B(n_1641),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1720),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1723),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1721),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1724),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1730),
.B(n_1641),
.Y(n_1732)
);

BUFx12f_ASAP7_75t_L g1733 ( 
.A(n_1729),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1726),
.A2(n_1611),
.B1(n_1585),
.B2(n_1599),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1726),
.B(n_1599),
.Y(n_1735)
);

OAI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1731),
.A2(n_1611),
.B(n_1596),
.Y(n_1736)
);

XNOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1732),
.B(n_1728),
.Y(n_1737)
);

AND2x2_ASAP7_75t_SL g1738 ( 
.A(n_1735),
.B(n_1727),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1735),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1738),
.Y(n_1740)
);

NOR4xp25_ASAP7_75t_L g1741 ( 
.A(n_1740),
.B(n_1739),
.C(n_1736),
.D(n_1737),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1741),
.Y(n_1742)
);

OAI22x1_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1733),
.B1(n_1734),
.B2(n_1595),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1606),
.B1(n_1598),
.B2(n_1596),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1743),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1745),
.B(n_1744),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1598),
.B(n_1556),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1746),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_R g1749 ( 
.A1(n_1748),
.A2(n_1747),
.B1(n_1549),
.B2(n_1540),
.C(n_1551),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1565),
.B1(n_1540),
.B2(n_1545),
.C(n_1549),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1274),
.B(n_1334),
.C(n_1322),
.Y(n_1751)
);


endmodule