module fake_jpeg_3154_n_707 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_707);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_707;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_7),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_61),
.Y(n_179)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_87),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_67),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_72),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_73),
.Y(n_184)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_21),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_99),
.Y(n_141)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_18),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_95),
.B(n_44),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_43),
.B(n_17),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_43),
.B(n_49),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_132),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx4f_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_49),
.B(n_17),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_50),
.B1(n_28),
.B2(n_39),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_150),
.B(n_123),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_72),
.A2(n_39),
.B1(n_50),
.B2(n_28),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_157),
.A2(n_195),
.B1(n_206),
.B2(n_207),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_65),
.A2(n_50),
.B1(n_39),
.B2(n_28),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_161),
.A2(n_176),
.B1(n_225),
.B2(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_174),
.B(n_192),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_68),
.A2(n_50),
.B1(n_36),
.B2(n_46),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_97),
.B(n_44),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_183),
.B(n_190),
.Y(n_282)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_121),
.B(n_36),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_100),
.B(n_46),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_112),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_117),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_117),
.A2(n_53),
.B1(n_42),
.B2(n_41),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_210),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_83),
.B(n_53),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_212),
.B(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_213),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_81),
.B(n_22),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_110),
.B(n_42),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_113),
.B(n_41),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_227),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_76),
.A2(n_70),
.B1(n_73),
.B2(n_88),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_93),
.B(n_30),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_134),
.B(n_33),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_82),
.B(n_85),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_130),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_101),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_111),
.A2(n_27),
.B1(n_22),
.B2(n_17),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_146),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_233),
.B(n_245),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_234),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_176),
.A2(n_108),
.B1(n_96),
.B2(n_104),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_235),
.A2(n_243),
.B1(n_268),
.B2(n_184),
.Y(n_344)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_236),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_183),
.A2(n_94),
.B(n_105),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_238),
.A2(n_266),
.B(n_288),
.Y(n_379)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_136),
.A2(n_115),
.B1(n_131),
.B2(n_126),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_246),
.B(n_250),
.Y(n_322)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_247),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_248),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_150),
.Y(n_249)
);

BUFx24_ASAP7_75t_L g357 ( 
.A(n_249),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_164),
.B(n_125),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_254),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_257),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_256),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_203),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_152),
.B(n_0),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_287),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_260),
.Y(n_356)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_261),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_218),
.A2(n_102),
.B1(n_16),
.B2(n_15),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_157),
.A2(n_14),
.B(n_13),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_269),
.A2(n_230),
.B(n_191),
.C(n_172),
.Y(n_336)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_162),
.Y(n_270)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_271),
.A2(n_276),
.B1(n_289),
.B2(n_291),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_141),
.A2(n_14),
.B1(n_13),
.B2(n_5),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_164),
.B(n_13),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_278),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_203),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_281),
.Y(n_345)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_215),
.Y(n_285)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_189),
.Y(n_286)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_141),
.B(n_1),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_139),
.B(n_4),
.C(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_295),
.C(n_307),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_140),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_160),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_148),
.B(n_7),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_304),
.Y(n_347)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_186),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_144),
.B(n_9),
.C(n_10),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_221),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_300),
.B1(n_256),
.B2(n_301),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_195),
.A2(n_231),
.B1(n_207),
.B2(n_206),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_298),
.A2(n_299),
.B1(n_303),
.B2(n_314),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_193),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_200),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_179),
.Y(n_301)
);

OR2x6_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_205),
.Y(n_320)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_302),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_142),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_151),
.B(n_12),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_142),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_305),
.B(n_308),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_154),
.B(n_12),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_147),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_143),
.B(n_145),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_309),
.B(n_315),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_229),
.A2(n_216),
.B1(n_149),
.B2(n_193),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_191),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_159),
.A2(n_217),
.B(n_199),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_223),
.C(n_166),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_167),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_313),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_175),
.A2(n_197),
.B1(n_155),
.B2(n_177),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_205),
.B(n_179),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_180),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_316),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_320),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_249),
.A2(n_184),
.B1(n_177),
.B2(n_138),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g422 ( 
.A1(n_325),
.A2(n_336),
.B1(n_344),
.B2(n_320),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_237),
.B(n_208),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_327),
.B(n_265),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_363),
.C(n_379),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_239),
.B(n_211),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_361),
.C(n_301),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_153),
.B(n_168),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_275),
.B(n_281),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_239),
.B(n_307),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_264),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_272),
.B(n_182),
.C(n_211),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_267),
.A2(n_228),
.B1(n_185),
.B2(n_181),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_240),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_SL g365 ( 
.A(n_287),
.B(n_181),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_SL g419 ( 
.A(n_365),
.B(n_316),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_SL g366 ( 
.A(n_268),
.B(n_194),
.C(n_147),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_SL g416 ( 
.A(n_366),
.B(n_270),
.C(n_279),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_238),
.A2(n_194),
.B1(n_282),
.B2(n_241),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_373),
.B1(n_378),
.B2(n_308),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_256),
.A2(n_235),
.B1(n_306),
.B2(n_236),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_370),
.A2(n_280),
.B1(n_286),
.B2(n_260),
.Y(n_413)
);

OA22x2_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_306),
.B1(n_269),
.B2(n_291),
.Y(n_371)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_258),
.A2(n_245),
.B1(n_304),
.B2(n_292),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_266),
.A2(n_306),
.B1(n_284),
.B2(n_312),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_295),
.B(n_297),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g446 ( 
.A1(n_383),
.A2(n_397),
.B(n_401),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_384),
.B(n_385),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_358),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_386),
.B(n_394),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_234),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_387),
.B(n_388),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_327),
.B(n_242),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_263),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_399),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_390),
.A2(n_413),
.B(n_331),
.Y(n_450)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_416),
.Y(n_461)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_378),
.B(n_317),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_396),
.B(n_326),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_333),
.B(n_274),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_403),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_244),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_305),
.B1(n_290),
.B2(n_293),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_400),
.A2(n_408),
.B1(n_409),
.B2(n_320),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_273),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_320),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_360),
.B(n_253),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_415),
.Y(n_453)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_332),
.B1(n_371),
.B2(n_363),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_359),
.A2(n_294),
.B1(n_310),
.B2(n_259),
.Y(n_409)
);

OR2x2_ASAP7_75t_SL g410 ( 
.A(n_365),
.B(n_251),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_L g470 ( 
.A1(n_410),
.A2(n_353),
.B(n_345),
.Y(n_470)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_252),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_318),
.C(n_361),
.Y(n_437)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_322),
.B(n_247),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_283),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_343),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_336),
.B(n_357),
.Y(n_441)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_420),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_364),
.A2(n_261),
.B1(n_254),
.B2(n_248),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_422),
.B1(n_427),
.B2(n_371),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_426),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_285),
.B1(n_313),
.B2(n_302),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_425),
.A2(n_376),
.B1(n_320),
.B2(n_331),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_344),
.A2(n_316),
.B1(n_371),
.B2(n_357),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_318),
.B(n_328),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_324),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_429),
.B(n_348),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_418),
.A2(n_357),
.B(n_321),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_463),
.B(n_468),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_462),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_438),
.A2(n_427),
.B1(n_421),
.B2(n_395),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_351),
.C(n_328),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_447),
.C(n_415),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_441),
.A2(n_443),
.B(n_450),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_469),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_380),
.A2(n_321),
.B1(n_320),
.B2(n_376),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_445),
.A2(n_449),
.B1(n_452),
.B2(n_467),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_324),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_382),
.A2(n_366),
.B1(n_372),
.B2(n_341),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_472),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_382),
.A2(n_372),
.B1(n_341),
.B2(n_362),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_382),
.A2(n_362),
.B1(n_335),
.B2(n_329),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_343),
.B(n_330),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_459),
.A2(n_418),
.B(n_424),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_403),
.A2(n_408),
.B(n_419),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_464),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_335),
.B1(n_337),
.B2(n_348),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_381),
.A2(n_345),
.B(n_369),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_470),
.A2(n_471),
.B(n_409),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_381),
.A2(n_375),
.B(n_330),
.Y(n_471)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_473),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_451),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_474),
.B(n_486),
.Y(n_515)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_430),
.Y(n_476)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_430),
.Y(n_478)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_479),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_480),
.A2(n_496),
.B(n_498),
.Y(n_530)
);

OAI22x1_ASAP7_75t_L g525 ( 
.A1(n_481),
.A2(n_455),
.B1(n_441),
.B2(n_468),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_445),
.A2(n_395),
.B1(n_410),
.B2(n_400),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_504),
.Y(n_524)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

AOI32xp33_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_388),
.A3(n_395),
.B1(n_410),
.B2(n_402),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_451),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_458),
.Y(n_516)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_436),
.Y(n_490)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_490),
.Y(n_523)
);

XOR2x1_ASAP7_75t_SL g491 ( 
.A(n_463),
.B(n_383),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_SL g545 ( 
.A1(n_491),
.A2(n_495),
.B(n_466),
.Y(n_545)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_439),
.Y(n_494)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_416),
.Y(n_495)
);

A2O1A1O1Ixp25_ASAP7_75t_L g496 ( 
.A1(n_440),
.A2(n_385),
.B(n_404),
.C(n_399),
.D(n_389),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_439),
.Y(n_497)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_437),
.B(n_384),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_507),
.Y(n_521)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_500),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_437),
.B(n_417),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_502),
.C(n_505),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_438),
.A2(n_387),
.B1(n_397),
.B2(n_401),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_461),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_431),
.B(n_391),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_462),
.B(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_506),
.B(n_508),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_440),
.B(n_405),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_426),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_434),
.A2(n_390),
.B1(n_407),
.B2(n_414),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_434),
.B(n_420),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_511),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_461),
.A2(n_390),
.B1(n_411),
.B2(n_398),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_369),
.C(n_326),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_447),
.C(n_454),
.Y(n_541)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_516),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_504),
.B(n_453),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_520),
.B(n_532),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_525),
.A2(n_528),
.B1(n_538),
.B2(n_546),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_481),
.A2(n_461),
.B1(n_469),
.B2(n_435),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_489),
.B(n_453),
.Y(n_529)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_508),
.B(n_446),
.Y(n_531)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_510),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_533),
.A2(n_537),
.B(n_480),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_477),
.Y(n_535)
);

INVx13_ASAP7_75t_L g567 ( 
.A(n_535),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_484),
.A2(n_455),
.B(n_433),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_503),
.A2(n_477),
.B1(n_488),
.B2(n_495),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_542),
.C(n_491),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_454),
.C(n_447),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_464),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_543),
.B(n_484),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_477),
.A2(n_459),
.B1(n_452),
.B2(n_449),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_544),
.A2(n_547),
.B1(n_492),
.B2(n_490),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_545),
.B(n_493),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_488),
.A2(n_443),
.B1(n_466),
.B2(n_448),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_475),
.A2(n_467),
.B1(n_433),
.B2(n_458),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_495),
.A2(n_450),
.B1(n_456),
.B2(n_457),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_498),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_499),
.B(n_507),
.Y(n_549)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_511),
.B(n_457),
.Y(n_550)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_550),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_552),
.B(n_560),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_501),
.C(n_502),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_557),
.C(n_565),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_512),
.C(n_505),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_558),
.B(n_571),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_561),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_483),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_524),
.A2(n_493),
.B1(n_496),
.B2(n_497),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_562),
.A2(n_569),
.B1(n_570),
.B2(n_550),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_506),
.C(n_500),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_479),
.C(n_476),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_566),
.B(n_572),
.C(n_579),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_524),
.A2(n_478),
.B1(n_494),
.B2(n_456),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_536),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_472),
.C(n_465),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_537),
.A2(n_442),
.B(n_460),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_573),
.B(n_576),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_334),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_574),
.B(n_575),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_530),
.B(n_334),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_535),
.A2(n_386),
.B(n_394),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_576),
.B(n_577),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_551),
.A2(n_473),
.B(n_460),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_406),
.C(n_353),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_531),
.B(n_367),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_582),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_538),
.B(n_423),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g583 ( 
.A1(n_551),
.A2(n_423),
.B(n_356),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_514),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_533),
.B(n_406),
.C(n_356),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_584),
.B(n_585),
.C(n_544),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_337),
.C(n_367),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_515),
.B(n_323),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_586),
.B(n_539),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_589),
.A2(n_602),
.B1(n_613),
.B2(n_567),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_520),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_591),
.B(n_600),
.Y(n_626)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_564),
.Y(n_594)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_594),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_554),
.B(n_563),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_598),
.B(n_604),
.Y(n_617)
);

FAx1_ASAP7_75t_SL g600 ( 
.A(n_562),
.B(n_528),
.CI(n_558),
.CON(n_600),
.SN(n_600)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_601),
.B(n_607),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_580),
.A2(n_546),
.B1(n_547),
.B2(n_568),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_568),
.A2(n_532),
.B1(n_522),
.B2(n_529),
.Y(n_603)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_603),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_556),
.B(n_548),
.C(n_525),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_605),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_565),
.B(n_536),
.C(n_527),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_606),
.B(n_574),
.C(n_585),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_527),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_567),
.Y(n_634)
);

FAx1_ASAP7_75t_SL g609 ( 
.A(n_559),
.B(n_539),
.CI(n_513),
.CON(n_609),
.SN(n_609)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_609),
.B(n_614),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_566),
.B(n_519),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_610),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_611),
.A2(n_583),
.B(n_577),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_572),
.B(n_519),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_581),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_555),
.A2(n_518),
.B1(n_513),
.B2(n_514),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_592),
.A2(n_573),
.B(n_553),
.Y(n_615)
);

OAI21x1_ASAP7_75t_SL g654 ( 
.A1(n_615),
.A2(n_627),
.B(n_635),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_619),
.B(n_622),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_613),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_635),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_552),
.C(n_561),
.Y(n_622)
);

BUFx24_ASAP7_75t_SL g623 ( 
.A(n_609),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_623),
.B(n_632),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_588),
.B(n_579),
.C(n_584),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_625),
.B(n_628),
.C(n_629),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_588),
.B(n_582),
.C(n_575),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_586),
.C(n_560),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_526),
.Y(n_630)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_630),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_631),
.A2(n_587),
.B1(n_614),
.B2(n_607),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_634),
.B(n_638),
.C(n_597),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_603),
.B(n_518),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_590),
.B(n_523),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_597),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_523),
.C(n_526),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_641),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_626),
.A2(n_589),
.B1(n_602),
.B2(n_599),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_616),
.B(n_601),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_642),
.B(n_648),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_SL g644 ( 
.A(n_627),
.B(n_590),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_644),
.B(n_658),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_620),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_638),
.C(n_619),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_626),
.B(n_599),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_649),
.B(n_650),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_604),
.C(n_587),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_624),
.B(n_517),
.Y(n_651)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_651),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_652),
.A2(n_654),
.B1(n_633),
.B2(n_621),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_517),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_653),
.B(n_655),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_617),
.B(n_593),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_630),
.B(n_534),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_656),
.A2(n_615),
.B(n_618),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_659),
.B(n_664),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_660),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_620),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_SL g680 ( 
.A(n_663),
.B(n_659),
.Y(n_680)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_650),
.B(n_628),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_665),
.B(n_657),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_646),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_666),
.B(n_667),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_637),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_640),
.B(n_637),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_674),
.Y(n_677)
);

XOR2xp5_ASAP7_75t_L g669 ( 
.A(n_647),
.B(n_636),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_669),
.B(n_673),
.Y(n_678)
);

XOR2xp5_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_631),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_671),
.B(n_661),
.Y(n_679)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_680),
.A2(n_681),
.B(n_658),
.Y(n_687)
);

NOR2x1_ASAP7_75t_SL g681 ( 
.A(n_663),
.B(n_657),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_682),
.B(n_684),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_670),
.B(n_654),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_686),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_664),
.B(n_640),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_669),
.B(n_622),
.C(n_633),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_687),
.A2(n_688),
.B(n_691),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_685),
.A2(n_677),
.B(n_675),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_685),
.A2(n_676),
.B(n_686),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_678),
.B(n_662),
.Y(n_693)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_693),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_675),
.A2(n_674),
.B(n_656),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_694),
.A2(n_645),
.B(n_652),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_672),
.Y(n_696)
);

OAI21x1_ASAP7_75t_SL g702 ( 
.A1(n_696),
.A2(n_697),
.B(n_534),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_689),
.B(n_645),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g701 ( 
.A1(n_698),
.A2(n_629),
.B(n_673),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_699),
.A2(n_692),
.B(n_690),
.Y(n_700)
);

OAI321xp33_ASAP7_75t_L g704 ( 
.A1(n_700),
.A2(n_701),
.A3(n_600),
.B1(n_595),
.B2(n_593),
.C(n_340),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_702),
.A2(n_695),
.B(n_609),
.Y(n_703)
);

BUFx24_ASAP7_75t_SL g705 ( 
.A(n_703),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_705),
.B(n_704),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_706),
.A2(n_600),
.B(n_595),
.Y(n_707)
);


endmodule