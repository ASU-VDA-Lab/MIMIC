module fake_jpeg_20172_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_15),
.B1(n_33),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_53),
.B1(n_29),
.B2(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_15),
.B1(n_33),
.B2(n_16),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_31),
.B1(n_19),
.B2(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_64),
.B1(n_25),
.B2(n_24),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_57),
.B1(n_42),
.B2(n_38),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_104),
.B(n_3),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_70),
.B(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_73),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_32),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_84),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_39),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_44),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_87),
.B1(n_98),
.B2(n_62),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_37),
.B1(n_20),
.B2(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_106),
.B1(n_0),
.B2(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_13),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_97),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_31),
.B1(n_19),
.B2(n_2),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_19),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_1),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_62),
.B1(n_5),
.B2(n_2),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_5),
.C(n_11),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_112),
.C(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_117),
.B1(n_132),
.B2(n_119),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_5),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_84),
.B(n_99),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_4),
.B(n_8),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_106),
.B(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_10),
.B1(n_12),
.B2(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_101),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_10),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_10),
.C(n_12),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_160),
.B(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_147),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_138),
.C(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_121),
.B1(n_110),
.B2(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_100),
.B1(n_113),
.B2(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_74),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_108),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_91),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_121),
.B1(n_114),
.B2(n_122),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_159),
.B1(n_108),
.B2(n_123),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_105),
.B1(n_95),
.B2(n_71),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_89),
.B(n_90),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_88),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_165),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_95),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_71),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_127),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_119),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_182),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_120),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_151),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_159),
.B1(n_146),
.B2(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_131),
.B(n_100),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_192),
.B1(n_181),
.B2(n_171),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_162),
.C(n_146),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_200),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_145),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_146),
.C(n_164),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_164),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.C(n_186),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_141),
.C(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_161),
.B1(n_141),
.B2(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_178),
.B1(n_172),
.B2(n_166),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_216),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_200),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_184),
.B1(n_161),
.B2(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_211),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_196),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_168),
.B1(n_171),
.B2(n_182),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_212),
.Y(n_227)
);

FAx1_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_175),
.CI(n_167),
.CON(n_213),
.SN(n_213)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_194),
.B(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_185),
.B1(n_166),
.B2(n_178),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_192),
.B1(n_197),
.B2(n_194),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_168),
.B1(n_173),
.B2(n_170),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_170),
.A3(n_180),
.B1(n_154),
.B2(n_183),
.C1(n_157),
.C2(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_193),
.C(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.C(n_215),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_202),
.C(n_190),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_217),
.B(n_209),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_154),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_236),
.B(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_217),
.B(n_213),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_213),
.B(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_229),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_218),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_219),
.B(n_225),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_225),
.B1(n_227),
.B2(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_218),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_215),
.B(n_228),
.C(n_243),
.D(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_250),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_252),
.B1(n_254),
.B2(n_241),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_259),
.A2(n_257),
.B(n_226),
.C(n_150),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_131),
.Y(n_261)
);


endmodule