module fake_jpeg_5157_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_39),
.B(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_7),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_44),
.B(n_50),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_52),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_10),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_17),
.Y(n_70)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_28),
.B1(n_16),
.B2(n_18),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_37),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_71),
.B1(n_96),
.B2(n_98),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_69),
.B(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_27),
.B1(n_37),
.B2(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_27),
.B(n_19),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_91),
.B(n_17),
.Y(n_109)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_79),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_90),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_33),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_97),
.Y(n_112)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_16),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_18),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_1),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_26),
.B1(n_35),
.B2(n_32),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_42),
.A2(n_35),
.B1(n_29),
.B2(n_20),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_17),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_29),
.B1(n_32),
.B2(n_20),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_111),
.B1(n_115),
.B2(n_117),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_125),
.B(n_92),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_22),
.B1(n_17),
.B2(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_22),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_122),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_8),
.B1(n_13),
.B2(n_3),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_126),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_68),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_128),
.B1(n_68),
.B2(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_2),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_4),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_9),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_63),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_98),
.B1(n_60),
.B2(n_85),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_58),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_144),
.C(n_106),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_145),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_125),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_147),
.B1(n_157),
.B2(n_141),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_106),
.B(n_112),
.Y(n_166)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_140),
.Y(n_184)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_143),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_84),
.C(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_59),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_160),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_153),
.B1(n_155),
.B2(n_157),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_84),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_156),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_69),
.B1(n_66),
.B2(n_73),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_111),
.B1(n_120),
.B2(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_73),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_75),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_110),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_80),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_67),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_62),
.CI(n_59),
.CON(n_164),
.SN(n_164)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_135),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_169),
.B(n_159),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_177),
.CI(n_180),
.CON(n_198),
.SN(n_198)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_188),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_132),
.B1(n_119),
.B2(n_121),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_127),
.B1(n_114),
.B2(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_114),
.B(n_120),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_104),
.B1(n_108),
.B2(n_65),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_62),
.C(n_67),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_136),
.C(n_155),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_108),
.B1(n_131),
.B2(n_65),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_12),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_93),
.B1(n_15),
.B2(n_13),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_145),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_211),
.B(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_204),
.C(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_164),
.C(n_143),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_180),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_167),
.A2(n_139),
.B1(n_140),
.B2(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_162),
.C(n_131),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_166),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_175),
.C(n_177),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_165),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_171),
.B1(n_170),
.B2(n_178),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_186),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_224),
.C(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_191),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_196),
.B(n_199),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_190),
.A3(n_182),
.B1(n_169),
.B2(n_173),
.Y(n_227)
);

AOI321xp33_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_230),
.A3(n_205),
.B1(n_198),
.B2(n_213),
.C(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_172),
.C(n_169),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_173),
.C(n_189),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_214),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_223),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_208),
.B1(n_176),
.B2(n_204),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_208),
.B(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_222),
.B1(n_229),
.B2(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_232),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_246),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_237),
.B(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_218),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_220),
.C(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_242),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_223),
.C(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_238),
.C(n_245),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_254),
.CI(n_255),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_249),
.C(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_260),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_244),
.C(n_217),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_259),
.C(n_262),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_252),
.Y(n_265)
);


endmodule