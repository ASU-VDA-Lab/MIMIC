module fake_jpeg_29613_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_2),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_42),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_3),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_3),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_70),
.B1(n_24),
.B2(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_4),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_22),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_13),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_15),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_21),
.C(n_23),
.Y(n_85)
);

AO21x2_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_18),
.B(n_19),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_87),
.B1(n_65),
.B2(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_26),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_91),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_83),
.B(n_66),
.C(n_82),
.D(n_86),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_86),
.C(n_82),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_79),
.C(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_84),
.C(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_97),
.C(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_79),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

AOI21x1_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_88),
.B(n_29),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_27),
.Y(n_103)
);


endmodule