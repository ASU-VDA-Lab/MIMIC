module fake_aes_8247_n_29 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_6), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g11 ( .A(n_7), .B(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_0), .B(n_1), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_SL g19 ( .A1(n_14), .A2(n_0), .B(n_2), .C(n_3), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_16), .B(n_14), .Y(n_20) );
AO31x2_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_15), .A3(n_14), .B(n_11), .Y(n_21) );
NOR2xp67_ASAP7_75t_R g22 ( .A(n_18), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_12), .C(n_10), .Y(n_25) );
A2O1A1Ixp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_23), .B(n_24), .C(n_15), .Y(n_26) );
AOI222xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_22), .B1(n_18), .B2(n_19), .C1(n_21), .C2(n_4), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B1(n_22), .B2(n_7), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_18), .B1(n_6), .B2(n_8), .Y(n_29) );
endmodule