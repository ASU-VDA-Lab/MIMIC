module fake_jpeg_1046_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_0),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_17),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_15),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_0),
.B(n_3),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_36),
.B1(n_37),
.B2(n_17),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_73),
.B1(n_84),
.B2(n_86),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_21),
.B1(n_29),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_75),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_36),
.B1(n_30),
.B2(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_87),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_16),
.B1(n_23),
.B2(n_19),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_41),
.A2(n_38),
.B1(n_24),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_26),
.B1(n_34),
.B2(n_18),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_98),
.B1(n_108),
.B2(n_110),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_24),
.B1(n_40),
.B2(n_38),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_99),
.B1(n_107),
.B2(n_7),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_31),
.B1(n_28),
.B2(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_26),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_9),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_31),
.B1(n_28),
.B2(n_22),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_31),
.B1(n_28),
.B2(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_0),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_48),
.A2(n_39),
.B1(n_1),
.B2(n_3),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_39),
.B1(n_32),
.B2(n_8),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_32),
.B1(n_14),
.B2(n_11),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_51),
.A2(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_128),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_123),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_0),
.B(n_3),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_125),
.B(n_145),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_121),
.B(n_127),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_67),
.B(n_5),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_32),
.B1(n_8),
.B2(n_10),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_137),
.B(n_77),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_7),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_76),
.B1(n_106),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_110),
.B1(n_102),
.B2(n_66),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_77),
.B1(n_83),
.B2(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

AO22x2_ASAP7_75t_L g137 ( 
.A1(n_69),
.A2(n_90),
.B1(n_79),
.B2(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_68),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_70),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_66),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_69),
.A2(n_68),
.B(n_82),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_152),
.B1(n_148),
.B2(n_126),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_79),
.B1(n_88),
.B2(n_76),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_101),
.C(n_93),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_181),
.C(n_143),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_100),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_159),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_109),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_119),
.B(n_117),
.C(n_121),
.D(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_109),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_134),
.B1(n_131),
.B2(n_137),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_109),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_83),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_147),
.Y(n_212)
);

CKINVDCx10_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_106),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_132),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_130),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_204),
.B1(n_162),
.B2(n_149),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_190),
.A2(n_220),
.B(n_186),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_199),
.Y(n_248)
);

NOR2x1p5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_216),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_162),
.B1(n_173),
.B2(n_175),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_125),
.B1(n_137),
.B2(n_123),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_147),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_130),
.Y(n_210)
);

AOI31xp33_ASAP7_75t_SL g249 ( 
.A1(n_210),
.A2(n_218),
.A3(n_190),
.B(n_220),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_213),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_144),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_151),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_158),
.B(n_113),
.C(n_144),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_176),
.A2(n_179),
.B(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_146),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_162),
.B1(n_160),
.B2(n_173),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_195),
.B1(n_187),
.B2(n_193),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_228),
.A2(n_201),
.B1(n_214),
.B2(n_222),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_155),
.C(n_161),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_235),
.C(n_213),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_161),
.C(n_173),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_195),
.A2(n_185),
.B1(n_165),
.B2(n_184),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_239),
.B(n_247),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_168),
.B(n_171),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_209),
.A2(n_151),
.B(n_154),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_211),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_154),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_204),
.A2(n_194),
.B1(n_207),
.B2(n_203),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_253),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_245),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_231),
.B(n_247),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_269),
.C(n_230),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_258),
.Y(n_286)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_227),
.B1(n_250),
.B2(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_272),
.B1(n_229),
.B2(n_228),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_191),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_268),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_218),
.B1(n_194),
.B2(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_244),
.B1(n_229),
.B2(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_212),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_200),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_234),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_265),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_282),
.C(n_289),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_248),
.C(n_235),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_233),
.B1(n_225),
.B2(n_246),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_251),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_246),
.B1(n_239),
.B2(n_216),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_243),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_243),
.C(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_243),
.C(n_189),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_266),
.C(n_257),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_262),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_300),
.Y(n_313)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_262),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_SL g300 ( 
.A(n_274),
.B(n_271),
.C(n_268),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_236),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_271),
.C(n_263),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_282),
.C(n_290),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_291),
.A2(n_278),
.B(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_307),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_289),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_253),
.B1(n_252),
.B2(n_258),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_316),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_267),
.B1(n_261),
.B2(n_264),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_299),
.B(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_261),
.B1(n_238),
.B2(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_301),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_324),
.B1(n_314),
.B2(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_297),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_293),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_312),
.B(n_309),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_327),
.B(n_306),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_307),
.B(n_311),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_298),
.C(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_288),
.B1(n_303),
.B2(n_272),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_306),
.C(n_321),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_321),
.B(n_319),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_328),
.A3(n_198),
.B1(n_202),
.B2(n_189),
.C1(n_219),
.C2(n_205),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_198),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_198),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_336),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_205),
.Y(n_341)
);


endmodule