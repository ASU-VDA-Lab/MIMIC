module fake_jpeg_13572_n_497 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_3),
.B(n_4),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_64),
.Y(n_132)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_65),
.B(n_75),
.Y(n_167)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_66),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_10),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_10),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_68),
.B(n_71),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_17),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_76),
.B(n_80),
.Y(n_147)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_8),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_11),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_82),
.B(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_22),
.B(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_11),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_26),
.B(n_17),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_100),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_91),
.Y(n_188)
);

BUFx6f_ASAP7_75t_SL g92 ( 
.A(n_28),
.Y(n_92)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_28),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_94),
.Y(n_191)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_26),
.B(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx3_ASAP7_75t_SL g104 ( 
.A(n_56),
.Y(n_104)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_109),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g109 ( 
.A(n_56),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_25),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_113),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_35),
.Y(n_111)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_27),
.B(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_19),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g121 ( 
.A(n_50),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_56),
.B(n_42),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_41),
.C(n_56),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_124),
.B(n_146),
.C(n_186),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_58),
.B1(n_52),
.B2(n_40),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_127),
.A2(n_137),
.B1(n_157),
.B2(n_160),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_65),
.A2(n_18),
.B1(n_51),
.B2(n_59),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_133),
.A2(n_154),
.B1(n_159),
.B2(n_163),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_40),
.B1(n_58),
.B2(n_52),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_111),
.C(n_95),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_72),
.A2(n_18),
.B1(n_51),
.B2(n_40),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_150),
.A2(n_173),
.B1(n_177),
.B2(n_194),
.Y(n_229)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_151),
.B(n_191),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_69),
.A2(n_51),
.B1(n_58),
.B2(n_35),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_34),
.B1(n_49),
.B2(n_48),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_94),
.A2(n_35),
.B1(n_43),
.B2(n_38),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_61),
.A2(n_53),
.B1(n_43),
.B2(n_38),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_30),
.B1(n_53),
.B2(n_25),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_74),
.A2(n_112),
.B1(n_83),
.B2(n_79),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_164),
.A2(n_168),
.B1(n_183),
.B2(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_66),
.B(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_182),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_105),
.A2(n_32),
.B1(n_49),
.B2(n_48),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_78),
.A2(n_29),
.B1(n_47),
.B2(n_34),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_176),
.B1(n_181),
.B2(n_186),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_84),
.A2(n_57),
.B1(n_47),
.B2(n_29),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_91),
.A2(n_32),
.B1(n_57),
.B2(n_42),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_106),
.A2(n_42),
.B1(n_50),
.B2(n_19),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_119),
.A2(n_19),
.B1(n_1),
.B2(n_0),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_102),
.B(n_0),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_60),
.A2(n_4),
.B1(n_13),
.B2(n_14),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_120),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_60),
.A2(n_13),
.B1(n_0),
.B2(n_1),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_104),
.B(n_0),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_167),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_104),
.A2(n_1),
.B1(n_63),
.B2(n_116),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_104),
.B1(n_121),
.B2(n_99),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g262 ( 
.A1(n_195),
.A2(n_213),
.B(n_252),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_121),
.B1(n_1),
.B2(n_96),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_196),
.A2(n_223),
.B1(n_249),
.B2(n_252),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_197),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_136),
.B(n_1),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_198),
.B(n_206),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_199),
.B(n_230),
.Y(n_295)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_203),
.B(n_217),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_146),
.B1(n_177),
.B2(n_124),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_205),
.A2(n_242),
.B1(n_251),
.B2(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_138),
.B(n_180),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_207),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_167),
.B(n_134),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_209),
.A2(n_238),
.B(n_244),
.Y(n_310)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_144),
.A2(n_182),
.B1(n_126),
.B2(n_147),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_211),
.A2(n_245),
.B1(n_256),
.B2(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_212),
.B(n_215),
.Y(n_278)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_122),
.B1(n_170),
.B2(n_166),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_184),
.Y(n_215)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_130),
.B(n_153),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_218),
.B(n_225),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_143),
.Y(n_221)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_127),
.A2(n_144),
.B1(n_126),
.B2(n_179),
.Y(n_223)
);

OR2x2_ASAP7_75t_SL g224 ( 
.A(n_123),
.B(n_125),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_132),
.B(n_169),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_170),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_227),
.Y(n_296)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_143),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_233),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g232 ( 
.A(n_141),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_232),
.Y(n_286)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

CKINVDCx12_ASAP7_75t_R g234 ( 
.A(n_140),
.Y(n_234)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_234),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_162),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_239),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_123),
.B(n_125),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_236),
.B(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_178),
.A2(n_172),
.B(n_128),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_129),
.B(n_148),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_129),
.B(n_148),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_149),
.B(n_152),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_140),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_246),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_149),
.A2(n_152),
.B(n_156),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_155),
.A2(n_179),
.B1(n_156),
.B2(n_188),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_145),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_248),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_141),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_193),
.A2(n_155),
.B1(n_189),
.B2(n_145),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_135),
.B(n_189),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_161),
.B(n_178),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_193),
.B1(n_139),
.B2(n_172),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_161),
.B(n_139),
.Y(n_253)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_254),
.A2(n_239),
.B1(n_232),
.B2(n_214),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_138),
.A2(n_146),
.B1(n_144),
.B2(n_182),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_180),
.B(n_147),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_257),
.A2(n_225),
.B1(n_251),
.B2(n_253),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_146),
.A2(n_165),
.B(n_167),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_212),
.B(n_204),
.C(n_217),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_136),
.B(n_153),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_259),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_204),
.B(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_266),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_262),
.A2(n_235),
.B(n_216),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_263),
.A2(n_282),
.B(n_278),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_219),
.B1(n_202),
.B2(n_208),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_267),
.A2(n_288),
.B1(n_234),
.B2(n_257),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_270),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_271),
.B(n_265),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_277),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_237),
.Y(n_277)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_203),
.A2(n_219),
.B1(n_213),
.B2(n_229),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_291),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_202),
.A2(n_255),
.B1(n_195),
.B2(n_213),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_227),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_245),
.A2(n_201),
.B1(n_207),
.B2(n_218),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_292),
.A2(n_308),
.B1(n_286),
.B2(n_291),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_199),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_280),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_228),
.A2(n_233),
.B1(n_221),
.B2(n_210),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_325),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_238),
.C(n_246),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_318),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_231),
.B1(n_232),
.B2(n_248),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_313),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_315),
.A2(n_336),
.B1(n_343),
.B2(n_264),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_316),
.A2(n_326),
.B(n_312),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_269),
.B1(n_267),
.B2(n_287),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_317),
.A2(n_334),
.B(n_335),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_197),
.C(n_254),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_197),
.C(n_200),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_324),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_197),
.C(n_220),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_310),
.A2(n_220),
.B(n_269),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_348),
.B(n_346),
.Y(n_362)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g328 ( 
.A1(n_261),
.A2(n_220),
.A3(n_268),
.B1(n_263),
.B2(n_270),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_330),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_279),
.A2(n_282),
.B1(n_260),
.B2(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_279),
.B1(n_260),
.B2(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_278),
.B(n_293),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_342),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_293),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_282),
.A2(n_262),
.B(n_295),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_265),
.A2(n_262),
.B1(n_285),
.B2(n_309),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_307),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_345),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_306),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_338),
.B(n_347),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_341),
.A2(n_286),
.B1(n_273),
.B2(n_280),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_262),
.A2(n_300),
.B1(n_284),
.B2(n_275),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_306),
.A2(n_284),
.B1(n_296),
.B2(n_294),
.Y(n_343)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_303),
.B(n_296),
.C(n_272),
.D(n_274),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_346),
.A2(n_274),
.B(n_304),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_272),
.A2(n_273),
.B(n_274),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_350),
.A2(n_358),
.B(n_362),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_351),
.B(n_353),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_338),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_334),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_317),
.A2(n_264),
.B1(n_304),
.B2(n_305),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_357),
.A2(n_370),
.B1(n_377),
.B2(n_334),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_333),
.B(n_289),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_365),
.B(n_366),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_322),
.B(n_305),
.Y(n_366)
);

O2A1O1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_290),
.B(n_283),
.C(n_302),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_321),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_335),
.B(n_341),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_368),
.A2(n_374),
.B(n_312),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_322),
.B(n_302),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_371),
.B(n_372),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_302),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_290),
.B(n_264),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_314),
.A2(n_290),
.B1(n_313),
.B2(n_342),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_376),
.A2(n_318),
.B1(n_323),
.B2(n_324),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_330),
.A2(n_336),
.B1(n_315),
.B2(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_340),
.B(n_319),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_379),
.B(n_334),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_352),
.C(n_350),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_383),
.C(n_391),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_373),
.A2(n_325),
.B1(n_339),
.B2(n_332),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_381),
.A2(n_393),
.B1(n_370),
.B2(n_377),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_328),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_387),
.Y(n_408)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_340),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_388),
.A2(n_373),
.B1(n_386),
.B2(n_354),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_390),
.Y(n_409)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_339),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_344),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_396),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_398),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_356),
.A2(n_344),
.B(n_320),
.C(n_348),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_399),
.Y(n_417)
);

NOR4xp25_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_346),
.C(n_329),
.D(n_327),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_400),
.A2(n_367),
.B(n_368),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_366),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_403),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_369),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_352),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_412),
.C(n_413),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_418),
.B1(n_400),
.B2(n_355),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_352),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_361),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_350),
.C(n_361),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_421),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_373),
.B1(n_349),
.B2(n_376),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_422),
.Y(n_427)
);

AOI322xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_356),
.A3(n_364),
.B1(n_365),
.B2(n_360),
.C1(n_357),
.C2(n_371),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_360),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_356),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_389),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_367),
.B1(n_374),
.B2(n_357),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_426),
.B1(n_368),
.B2(n_362),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_389),
.A2(n_374),
.B1(n_355),
.B2(n_349),
.Y(n_426)
);

OAI321xp33_ASAP7_75t_L g428 ( 
.A1(n_411),
.A2(n_387),
.A3(n_385),
.B1(n_401),
.B2(n_392),
.C(n_402),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_432),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_422),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_425),
.Y(n_431)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_408),
.B(n_401),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_425),
.Y(n_433)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_437),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_411),
.B(n_403),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_416),
.B(n_364),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_443),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_384),
.Y(n_440)
);

AOI21x1_ASAP7_75t_SL g453 ( 
.A1(n_440),
.A2(n_382),
.B(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_414),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_418),
.B1(n_423),
.B2(n_400),
.Y(n_454)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_440),
.A2(n_419),
.B(n_409),
.Y(n_447)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_447),
.A2(n_437),
.B(n_358),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_454),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_407),
.C(n_405),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_457),
.Y(n_464)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_453),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_407),
.C(n_412),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_372),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_458),
.B(n_369),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_466),
.Y(n_470)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_467),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_462),
.B(n_428),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_449),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_432),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_439),
.C(n_444),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_469),
.Y(n_475)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_464),
.A2(n_449),
.B(n_447),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_474),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_473),
.A2(n_433),
.B(n_431),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_463),
.A2(n_435),
.B1(n_451),
.B2(n_429),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_455),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_476),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_478),
.C(n_453),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_463),
.A2(n_451),
.B1(n_446),
.B2(n_427),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_475),
.A2(n_468),
.B(n_455),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_480),
.C(n_481),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_466),
.C(n_454),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_483),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g485 ( 
.A1(n_472),
.A2(n_427),
.B(n_456),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g487 ( 
.A1(n_485),
.A2(n_358),
.A3(n_394),
.B1(n_398),
.B2(n_474),
.C1(n_382),
.C2(n_390),
.Y(n_487)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g486 ( 
.A1(n_483),
.A2(n_434),
.B(n_443),
.C(n_441),
.D(n_478),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_487),
.Y(n_493)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_484),
.A2(n_470),
.A3(n_400),
.B1(n_430),
.B2(n_406),
.C1(n_424),
.C2(n_417),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_489),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_488),
.A2(n_482),
.B(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_491),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_490),
.C(n_448),
.Y(n_495)
);

OAI31xp33_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_493),
.A3(n_415),
.B(n_426),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_494),
.C(n_421),
.Y(n_497)
);


endmodule