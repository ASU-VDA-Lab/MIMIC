module fake_netlist_1_9417_n_628 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_628);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_628;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_35), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_65), .Y(n_76) );
BUFx6f_ASAP7_75t_L g77 ( .A(n_46), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_70), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_68), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_67), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_73), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_24), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_72), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_51), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_17), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_25), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_74), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_19), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_37), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_62), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_64), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
NAND2xp33_ASAP7_75t_R g98 ( .A(n_58), .B(n_4), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_54), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_15), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_1), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_48), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_41), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_43), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_53), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_55), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_61), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_104), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_104), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_88), .B(n_0), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_106), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_119), .B(n_0), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
NAND2xp33_ASAP7_75t_R g133 ( .A(n_118), .B(n_44), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_75), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_75), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
OR2x2_ASAP7_75t_L g140 ( .A(n_94), .B(n_2), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_77), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_76), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_92), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_98), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_95), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_78), .B(n_2), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_79), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_77), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_77), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_100), .B(n_3), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_80), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_90), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_96), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_77), .Y(n_159) );
BUFx4f_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_148), .B(n_91), .Y(n_163) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_148), .B(n_100), .C(n_101), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
OAI221xp5_ASAP7_75t_L g169 ( .A1(n_132), .A2(n_105), .B1(n_111), .B2(n_101), .C(n_108), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_124), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_148), .B(n_91), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_136), .B(n_105), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_140), .B(n_108), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_137), .B(n_111), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_143), .A2(n_117), .B1(n_116), .B2(n_99), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_128), .B(n_117), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_149), .B(n_116), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
AO22x2_ASAP7_75t_L g187 ( .A1(n_149), .A2(n_99), .B1(n_83), .B2(n_86), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_147), .B(n_103), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_150), .B(n_107), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_128), .B(n_81), .C(n_83), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_157), .B(n_103), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_122), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_154), .B(n_110), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_156), .B(n_81), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_156), .B(n_86), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_122), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_122), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_139), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_120), .B(n_109), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_131), .A2(n_109), .B1(n_93), .B2(n_97), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_145), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_155), .B(n_112), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_178), .B(n_129), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
AO22x1_ASAP7_75t_L g218 ( .A1(n_178), .A2(n_82), .B1(n_102), .B2(n_155), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_170), .Y(n_219) );
OR2x2_ASAP7_75t_SL g220 ( .A(n_163), .B(n_146), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_178), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_174), .B(n_161), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_192), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_203), .Y(n_224) );
NOR2x2_ASAP7_75t_L g225 ( .A(n_180), .B(n_121), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_160), .B(n_134), .Y(n_226) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_160), .B(n_93), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_207), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_192), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_160), .B(n_97), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_184), .B(n_120), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_180), .B(n_173), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
AOI221xp5_ASAP7_75t_L g234 ( .A1(n_169), .A2(n_125), .B1(n_142), .B2(n_151), .C(n_112), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_184), .B(n_212), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_203), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_204), .Y(n_238) );
NAND3xp33_ASAP7_75t_SL g239 ( .A(n_172), .B(n_125), .C(n_151), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_186), .Y(n_242) );
BUFx2_ASAP7_75t_SL g243 ( .A(n_197), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_184), .B(n_142), .Y(n_245) );
INVx6_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_184), .B(n_151), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_212), .B(n_190), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_180), .B(n_133), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_211), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_212), .B(n_159), .Y(n_255) );
NOR3xp33_ASAP7_75t_SL g256 ( .A(n_172), .B(n_3), .C(n_4), .Y(n_256) );
NOR3xp33_ASAP7_75t_SL g257 ( .A(n_189), .B(n_5), .C(n_6), .Y(n_257) );
NOR3xp33_ASAP7_75t_SL g258 ( .A(n_164), .B(n_5), .C(n_7), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_193), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_181), .B(n_7), .Y(n_261) );
BUFx12f_ASAP7_75t_SL g262 ( .A(n_176), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_175), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_205), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_176), .B(n_123), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_181), .B(n_9), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_168), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_198), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_228), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_228), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
OR2x6_ASAP7_75t_L g273 ( .A(n_253), .B(n_187), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_222), .B(n_165), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_232), .A2(n_187), .B1(n_182), .B2(n_191), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_269), .B(n_188), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_213), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_250), .A2(n_183), .B(n_196), .Y(n_278) );
CKINVDCx8_ASAP7_75t_R g279 ( .A(n_243), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_253), .B(n_177), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_214), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_253), .B(n_194), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_219), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_236), .A2(n_210), .B1(n_200), .B2(n_179), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_215), .B(n_209), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_244), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_253), .B(n_171), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_231), .A2(n_185), .B(n_199), .Y(n_291) );
AO21x1_ASAP7_75t_L g292 ( .A1(n_261), .A2(n_159), .B(n_152), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_232), .B(n_199), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_213), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_261), .B(n_187), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_221), .B(n_187), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_261), .A2(n_182), .B1(n_185), .B2(n_206), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_223), .B(n_159), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_223), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_259), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_223), .Y(n_307) );
NOR2xp33_ASAP7_75t_SL g308 ( .A(n_262), .B(n_182), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_254), .Y(n_309) );
BUFx10_ASAP7_75t_L g310 ( .A(n_247), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_217), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_217), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_223), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_243), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_246), .A2(n_182), .B1(n_152), .B2(n_153), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_283), .B(n_267), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_283), .B(n_267), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_283), .A2(n_252), .B1(n_227), .B2(n_267), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_296), .B(n_267), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
BUFx10_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_303), .A2(n_252), .B1(n_227), .B2(n_245), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_286), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_288), .A2(n_252), .B1(n_227), .B2(n_246), .Y(n_324) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_314), .B(n_256), .C(n_257), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_308), .B(n_229), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_252), .B1(n_246), .B2(n_249), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_293), .A2(n_252), .B1(n_246), .B2(n_239), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_278), .A2(n_264), .B(n_268), .C(n_260), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_229), .B1(n_216), .B2(n_234), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_273), .A2(n_268), .B1(n_258), .B2(n_237), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_224), .B1(n_217), .B2(n_237), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_276), .B(n_218), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_287), .A2(n_218), .B1(n_226), .B2(n_230), .C(n_255), .Y(n_336) );
OAI222xp33_ASAP7_75t_L g337 ( .A1(n_273), .A2(n_225), .B1(n_220), .B2(n_260), .C1(n_233), .C2(n_235), .Y(n_337) );
NAND2xp33_ASAP7_75t_SL g338 ( .A(n_296), .B(n_229), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_273), .A2(n_229), .B1(n_224), .B2(n_237), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_275), .A2(n_229), .B1(n_224), .B2(n_238), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_293), .A2(n_233), .B1(n_235), .B2(n_248), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_279), .A2(n_238), .B1(n_265), .B2(n_263), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g344 ( .A(n_284), .B(n_242), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_322), .A2(n_282), .B1(n_293), .B2(n_306), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_318), .A2(n_299), .B1(n_271), .B2(n_289), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_343), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_333), .B(n_315), .C(n_297), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_340), .A2(n_292), .B(n_304), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_326), .B(n_271), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_331), .A2(n_291), .B(n_289), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_322), .A2(n_299), .B1(n_298), .B2(n_309), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_319), .B(n_274), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_321), .A2(n_282), .B1(n_309), .B2(n_298), .Y(n_354) );
OA21x2_ASAP7_75t_L g355 ( .A1(n_334), .A2(n_292), .B(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_333), .B(n_284), .C(n_294), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_282), .B1(n_290), .B2(n_302), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_319), .B(n_311), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_337), .B(n_220), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_324), .A2(n_290), .B1(n_280), .B2(n_301), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_334), .A2(n_279), .B1(n_311), .B2(n_312), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_285), .B(n_312), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_316), .B(n_281), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
AOI21x1_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_152), .B(n_153), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_290), .B1(n_301), .B2(n_235), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_316), .A2(n_285), .B1(n_300), .B2(n_290), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_317), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_364), .Y(n_371) );
NOR4xp25_ASAP7_75t_SL g372 ( .A(n_356), .B(n_338), .C(n_336), .D(n_321), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_353), .B(n_323), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_362), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_347), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_356), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_360), .A2(n_328), .B1(n_332), .B2(n_330), .C(n_317), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_365), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_365), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_364), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_339), .B1(n_341), .B2(n_342), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_353), .B(n_321), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_368), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_368), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_370), .B(n_321), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_349), .A2(n_320), .B(n_304), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_346), .A2(n_320), .B1(n_300), .B2(n_277), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_320), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_359), .B(n_301), .Y(n_391) );
OAI33xp33_ASAP7_75t_L g392 ( .A1(n_346), .A2(n_153), .A3(n_266), .B1(n_251), .B2(n_12), .B3(n_13), .Y(n_392) );
NAND2xp33_ASAP7_75t_R g393 ( .A(n_355), .B(n_295), .Y(n_393) );
OAI31xp33_ASAP7_75t_SL g394 ( .A1(n_352), .A2(n_251), .A3(n_238), .B(n_310), .Y(n_394) );
NAND2xp33_ASAP7_75t_R g395 ( .A(n_355), .B(n_295), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_233), .B1(n_248), .B2(n_235), .C(n_251), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_370), .A2(n_358), .B1(n_354), .B2(n_359), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_350), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_357), .B(n_277), .C(n_344), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g401 ( .A(n_357), .B(n_277), .Y(n_401) );
OAI33xp33_ASAP7_75t_L g402 ( .A1(n_348), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_380), .B(n_355), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_394), .B(n_351), .C(n_367), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_390), .B(n_348), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_390), .B(n_351), .Y(n_412) );
OAI33xp33_ASAP7_75t_L g413 ( .A1(n_373), .A2(n_11), .A3(n_14), .B1(n_16), .B2(n_18), .B3(n_19), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_391), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_398), .B(n_369), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_378), .B(n_355), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_379), .B(n_363), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_379), .B(n_363), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_374), .B(n_349), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_402), .A2(n_361), .B1(n_369), .B2(n_248), .C(n_233), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_399), .B(n_272), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_391), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_385), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_386), .B(n_14), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_392), .A2(n_248), .B1(n_123), .B2(n_122), .C(n_141), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_384), .B(n_310), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_388), .B(n_366), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
NAND2xp67_ASAP7_75t_L g440 ( .A(n_372), .B(n_18), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g442 ( .A1(n_397), .A2(n_304), .A3(n_272), .B(n_307), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_387), .B(n_20), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_377), .B(n_284), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_382), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_393), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_395), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_396), .B(n_284), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_404), .B(n_20), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_418), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_414), .B(n_21), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_443), .B(n_123), .C(n_122), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_420), .B(n_366), .Y(n_453) );
CKINVDCx8_ASAP7_75t_R g454 ( .A(n_418), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_445), .A2(n_123), .B(n_141), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_438), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_425), .B(n_21), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_443), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_123), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_413), .B(n_313), .C(n_305), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_433), .B(n_22), .Y(n_465) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_446), .B(n_294), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_433), .B(n_22), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_436), .B(n_23), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_428), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_445), .B(n_23), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_436), .B(n_277), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_435), .Y(n_473) );
AOI21xp5_ASAP7_75t_SL g474 ( .A1(n_428), .A2(n_284), .B(n_294), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_277), .Y(n_475) );
NOR3xp33_ASAP7_75t_SL g476 ( .A(n_407), .B(n_26), .C(n_28), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_409), .B(n_123), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_430), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_403), .Y(n_479) );
NAND5xp2_ASAP7_75t_L g480 ( .A(n_442), .B(n_310), .C(n_30), .D(n_33), .E(n_34), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_405), .B(n_307), .C(n_313), .D(n_305), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_410), .B(n_141), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_405), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_410), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_446), .B(n_294), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_411), .B(n_294), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_411), .B(n_313), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_423), .B(n_122), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_430), .Y(n_489) );
OAI21x1_ASAP7_75t_SL g490 ( .A1(n_424), .A2(n_29), .B(n_38), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_423), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_427), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_427), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_416), .B(n_305), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_417), .B(n_295), .Y(n_495) );
INVx5_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
NAND2xp33_ASAP7_75t_R g497 ( .A(n_435), .B(n_39), .Y(n_497) );
NOR3xp33_ASAP7_75t_SL g498 ( .A(n_434), .B(n_49), .C(n_50), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_415), .B(n_141), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_417), .B(n_141), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_432), .B(n_52), .C(n_56), .D(n_57), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_474), .B(n_424), .C(n_422), .D(n_447), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_480), .A2(n_447), .A3(n_441), .B(n_444), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_456), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_458), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_474), .A2(n_437), .B(n_441), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_491), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_469), .B(n_419), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_470), .A2(n_412), .B1(n_420), .B2(n_444), .C1(n_419), .C2(n_439), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_458), .B(n_406), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_457), .B(n_406), .Y(n_511) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_481), .B(n_431), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_473), .B(n_420), .C(n_431), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_452), .A2(n_448), .B(n_437), .Y(n_514) );
NAND2xp33_ASAP7_75t_SL g515 ( .A(n_497), .B(n_412), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_459), .B(n_412), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_471), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_451), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_492), .Y(n_519) );
AOI322xp5_ASAP7_75t_L g520 ( .A1(n_461), .A2(n_412), .A3(n_420), .B1(n_439), .B2(n_448), .C1(n_431), .C2(n_437), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_479), .B(n_408), .Y(n_521) );
AOI21xp33_ASAP7_75t_SL g522 ( .A1(n_497), .A2(n_408), .B(n_431), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_494), .B(n_408), .Y(n_523) );
AOI21xp33_ASAP7_75t_SL g524 ( .A1(n_466), .A2(n_408), .B(n_440), .Y(n_524) );
AND3x2_ASAP7_75t_L g525 ( .A(n_450), .B(n_440), .C(n_408), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_454), .A2(n_476), .B1(n_498), .B2(n_466), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_483), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_478), .B(n_141), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_454), .A2(n_242), .B1(n_241), .B2(n_240), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_496), .B(n_59), .Y(n_530) );
NOR4xp25_ASAP7_75t_L g531 ( .A(n_449), .B(n_265), .C(n_263), .D(n_69), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
AOI32xp33_ASAP7_75t_L g533 ( .A1(n_460), .A2(n_240), .A3(n_60), .B1(n_63), .B2(n_265), .Y(n_533) );
OAI22xp33_ASAP7_75t_SL g534 ( .A1(n_467), .A2(n_240), .B1(n_263), .B2(n_242), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_489), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_495), .A2(n_242), .B1(n_241), .B2(n_201), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_465), .A2(n_242), .B(n_241), .C(n_202), .Y(n_537) );
NOR4xp25_ASAP7_75t_SL g538 ( .A(n_450), .B(n_166), .C(n_202), .D(n_201), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_468), .B(n_166), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_473), .B(n_166), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_462), .B(n_241), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_500), .A2(n_166), .B1(n_202), .B2(n_201), .C(n_195), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_462), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_464), .Y(n_545) );
NOR2xp33_ASAP7_75t_SL g546 ( .A(n_490), .B(n_241), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_493), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_476), .A2(n_241), .B(n_202), .C(n_166), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_487), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_541), .Y(n_551) );
AND4x1_ASAP7_75t_L g552 ( .A(n_546), .B(n_498), .C(n_463), .D(n_475), .Y(n_552) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_518), .A2(n_499), .B(n_485), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_523), .B(n_496), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_508), .B(n_484), .Y(n_556) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_522), .A2(n_463), .B(n_455), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_517), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_547), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_505), .B(n_484), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_507), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_510), .B(n_486), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_532), .Y(n_565) );
OAI21xp33_ASAP7_75t_L g566 ( .A1(n_520), .A2(n_485), .B(n_501), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_545), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_535), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_512), .A2(n_485), .B(n_472), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_549), .B(n_496), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_511), .Y(n_572) );
NOR2xp67_ASAP7_75t_SL g573 ( .A(n_506), .B(n_496), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_515), .A2(n_453), .B(n_482), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_509), .B(n_477), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_521), .B(n_488), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_503), .B(n_453), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_514), .B(n_453), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_526), .B(n_202), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_581), .B(n_502), .C(n_524), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_554), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_576), .A2(n_539), .B1(n_513), .B2(n_525), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_558), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_560), .Y(n_587) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_570), .A2(n_533), .B(n_531), .C(n_548), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
XNOR2xp5_ASAP7_75t_L g591 ( .A(n_552), .B(n_525), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_557), .A2(n_548), .B(n_534), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_578), .B(n_540), .C(n_537), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_566), .A2(n_537), .B(n_530), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g595 ( .A1(n_559), .A2(n_529), .B(n_539), .C(n_540), .Y(n_595) );
XNOR2x2_ASAP7_75t_L g596 ( .A(n_574), .B(n_542), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_563), .A2(n_529), .B(n_543), .C(n_538), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_556), .Y(n_598) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_580), .A2(n_536), .B1(n_195), .B2(n_201), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_573), .B(n_195), .C(n_568), .Y(n_600) );
NOR2xp33_ASAP7_75t_R g601 ( .A(n_591), .B(n_580), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_591), .A2(n_579), .B1(n_572), .B2(n_569), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_584), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_598), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_592), .A2(n_579), .B1(n_575), .B2(n_573), .C1(n_565), .C2(n_550), .Y(n_605) );
NOR2x1_ASAP7_75t_R g606 ( .A(n_596), .B(n_580), .Y(n_606) );
NAND2xp33_ASAP7_75t_SL g607 ( .A(n_585), .B(n_555), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_596), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_588), .B(n_553), .C(n_582), .Y(n_609) );
XOR2x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_571), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_594), .A2(n_597), .B(n_593), .C(n_600), .Y(n_611) );
AO22x1_ASAP7_75t_L g612 ( .A1(n_590), .A2(n_561), .B1(n_562), .B2(n_551), .Y(n_612) );
AND4x1_ASAP7_75t_L g613 ( .A(n_585), .B(n_595), .C(n_599), .D(n_586), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_590), .A2(n_564), .B1(n_577), .B2(n_567), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_587), .A2(n_577), .B1(n_551), .B2(n_567), .C(n_195), .Y(n_615) );
OAI311xp33_ASAP7_75t_L g616 ( .A1(n_589), .A2(n_585), .A3(n_592), .B1(n_566), .C1(n_593), .Y(n_616) );
OAI21x1_ASAP7_75t_SL g617 ( .A1(n_611), .A2(n_602), .B(n_606), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_604), .Y(n_618) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_608), .B(n_611), .C(n_613), .Y(n_619) );
NAND4xp25_ASAP7_75t_SL g620 ( .A(n_605), .B(n_609), .C(n_616), .D(n_601), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g621 ( .A(n_620), .B(n_603), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_618), .B(n_607), .Y(n_622) );
OAI222xp33_ASAP7_75t_L g623 ( .A1(n_617), .A2(n_607), .B1(n_615), .B2(n_610), .C1(n_614), .C2(n_601), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_622), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_621), .Y(n_625) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_625), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_626), .A2(n_619), .B1(n_624), .B2(n_623), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_627), .A2(n_624), .B(n_612), .Y(n_628) );
endmodule