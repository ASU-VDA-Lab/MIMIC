module fake_ariane_2303_n_106 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_106);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_106;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_81;
wire n_87;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

BUFx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_R g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_R g46 ( 
.A(n_31),
.B(n_12),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_29),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_27),
.B(n_26),
.C(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_45),
.B1(n_42),
.B2(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_47),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_39),
.B(n_44),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_44),
.B(n_33),
.C(n_30),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_55),
.B(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_50),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_48),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_65),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_62),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_73),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_35),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_77),
.Y(n_82)
);

OR2x6_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_69),
.B(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_91),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_86),
.B(n_51),
.C(n_43),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_51),
.B1(n_43),
.B2(n_46),
.C(n_41),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_41),
.B1(n_23),
.B2(n_55),
.C(n_6),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_95),
.B(n_92),
.C(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.C(n_98),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI211xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_23),
.B(n_3),
.C(n_5),
.Y(n_104)
);

AOI222xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.C1(n_2),
.C2(n_83),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_23),
.B1(n_7),
.B2(n_2),
.C(n_13),
.Y(n_106)
);


endmodule