module fake_jpeg_535_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_30),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_75),
.Y(n_95)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_60),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_68),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_1),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_66),
.Y(n_92)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_16),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_76),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_28),
.Y(n_88)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_12),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_36),
.B1(n_40),
.B2(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_91),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_36),
.B1(n_38),
.B2(n_29),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_97),
.B1(n_113),
.B2(n_69),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_100),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_40),
.B1(n_43),
.B2(n_38),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_27),
.CON(n_98),
.SN(n_98)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_43),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_32),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_26),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_124),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_34),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_4),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_5),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_128),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_44),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_144),
.C(n_149),
.Y(n_176)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_143),
.Y(n_161)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_141),
.C(n_147),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_79),
.A2(n_64),
.B1(n_74),
.B2(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_5),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_22),
.B1(n_34),
.B2(n_80),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_98),
.A2(n_34),
.B(n_97),
.C(n_112),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_34),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_101),
.Y(n_165)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_119),
.B(n_87),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_128),
.B(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_92),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_105),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_146),
.C(n_114),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_122),
.B1(n_96),
.B2(n_86),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_156),
.B1(n_152),
.B2(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_85),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_83),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_177),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_93),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_102),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_102),
.B1(n_96),
.B2(n_123),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_128),
.B1(n_154),
.B2(n_142),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_132),
.B(n_149),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_114),
.A3(n_81),
.B1(n_115),
.B2(n_118),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_123),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_196),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_192),
.B1(n_197),
.B2(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_195),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_145),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_194),
.B(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_176),
.C(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_118),
.B1(n_133),
.B2(n_81),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_137),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_82),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_195),
.C(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_160),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_159),
.B(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_191),
.B(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_209),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_188),
.B(n_202),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_211),
.C(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_212),
.A2(n_170),
.B1(n_205),
.B2(n_159),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_232),
.B1(n_223),
.B2(n_225),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_170),
.B(n_191),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_198),
.B1(n_199),
.B2(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_240),
.B(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_207),
.C(n_213),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_222),
.B1(n_221),
.B2(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_226),
.B1(n_236),
.B2(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_190),
.C(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_250),
.B1(n_247),
.B2(n_246),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_236),
.B1(n_230),
.B2(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_254),
.B(n_246),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_229),
.B(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_251),
.C(n_248),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_249),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_250),
.A2(n_228),
.B1(n_235),
.B2(n_242),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

NAND4xp25_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.C(n_187),
.D(n_180),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.C(n_162),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_217),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_220),
.B(n_210),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_269),
.B(n_267),
.C(n_161),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_266),
.A2(n_206),
.B1(n_178),
.B2(n_167),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_262),
.C(n_197),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_272),
.A3(n_161),
.B1(n_178),
.B2(n_183),
.C1(n_169),
.C2(n_175),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_270),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_274),
.B(n_175),
.C(n_82),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_106),
.Y(n_276)
);


endmodule