module fake_jpeg_16223_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_62),
.B1(n_41),
.B2(n_54),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_56),
.B(n_2),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_61),
.B1(n_44),
.B2(n_49),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_92),
.B(n_94),
.C(n_108),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_45),
.B1(n_52),
.B2(n_50),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_5),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_56),
.B1(n_48),
.B2(n_60),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_58),
.B1(n_53),
.B2(n_57),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_16),
.B1(n_36),
.B2(n_35),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_113),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_124),
.B(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_106),
.Y(n_133)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_105),
.B(n_97),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_119),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_130),
.B1(n_122),
.B2(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_140),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_116),
.B(n_101),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_116),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_144),
.C(n_137),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_151),
.B1(n_117),
.B2(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_7),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_103),
.B(n_104),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_22),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_20),
.C(n_8),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_24),
.C(n_10),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_31),
.B(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_32),
.B(n_12),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_111),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule