module fake_netlist_5_1005_n_919 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_919);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_919;

wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_443;
wire n_372;
wire n_293;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_449;
wire n_325;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_894;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_338;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_846;
wire n_586;
wire n_748;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_217;
wire n_440;
wire n_793;
wire n_478;
wire n_726;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_237;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_491;
wire n_272;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_8),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_7),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_42),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_161),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_31),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_73),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_97),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_124),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_22),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_68),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_70),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_85),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_57),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_191),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_60),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_41),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_166),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_64),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_162),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_66),
.B(n_198),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_190),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_74),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_87),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_89),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_63),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_133),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_86),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_20),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_193),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_48),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_33),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_128),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_91),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_131),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_179),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_117),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_37),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_81),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_1),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_201),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_126),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_78),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_98),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_160),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_92),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_93),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_62),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_50),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_157),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_16),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_111),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_199),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_65),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_11),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_156),
.B(n_186),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_110),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_25),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_167),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_56),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_205),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_187),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_100),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_189),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_132),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_90),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_144),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_135),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_134),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_47),
.B(n_178),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_125),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_113),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_88),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_171),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_202),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_195),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_159),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_83),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_137),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_53),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_183),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_103),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_149),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_17),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_109),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_43),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_143),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_19),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_145),
.B(n_23),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_44),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_123),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_152),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_174),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_112),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_54),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_79),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_163),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_172),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_3),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_138),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_27),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_11),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_95),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_36),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_94),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_177),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_4),
.Y(n_362)
);

BUFx2_ASAP7_75t_SL g363 ( 
.A(n_168),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_67),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_216),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_210),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_0),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_212),
.B(n_0),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_214),
.B(n_1),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_288),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_216),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_342),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_232),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_257),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_216),
.B(n_28),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_244),
.A2(n_104),
.B(n_206),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_240),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_250),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_265),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_222),
.B(n_2),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_250),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_234),
.B(n_29),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_268),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_250),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_327),
.B(n_2),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_235),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_266),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_240),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_265),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

OAI22x1_ASAP7_75t_SL g398 ( 
.A1(n_299),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_240),
.Y(n_399)
);

AOI22x1_ASAP7_75t_SL g400 ( 
.A1(n_306),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_281),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_266),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_242),
.B(n_6),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_309),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_217),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_9),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_362),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_290),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_218),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_208),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_290),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_223),
.B(n_10),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_290),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_295),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_233),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_224),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_295),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_258),
.B(n_12),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_225),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_295),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_230),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_326),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_311),
.B(n_12),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_259),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_231),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_209),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_211),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_241),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_247),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_251),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_13),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_271),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_312),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_253),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_213),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_256),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_314),
.B(n_14),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_317),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_349),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_261),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_336),
.B(n_15),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_263),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_360),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_343),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_215),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_264),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_269),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_275),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_270),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_276),
.B(n_21),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_277),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_278),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_367),
.B(n_323),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_379),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_369),
.B(n_239),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_425),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

NOR2x1p5_ASAP7_75t_L g477 ( 
.A(n_403),
.B(n_219),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_416),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_280),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_425),
.B(n_308),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

BUFx6f_ASAP7_75t_SL g487 ( 
.A(n_396),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_375),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g501 ( 
.A(n_376),
.B(n_363),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_368),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_449),
.B(n_254),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_420),
.Y(n_511)
);

AND2x2_ASAP7_75t_SL g512 ( 
.A(n_431),
.B(n_307),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_372),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_401),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_373),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_427),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_461),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_447),
.B(n_283),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_220),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

AO21x2_ASAP7_75t_L g527 ( 
.A1(n_430),
.A2(n_453),
.B(n_392),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_413),
.B(n_284),
.Y(n_528)
);

AO22x2_ASAP7_75t_L g529 ( 
.A1(n_456),
.A2(n_364),
.B1(n_361),
.B2(n_359),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_449),
.B(n_273),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_386),
.B(n_334),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_436),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_378),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_286),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_378),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_374),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_374),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_383),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_370),
.B(n_282),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_287),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_417),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_387),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_514),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_512),
.A2(n_451),
.B1(n_421),
.B2(n_462),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_500),
.B(n_541),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_417),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_533),
.B(n_408),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_472),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_433),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_433),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_475),
.B(n_433),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_537),
.B(n_380),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_475),
.B(n_381),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_512),
.A2(n_304),
.B1(n_310),
.B2(n_285),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_475),
.B(n_455),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_426),
.C(n_422),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_467),
.B(n_479),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

NOR2x1p5_ASAP7_75t_L g566 ( 
.A(n_500),
.B(n_385),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_475),
.B(n_455),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_475),
.B(n_455),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_481),
.B(n_524),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_479),
.B(n_412),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_479),
.B(n_377),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_469),
.B(n_370),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_530),
.A2(n_348),
.B1(n_355),
.B2(n_347),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_469),
.B(n_460),
.Y(n_575)
);

O2A1O1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_483),
.A2(n_458),
.B(n_459),
.C(n_432),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_480),
.B(n_376),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_465),
.B(n_395),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_466),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_483),
.B(n_434),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_490),
.B(n_406),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_406),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_484),
.B(n_444),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_530),
.B(n_411),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_490),
.B(n_411),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_484),
.B(n_444),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_490),
.B(n_434),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_441),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_529),
.A2(n_356),
.B1(n_390),
.B2(n_402),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_482),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_529),
.A2(n_410),
.B1(n_428),
.B2(n_415),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_488),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_501),
.B(n_221),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_488),
.B(n_444),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_L g600 ( 
.A1(n_529),
.A2(n_398),
.B1(n_402),
.B2(n_410),
.C(n_415),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_489),
.B(n_445),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_489),
.B(n_445),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_534),
.B(n_442),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_521),
.B(n_226),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_542),
.B(n_446),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_487),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_466),
.B(n_227),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_445),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_538),
.B(n_393),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_487),
.B(n_400),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_477),
.A2(n_319),
.B1(n_229),
.B2(n_236),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_294),
.C(n_293),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_513),
.A2(n_428),
.B(n_440),
.C(n_382),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_525),
.B(n_404),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_471),
.B(n_440),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_450),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_544),
.A2(n_389),
.B(n_492),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_548),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_543),
.A2(n_494),
.B(n_493),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_583),
.B(n_450),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_585),
.B(n_494),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_584),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_589),
.B(n_496),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_558),
.A2(n_498),
.B(n_496),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_603),
.B(n_498),
.Y(n_625)
);

OAI21xp33_ASAP7_75t_SL g626 ( 
.A1(n_573),
.A2(n_298),
.B(n_297),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_554),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_588),
.B(n_228),
.Y(n_628)
);

AO21x1_ASAP7_75t_L g629 ( 
.A1(n_546),
.A2(n_305),
.B(n_303),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_555),
.B(n_502),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_502),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_606),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_561),
.B(n_237),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_564),
.A2(n_546),
.B1(n_614),
.B2(n_586),
.Y(n_634)
);

AO21x1_ASAP7_75t_L g635 ( 
.A1(n_591),
.A2(n_316),
.B(n_315),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_581),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_576),
.A2(n_452),
.B(n_454),
.C(n_448),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_552),
.B(n_504),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_614),
.B(n_516),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_553),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_582),
.B(n_609),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_329),
.B(n_324),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_556),
.A2(n_335),
.B(n_332),
.Y(n_644)
);

AND2x6_ASAP7_75t_SL g645 ( 
.A(n_547),
.B(n_400),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_560),
.A2(n_346),
.B(n_339),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g647 ( 
.A1(n_595),
.A2(n_351),
.A3(n_358),
.B1(n_495),
.B2(n_476),
.C(n_465),
.Y(n_647)
);

BUFx2_ASAP7_75t_SL g648 ( 
.A(n_545),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_587),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_611),
.B(n_238),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_567),
.A2(n_507),
.B(n_505),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_568),
.A2(n_508),
.B(n_507),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

AO21x1_ASAP7_75t_L g654 ( 
.A1(n_591),
.A2(n_407),
.B(n_399),
.Y(n_654)
);

BUFx4f_ASAP7_75t_L g655 ( 
.A(n_606),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_557),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_549),
.B(n_562),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_565),
.B(n_570),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_563),
.A2(n_464),
.B(n_454),
.C(n_452),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_578),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_577),
.A2(n_509),
.B(n_508),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_559),
.A2(n_325),
.B1(n_245),
.B2(n_246),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_599),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_563),
.A2(n_338),
.B1(n_248),
.B2(n_249),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_572),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_579),
.A2(n_511),
.B(n_509),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_547),
.A2(n_340),
.B1(n_252),
.B2(n_255),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_601),
.A2(n_608),
.B(n_602),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_448),
.B(n_464),
.C(n_539),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_598),
.A2(n_381),
.B(n_515),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_590),
.B(n_517),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_592),
.B(n_517),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_593),
.A2(n_519),
.B(n_518),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_571),
.B(n_243),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_518),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_550),
.B(n_260),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_580),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_547),
.B(n_404),
.Y(n_679)
);

OAI21xp33_ASAP7_75t_L g680 ( 
.A1(n_641),
.A2(n_594),
.B(n_600),
.Y(n_680)
);

AO21x1_ASAP7_75t_L g681 ( 
.A1(n_642),
.A2(n_597),
.B(n_612),
.Y(n_681)
);

AOI21x1_ASAP7_75t_SL g682 ( 
.A1(n_627),
.A2(n_630),
.B(n_657),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

AO31x2_ASAP7_75t_L g684 ( 
.A1(n_654),
.A2(n_526),
.A3(n_520),
.B(n_535),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_634),
.A2(n_607),
.B(n_262),
.C(n_328),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_643),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_678),
.Y(n_687)
);

AOI221x1_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_463),
.B1(n_532),
.B2(n_522),
.C(n_523),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_624),
.A2(n_526),
.B(n_520),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_616),
.B(n_580),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_622),
.B(n_470),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_648),
.B(n_566),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_668),
.A2(n_536),
.B(n_470),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_619),
.A2(n_539),
.B(n_499),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_618),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_651),
.A2(n_499),
.B(n_497),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_649),
.B(n_267),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_665),
.A2(n_322),
.B(n_274),
.C(n_279),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_663),
.B(n_272),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_652),
.A2(n_506),
.B(n_497),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_631),
.B(n_289),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_617),
.A2(n_381),
.B(n_292),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_621),
.A2(n_296),
.B(n_291),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_625),
.B(n_620),
.Y(n_704)
);

AO21x2_ASAP7_75t_L g705 ( 
.A1(n_646),
.A2(n_381),
.B(n_32),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_679),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_610),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_679),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_661),
.A2(n_140),
.B(n_207),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_623),
.A2(n_321),
.B(n_353),
.Y(n_710)
);

AO21x2_ASAP7_75t_L g711 ( 
.A1(n_670),
.A2(n_344),
.B(n_352),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_674),
.A2(n_320),
.B(n_301),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_653),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_633),
.B(n_300),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_666),
.A2(n_130),
.B(n_203),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_647),
.A2(n_318),
.B(n_350),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_678),
.B(n_640),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_658),
.A2(n_129),
.B(n_194),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_638),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_463),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_660),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_721),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_704),
.A2(n_650),
.B(n_626),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_719),
.A2(n_669),
.B(n_672),
.Y(n_725)
);

NOR2x1_ASAP7_75t_R g726 ( 
.A(n_706),
.B(n_632),
.Y(n_726)
);

AO21x2_ASAP7_75t_L g727 ( 
.A1(n_681),
.A2(n_629),
.B(n_675),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_713),
.Y(n_728)
);

OA21x2_ASAP7_75t_L g729 ( 
.A1(n_688),
.A2(n_671),
.B(n_673),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_693),
.A2(n_637),
.B(n_659),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_687),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_719),
.B(n_635),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_687),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_702),
.A2(n_628),
.B(n_662),
.Y(n_734)
);

AO21x2_ASAP7_75t_L g735 ( 
.A1(n_711),
.A2(n_676),
.B(n_667),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_717),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_692),
.B(n_639),
.Y(n_737)
);

INVx6_ASAP7_75t_L g738 ( 
.A(n_713),
.Y(n_738)
);

OA21x2_ASAP7_75t_L g739 ( 
.A1(n_694),
.A2(n_664),
.B(n_639),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_686),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_709),
.A2(n_677),
.B(n_653),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_680),
.B(n_701),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_706),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_691),
.Y(n_745)
);

BUFx2_ASAP7_75t_SL g746 ( 
.A(n_683),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_711),
.A2(n_677),
.B(n_463),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_689),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_715),
.A2(n_677),
.B(n_121),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_720),
.B(n_655),
.Y(n_750)
);

OAI21x1_ASAP7_75t_L g751 ( 
.A1(n_682),
.A2(n_119),
.B(n_182),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_743),
.A2(n_714),
.B(n_710),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_732),
.A2(n_712),
.B1(n_734),
.B2(n_745),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_723),
.A2(n_697),
.B(n_699),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_738),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_731),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_732),
.B(n_695),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_731),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_733),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_733),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_738),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_722),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_724),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_736),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_736),
.B(n_684),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_750),
.A2(n_716),
.B1(n_707),
.B2(n_708),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_729),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_742),
.A2(n_700),
.B(n_696),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_750),
.B(n_684),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_727),
.B(n_684),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_729),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_725),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_746),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_744),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_746),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_741),
.Y(n_778)
);

AND2x4_ASAP7_75t_SL g779 ( 
.A(n_761),
.B(n_728),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_758),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_766),
.A2(n_735),
.B1(n_727),
.B2(n_705),
.Y(n_781)
);

CKINVDCx6p67_ASAP7_75t_R g782 ( 
.A(n_775),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_757),
.B(n_735),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_757),
.B(n_737),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_769),
.B(n_735),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_762),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_769),
.B(n_772),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_778),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_778),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_761),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_764),
.B(n_747),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_753),
.B(n_765),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_756),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_762),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_759),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_775),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_765),
.B(n_747),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_763),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_752),
.B(n_645),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_759),
.B(n_747),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_760),
.B(n_685),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_760),
.B(n_751),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_772),
.B(n_690),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_767),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_787),
.B(n_770),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_787),
.B(n_770),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_786),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_800),
.B(n_774),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_795),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_793),
.B(n_773),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_799),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_783),
.B(n_773),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_788),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_794),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_794),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_781),
.A2(n_754),
.B(n_698),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_796),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_791),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_791),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_784),
.B(n_789),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_784),
.B(n_777),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_784),
.B(n_761),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_780),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_783),
.B(n_767),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_790),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_790),
.B(n_755),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_793),
.B(n_780),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_805),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_785),
.B(n_771),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_792),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_792),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_831),
.B(n_798),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_807),
.B(n_798),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_832),
.B(n_801),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_821),
.Y(n_836)
);

AND2x4_ASAP7_75t_SL g837 ( 
.A(n_827),
.B(n_782),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_828),
.B(n_802),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_808),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_810),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_817),
.B(n_802),
.C(n_703),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_812),
.B(n_803),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_830),
.B(n_804),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_825),
.B(n_803),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_806),
.B(n_771),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_806),
.B(n_813),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_811),
.B(n_776),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_814),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_811),
.B(n_776),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_815),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_815),
.B(n_804),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_809),
.B(n_826),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_836),
.B(n_823),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_839),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_840),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_848),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_842),
.B(n_816),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_848),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_837),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_846),
.B(n_822),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_842),
.B(n_829),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_852),
.Y(n_862)
);

NOR2x1p5_ASAP7_75t_SL g863 ( 
.A(n_850),
.B(n_818),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_854),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_862),
.A2(n_841),
.B1(n_838),
.B2(n_834),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_860),
.B(n_843),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_855),
.Y(n_867)
);

NAND4xp75_ASAP7_75t_SL g868 ( 
.A(n_853),
.B(n_851),
.C(n_845),
.D(n_849),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_859),
.A2(n_833),
.B1(n_844),
.B2(n_797),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_865),
.B(n_857),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_864),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_867),
.Y(n_872)
);

OAI222xp33_ASAP7_75t_L g873 ( 
.A1(n_869),
.A2(n_861),
.B1(n_835),
.B2(n_858),
.C1(n_856),
.C2(n_850),
.Y(n_873)
);

OAI31xp33_ASAP7_75t_L g874 ( 
.A1(n_866),
.A2(n_849),
.A3(n_847),
.B(n_820),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_868),
.A2(n_726),
.B(n_819),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_865),
.A2(n_819),
.B(n_824),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_864),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_874),
.B(n_863),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_SL g879 ( 
.A(n_873),
.B(n_744),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_870),
.B(n_706),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_875),
.A2(n_718),
.B(n_749),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_779),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_871),
.B(n_779),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_877),
.B(n_739),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_871),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_SL g886 ( 
.A1(n_876),
.A2(n_683),
.B(n_49),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_882),
.B(n_749),
.Y(n_887)
);

NOR2x1_ASAP7_75t_L g888 ( 
.A(n_880),
.B(n_740),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_885),
.Y(n_889)
);

NAND5xp2_ASAP7_75t_L g890 ( 
.A(n_886),
.B(n_51),
.C(n_55),
.D(n_58),
.E(n_59),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_883),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_879),
.B(n_748),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_878),
.A2(n_739),
.B(n_730),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_889),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_888),
.B(n_884),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_893),
.B(n_881),
.Y(n_896)
);

NAND4xp25_ASAP7_75t_L g897 ( 
.A(n_890),
.B(n_75),
.C(n_76),
.D(n_77),
.Y(n_897)
);

NOR3x1_ASAP7_75t_L g898 ( 
.A(n_892),
.B(n_768),
.C(n_82),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_887),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_891),
.B(n_80),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_894),
.Y(n_901)
);

NOR3x1_ASAP7_75t_L g902 ( 
.A(n_900),
.B(n_897),
.C(n_896),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_898),
.B(n_895),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_899),
.B(n_84),
.Y(n_904)
);

AOI31xp33_ASAP7_75t_L g905 ( 
.A1(n_903),
.A2(n_102),
.A3(n_107),
.B(n_114),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_902),
.B(n_115),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_901),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_904),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_908),
.B(n_116),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_906),
.B(n_907),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_905),
.B(n_118),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_910),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_912),
.B(n_909),
.C(n_911),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_913),
.B(n_146),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_915),
.B(n_158),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_916),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_917),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_918),
.A2(n_169),
.B(n_170),
.Y(n_919)
);


endmodule