module fake_ariane_409_n_887 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_887);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_887;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_818;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_838;
wire n_623;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_278;
wire n_609;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_856;
wire n_782;
wire n_650;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_68),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_78),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_66),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_14),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_27),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_84),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_92),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_150),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_130),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_80),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_79),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_166),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_127),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_82),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_2),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_112),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_99),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_107),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_44),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_39),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_151),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_74),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_93),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_35),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_9),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g241 ( 
.A(n_105),
.B(n_26),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_178),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_40),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_184),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_23),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_63),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_49),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_119),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_67),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_41),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_60),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_111),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_165),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_117),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_115),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_45),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_195),
.A2(n_0),
.B(n_1),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_0),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_90),
.B(n_190),
.Y(n_285)
);

CKINVDCx6p67_ASAP7_75t_R g286 ( 
.A(n_221),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_223),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_200),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_201),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_263),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_225),
.A2(n_274),
.B(n_205),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_202),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_220),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_272),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_5),
.Y(n_311)
);

AOI22x1_ASAP7_75t_SL g312 ( 
.A1(n_222),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_258),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_204),
.B(n_7),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_232),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_207),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_209),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_210),
.Y(n_329)
);

BUFx8_ASAP7_75t_SL g330 ( 
.A(n_198),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_234),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_R g334 ( 
.A(n_324),
.B(n_273),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_R g335 ( 
.A(n_309),
.B(n_211),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_330),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_280),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_326),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_281),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_238),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_326),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_325),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_R g343 ( 
.A(n_307),
.B(n_304),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_294),
.B(n_248),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_245),
.Y(n_347)
);

AO21x2_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_252),
.B(n_246),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_289),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_320),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_320),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_317),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_309),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_R g357 ( 
.A(n_298),
.B(n_254),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_307),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_292),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_311),
.B(n_212),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_284),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_R g366 ( 
.A(n_328),
.B(n_213),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_323),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_323),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_214),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_290),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_283),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_283),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_295),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_308),
.A2(n_321),
.B1(n_306),
.B2(n_327),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_306),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_328),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_297),
.B(n_215),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_287),
.B(n_216),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_297),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_327),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_329),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_282),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_R g388 ( 
.A(n_287),
.B(n_218),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_219),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

AO221x1_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_363),
.B1(n_379),
.B2(n_335),
.C(n_378),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_287),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_287),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_347),
.B(n_314),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_276),
.C(n_267),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_389),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_276),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_374),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_383),
.Y(n_410)
);

BUFx6f_ASAP7_75t_SL g411 ( 
.A(n_340),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_337),
.B(n_314),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_266),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_314),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_10),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_285),
.C(n_227),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_346),
.B(n_224),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_314),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_315),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_345),
.B(n_315),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_315),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_346),
.B(n_228),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_357),
.A2(n_269),
.B1(n_230),
.B2(n_231),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_348),
.B(n_315),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_365),
.B(n_340),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_334),
.B(n_229),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_353),
.B(n_235),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_354),
.B(n_239),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_242),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_350),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_348),
.B(n_277),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_366),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_388),
.B(n_243),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_277),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_333),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_336),
.A2(n_241),
.B(n_251),
.C(n_253),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_338),
.B(n_255),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_332),
.B(n_259),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_369),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_342),
.B(n_261),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_358),
.B(n_262),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_277),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_361),
.B(n_265),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_342),
.B(n_270),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_342),
.B(n_271),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_347),
.B(n_279),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_386),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_349),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_11),
.C(n_12),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_396),
.Y(n_460)
);

AO22x1_ASAP7_75t_L g461 ( 
.A1(n_445),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_399),
.A2(n_408),
.B1(n_405),
.B2(n_395),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_410),
.B(n_13),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_394),
.B(n_15),
.C(n_16),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_431),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_15),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_16),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_322),
.B1(n_318),
.B2(n_316),
.Y(n_473)
);

NOR3xp33_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_449),
.C(n_428),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_455),
.A2(n_322),
.B1(n_318),
.B2(n_316),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_438),
.B(n_279),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_417),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_448),
.B(n_453),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_279),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_416),
.B(n_291),
.Y(n_482)
);

NOR2x2_ASAP7_75t_L g483 ( 
.A(n_411),
.B(n_17),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_291),
.Y(n_485)
);

NAND2x2_ASAP7_75t_L g486 ( 
.A(n_418),
.B(n_17),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_18),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_18),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_441),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_429),
.B(n_291),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_406),
.B(n_19),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_390),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_455),
.A2(n_322),
.B1(n_318),
.B2(n_316),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_400),
.B(n_293),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_436),
.B(n_421),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_447),
.A2(n_305),
.B1(n_302),
.B2(n_301),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_392),
.A2(n_305),
.B1(n_302),
.B2(n_301),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_293),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

BUFx4f_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_446),
.A2(n_305),
.B1(n_302),
.B2(n_301),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_400),
.B(n_293),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_404),
.B(n_293),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_404),
.B(n_296),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_414),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_432),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_450),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_401),
.Y(n_516)
);

NAND2x1p5_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_296),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_296),
.Y(n_518)
);

AO22x1_ASAP7_75t_L g519 ( 
.A1(n_427),
.A2(n_305),
.B1(n_302),
.B2(n_301),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_437),
.A2(n_299),
.B(n_21),
.C(n_22),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_402),
.B(n_299),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_437),
.A2(n_299),
.B1(n_24),
.B2(n_25),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_430),
.A2(n_299),
.B1(n_28),
.B2(n_29),
.Y(n_524)
);

BUFx8_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_415),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_490),
.B(n_439),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_471),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_479),
.B(n_422),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_498),
.A2(n_440),
.B(n_422),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_443),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_SL g535 ( 
.A1(n_472),
.A2(n_488),
.B(n_463),
.C(n_489),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_443),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_505),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_468),
.A2(n_443),
.B1(n_30),
.B2(n_31),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_499),
.A2(n_20),
.B(n_32),
.C(n_33),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_514),
.B(n_34),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_508),
.A2(n_36),
.B(n_37),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_38),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_507),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_509),
.A2(n_42),
.B(n_43),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_487),
.B(n_47),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_470),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_510),
.A2(n_53),
.B(n_54),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_477),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_525),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_R g552 ( 
.A(n_481),
.B(n_487),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_483),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_474),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_480),
.A2(n_59),
.B(n_61),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_462),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_495),
.B(n_69),
.Y(n_559)
);

AOI21xp33_ASAP7_75t_L g560 ( 
.A1(n_515),
.A2(n_71),
.B(n_72),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_523),
.A2(n_75),
.B(n_76),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_513),
.B(n_77),
.Y(n_562)
);

O2A1O1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_467),
.A2(n_81),
.B(n_83),
.C(n_87),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_88),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_485),
.A2(n_521),
.B(n_503),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_512),
.B(n_191),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_469),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_487),
.B(n_478),
.Y(n_569)
);

INVx6_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

O2A1O1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_476),
.A2(n_89),
.B(n_91),
.C(n_94),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_484),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_492),
.B(n_500),
.Y(n_573)
);

O2A1O1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_482),
.A2(n_96),
.B(n_97),
.C(n_100),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_522),
.A2(n_520),
.B(n_473),
.C(n_504),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_522),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_526),
.A2(n_104),
.B(n_106),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_494),
.B(n_109),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_461),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_473),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_524),
.B(n_118),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_517),
.B(n_120),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_497),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_528),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_565),
.A2(n_533),
.B(n_561),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_579),
.A2(n_556),
.B(n_564),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_539),
.B(n_494),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_531),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_546),
.Y(n_592)
);

AO21x2_ASAP7_75t_L g593 ( 
.A1(n_575),
.A2(n_491),
.B(n_518),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_582),
.Y(n_595)
);

BUFx6f_ASAP7_75t_SL g596 ( 
.A(n_551),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_582),
.Y(n_597)
);

AO21x2_ASAP7_75t_L g598 ( 
.A1(n_535),
.A2(n_497),
.B(n_475),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_568),
.Y(n_600)
);

AOI22x1_ASAP7_75t_L g601 ( 
.A1(n_554),
.A2(n_504),
.B1(n_493),
.B2(n_506),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_501),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_532),
.A2(n_519),
.B(n_123),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_534),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_542),
.A2(n_121),
.B(n_124),
.Y(n_605)
);

BUFx2_ASAP7_75t_R g606 ( 
.A(n_562),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_568),
.B(n_125),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_545),
.A2(n_126),
.B(n_128),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_572),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_189),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_549),
.A2(n_129),
.B(n_131),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_537),
.B(n_133),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_567),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_557),
.A2(n_134),
.B(n_135),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_536),
.B(n_569),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_583),
.A2(n_136),
.B(n_138),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_574),
.A2(n_577),
.B(n_540),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_569),
.B(n_140),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_571),
.A2(n_141),
.B(n_144),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_547),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_541),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_563),
.A2(n_145),
.B(n_146),
.Y(n_627)
);

OA21x2_ASAP7_75t_L g628 ( 
.A1(n_576),
.A2(n_148),
.B(n_152),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_543),
.B(n_153),
.Y(n_629)
);

BUFx2_ASAP7_75t_SL g630 ( 
.A(n_550),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_538),
.A2(n_155),
.B(n_158),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_584),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_618),
.A2(n_573),
.B1(n_566),
.B2(n_581),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_614),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_548),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_586),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_620),
.A2(n_570),
.B1(n_560),
.B2(n_163),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_633),
.B(n_570),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_589),
.B(n_159),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_599),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_614),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_596),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_597),
.Y(n_645)
);

BUFx6f_ASAP7_75t_SL g646 ( 
.A(n_595),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_624),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_619),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_600),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_588),
.A2(n_162),
.B(n_164),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_591),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_630),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

BUFx8_ASAP7_75t_SL g654 ( 
.A(n_596),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_619),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_604),
.B(n_188),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_600),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_588),
.A2(n_174),
.B(n_176),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_597),
.Y(n_659)
);

BUFx8_ASAP7_75t_L g660 ( 
.A(n_595),
.Y(n_660)
);

NOR2x1_ASAP7_75t_SL g661 ( 
.A(n_613),
.B(n_177),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_615),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_610),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_626),
.A2(n_632),
.B1(n_585),
.B2(n_608),
.Y(n_665)
);

AO21x2_ASAP7_75t_L g666 ( 
.A1(n_603),
.A2(n_183),
.B(n_185),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_613),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_617),
.B(n_186),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_626),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_632),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_593),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_602),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_592),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_632),
.Y(n_675)
);

AOI21x1_ASAP7_75t_L g676 ( 
.A1(n_587),
.A2(n_629),
.B(n_621),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_600),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_663),
.Y(n_678)
);

NAND2x1_ASAP7_75t_L g679 ( 
.A(n_636),
.B(n_625),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_637),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_653),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_R g682 ( 
.A(n_669),
.B(n_611),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_644),
.B(n_590),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_653),
.B(n_622),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_SL g685 ( 
.A(n_639),
.B(n_638),
.C(n_669),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_659),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_663),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_R g688 ( 
.A(n_659),
.B(n_660),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_634),
.A2(n_616),
.B(n_636),
.C(n_631),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_651),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_R g691 ( 
.A(n_647),
.B(n_628),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_643),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_647),
.B(n_667),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_674),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_664),
.B(n_641),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_654),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_657),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_662),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_654),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_648),
.Y(n_701)
);

AND2x6_ASAP7_75t_L g702 ( 
.A(n_636),
.B(n_607),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_653),
.B(n_602),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_645),
.B(n_607),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_646),
.B(n_641),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_657),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_655),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_670),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_643),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_673),
.B(n_602),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_640),
.B(n_590),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_643),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_640),
.B(n_606),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_673),
.A2(n_628),
.B1(n_601),
.B2(n_616),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

NOR3xp33_ASAP7_75t_SL g718 ( 
.A(n_652),
.B(n_627),
.C(n_621),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_R g719 ( 
.A(n_660),
.B(n_602),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_665),
.B(n_602),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_646),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_647),
.B(n_598),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_673),
.A2(n_598),
.B1(n_631),
.B2(n_627),
.Y(n_724)
);

INVx11_ASAP7_75t_L g725 ( 
.A(n_660),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_646),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_649),
.B(n_587),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_657),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_680),
.B(n_673),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_694),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_711),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_727),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_690),
.B(n_673),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_723),
.B(n_671),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_696),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_678),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_709),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_715),
.A2(n_721),
.B1(n_702),
.B2(n_703),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_717),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_687),
.B(n_649),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_711),
.B(n_677),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_701),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_720),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_699),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_706),
.B(n_676),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_714),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_683),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_706),
.B(n_677),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_679),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_708),
.B(n_677),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_681),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_708),
.B(n_677),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_728),
.B(n_672),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_728),
.B(n_661),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_686),
.B(n_656),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_681),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_703),
.B(n_635),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_702),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_702),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_704),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_722),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_738),
.B(n_686),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_732),
.B(n_689),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_730),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_736),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_761),
.B(n_704),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_758),
.B(n_684),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_743),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_743),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_744),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_744),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_745),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_732),
.B(n_724),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_745),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_755),
.B(n_718),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_749),
.B(n_722),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_748),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_740),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_748),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_761),
.B(n_762),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_746),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_735),
.B(n_704),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_735),
.B(n_758),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_746),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_755),
.B(n_698),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_741),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_741),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_766),
.B(n_734),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_786),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_770),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_780),
.B(n_747),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_765),
.B(n_751),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_789),
.B(n_734),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_765),
.B(n_705),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_788),
.B(n_731),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_779),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_770),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_790),
.B(n_762),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_772),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_788),
.B(n_764),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_774),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_779),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_774),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_767),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_793),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_797),
.A2(n_691),
.B1(n_778),
.B2(n_761),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_797),
.A2(n_775),
.B1(n_777),
.B2(n_693),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_795),
.A2(n_775),
.B1(n_777),
.B2(n_739),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_800),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_795),
.B(n_785),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_792),
.B(n_768),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_794),
.B(n_784),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_799),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_791),
.A2(n_759),
.B1(n_760),
.B2(n_684),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_809),
.A2(n_794),
.B(n_807),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_813),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_810),
.A2(n_769),
.B(n_808),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_819),
.Y(n_823)
);

AOI21xp33_ASAP7_75t_SL g824 ( 
.A1(n_815),
.A2(n_763),
.B(n_697),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_821),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_823),
.B(n_812),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_820),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_822),
.B(n_816),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_824),
.B(n_688),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_827),
.B(n_811),
.C(n_820),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_828),
.B(n_685),
.C(n_763),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_826),
.B(n_814),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_825),
.Y(n_833)
);

AOI211xp5_ASAP7_75t_L g834 ( 
.A1(n_830),
.A2(n_829),
.B(n_682),
.C(n_710),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_833),
.B(n_814),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_831),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_834),
.A2(n_832),
.B(n_716),
.C(n_713),
.Y(n_837)
);

NOR2x1p5_ASAP7_75t_L g838 ( 
.A(n_835),
.B(n_700),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_836),
.A2(n_692),
.B1(n_756),
.B2(n_726),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_838),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_837),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_836),
.Y(n_842)
);

AO211x2_ASAP7_75t_L g843 ( 
.A1(n_837),
.A2(n_760),
.B(n_787),
.C(n_783),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_836),
.A2(n_756),
.B1(n_818),
.B2(n_712),
.Y(n_844)
);

AOI222xp33_ASAP7_75t_L g845 ( 
.A1(n_841),
.A2(n_842),
.B1(n_843),
.B2(n_840),
.C1(n_716),
.C2(n_839),
.Y(n_845)
);

INVxp33_ASAP7_75t_L g846 ( 
.A(n_844),
.Y(n_846)
);

OAI211xp5_ASAP7_75t_L g847 ( 
.A1(n_842),
.A2(n_725),
.B(n_719),
.C(n_792),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_840),
.B(n_803),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_840),
.B(n_798),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_842),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_842),
.B(n_668),
.C(n_623),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_850),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_848),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_849),
.B(n_847),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_845),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_851),
.B(n_784),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_846),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_850),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_853),
.Y(n_859)
);

XOR2xp5_ASAP7_75t_L g860 ( 
.A(n_857),
.B(n_768),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_852),
.B(n_769),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_858),
.Y(n_862)
);

NAND4xp25_ASAP7_75t_L g863 ( 
.A(n_854),
.B(n_753),
.C(n_784),
.D(n_750),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_854),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_855),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_856),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_856),
.A2(n_776),
.B(n_773),
.Y(n_867)
);

AOI31xp33_ASAP7_75t_L g868 ( 
.A1(n_859),
.A2(n_796),
.A3(n_768),
.B(n_771),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_864),
.B(n_804),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_865),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_862),
.B(n_805),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_866),
.A2(n_817),
.B1(n_801),
.B2(n_750),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_860),
.Y(n_873)
);

OAI31xp33_ASAP7_75t_L g874 ( 
.A1(n_861),
.A2(n_729),
.A3(n_733),
.B(n_782),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_863),
.A2(n_666),
.B1(n_754),
.B2(n_752),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_867),
.A2(n_666),
.B1(n_754),
.B2(n_752),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_870),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_875),
.A2(n_733),
.B1(n_729),
.B2(n_698),
.Y(n_878)
);

OAI22x1_ASAP7_75t_L g879 ( 
.A1(n_873),
.A2(n_782),
.B1(n_742),
.B2(n_731),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_876),
.A2(n_698),
.B1(n_782),
.B2(n_806),
.Y(n_880)
);

AOI22x1_ASAP7_75t_L g881 ( 
.A1(n_869),
.A2(n_650),
.B1(n_658),
.B2(n_731),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_877),
.A2(n_871),
.B1(n_872),
.B2(n_868),
.Y(n_882)
);

AOI222xp33_ASAP7_75t_SL g883 ( 
.A1(n_879),
.A2(n_874),
.B1(n_658),
.B2(n_650),
.C1(n_623),
.C2(n_737),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_L g884 ( 
.A(n_883),
.B(n_878),
.C(n_880),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_884),
.A2(n_882),
.B1(n_881),
.B2(n_642),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_885),
.B(n_605),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_886),
.A2(n_609),
.B1(n_612),
.B2(n_781),
.Y(n_887)
);


endmodule