module real_aes_1460_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_784, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_784;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g178 ( .A(n_0), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_1), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_2), .B(n_184), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_3), .B(n_181), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_4), .A2(n_44), .B1(n_767), .B2(n_768), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_4), .Y(n_767) );
INVx1_ASAP7_75t_L g144 ( .A(n_5), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_6), .B(n_184), .Y(n_206) );
NAND2xp33_ASAP7_75t_SL g164 ( .A(n_7), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g135 ( .A(n_8), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_9), .Y(n_778) );
AND2x2_ASAP7_75t_L g204 ( .A(n_10), .B(n_187), .Y(n_204) );
AND2x2_ASAP7_75t_L g475 ( .A(n_11), .B(n_160), .Y(n_475) );
AND2x2_ASAP7_75t_L g526 ( .A(n_12), .B(n_215), .Y(n_526) );
INVx2_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_14), .B(n_181), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_15), .B(n_777), .C(n_779), .Y(n_776) );
AOI221x1_ASAP7_75t_L g156 ( .A1(n_16), .A2(n_157), .B1(n_159), .B2(n_160), .C(n_163), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_17), .B(n_184), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_18), .B(n_184), .Y(n_531) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_20), .A2(n_90), .B1(n_139), .B2(n_184), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_21), .A2(n_159), .B(n_208), .Y(n_207) );
AOI221xp5_ASAP7_75t_SL g251 ( .A1(n_22), .A2(n_36), .B1(n_159), .B2(n_184), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_23), .B(n_179), .Y(n_209) );
OR2x2_ASAP7_75t_L g137 ( .A(n_24), .B(n_89), .Y(n_137) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_24), .A2(n_89), .B(n_138), .Y(n_162) );
INVxp67_ASAP7_75t_L g155 ( .A(n_25), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_26), .B(n_181), .Y(n_246) );
AND2x2_ASAP7_75t_L g198 ( .A(n_27), .B(n_186), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_28), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_29), .A2(n_159), .B(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_30), .A2(n_160), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_31), .B(n_181), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_32), .A2(n_159), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_33), .B(n_181), .Y(n_507) );
AND2x2_ASAP7_75t_L g146 ( .A(n_34), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g150 ( .A(n_34), .Y(n_150) );
AND2x2_ASAP7_75t_L g165 ( .A(n_34), .B(n_144), .Y(n_165) );
OR2x6_ASAP7_75t_L g115 ( .A(n_35), .B(n_116), .Y(n_115) );
INVxp67_ASAP7_75t_L g779 ( .A(n_35), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_37), .B(n_184), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_38), .A2(n_81), .B1(n_148), .B2(n_159), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_39), .B(n_181), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_40), .A2(n_49), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_41), .B(n_184), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_42), .B(n_179), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_43), .A2(n_159), .B(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_44), .Y(n_768) );
AND2x2_ASAP7_75t_L g185 ( .A(n_45), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_46), .B(n_179), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_47), .B(n_186), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_48), .B(n_184), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_49), .Y(n_122) );
INVx1_ASAP7_75t_L g142 ( .A(n_50), .Y(n_142) );
INVx1_ASAP7_75t_L g169 ( .A(n_50), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_51), .B(n_181), .Y(n_473) );
AND2x2_ASAP7_75t_L g485 ( .A(n_52), .B(n_186), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_53), .B(n_184), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_54), .B(n_179), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_55), .B(n_179), .Y(n_506) );
AND2x2_ASAP7_75t_L g227 ( .A(n_56), .B(n_186), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_57), .B(n_184), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_58), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_59), .B(n_184), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_60), .A2(n_159), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_61), .B(n_179), .Y(n_225) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_62), .B(n_187), .Y(n_247) );
AND2x2_ASAP7_75t_L g537 ( .A(n_63), .B(n_187), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_64), .A2(n_159), .B(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_65), .B(n_181), .Y(n_210) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_66), .B(n_215), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_67), .B(n_179), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_68), .B(n_179), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_69), .A2(n_92), .B1(n_148), .B2(n_159), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_70), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_71), .B(n_181), .Y(n_534) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g171 ( .A(n_72), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_73), .B(n_179), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_74), .A2(n_159), .B(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_75), .A2(n_159), .B(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_76), .A2(n_159), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g509 ( .A(n_77), .B(n_187), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_78), .B(n_186), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_79), .A2(n_83), .B1(n_139), .B2(n_184), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_80), .B(n_184), .Y(n_226) );
INVx1_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_82), .B(n_117), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_84), .B(n_179), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_85), .B(n_179), .Y(n_254) );
AND2x2_ASAP7_75t_L g466 ( .A(n_86), .B(n_215), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_87), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_88), .A2(n_159), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_91), .B(n_181), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_93), .A2(n_159), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_94), .B(n_181), .Y(n_464) );
INVxp67_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_96), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_97), .B(n_181), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_98), .A2(n_159), .B(n_244), .Y(n_243) );
BUFx2_ASAP7_75t_L g536 ( .A(n_99), .Y(n_536) );
BUFx2_ASAP7_75t_L g107 ( .A(n_100), .Y(n_107) );
BUFx2_ASAP7_75t_SL g759 ( .A(n_100), .Y(n_759) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_770), .B(n_780), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_120), .B(n_757), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_109), .A2(n_761), .B(n_764), .Y(n_760) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_119), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_R g763 ( .A(n_112), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_113), .B(n_115), .Y(n_126) );
OR2x6_ASAP7_75t_SL g453 ( .A(n_113), .B(n_114), .Y(n_453) );
OR2x2_ASAP7_75t_L g756 ( .A(n_113), .B(n_115), .Y(n_756) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B(n_748), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_121), .A2(n_749), .B(n_752), .Y(n_748) );
OA22x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_127), .B1(n_450), .B2(n_454), .Y(n_124) );
OAI22x1_ASAP7_75t_L g749 ( .A1(n_125), .A2(n_451), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx11_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g750 ( .A(n_127), .Y(n_750) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_127), .A2(n_765), .B1(n_766), .B2(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_127), .Y(n_765) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_327), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_270), .C(n_309), .D(n_316), .Y(n_128) );
OAI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_188), .B1(n_228), .B2(n_237), .C(n_256), .Y(n_129) );
OR2x2_ASAP7_75t_L g400 ( .A(n_130), .B(n_262), .Y(n_400) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g315 ( .A(n_131), .B(n_240), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_131), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_131), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_172), .Y(n_131) );
AND2x4_ASAP7_75t_SL g239 ( .A(n_132), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g261 ( .A(n_132), .Y(n_261) );
AND2x2_ASAP7_75t_L g296 ( .A(n_132), .B(n_269), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_132), .B(n_173), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_132), .B(n_263), .Y(n_348) );
OR2x2_ASAP7_75t_L g426 ( .A(n_132), .B(n_240), .Y(n_426) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_156), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B1(n_148), .B2(n_154), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_136), .B(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_136), .B(n_158), .Y(n_157) );
NOR3xp33_ASAP7_75t_L g163 ( .A(n_136), .B(n_164), .C(n_166), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_136), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_136), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_136), .A2(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_137), .B(n_138), .Y(n_187) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g153 ( .A(n_142), .B(n_144), .Y(n_153) );
AND2x4_ASAP7_75t_L g181 ( .A(n_142), .B(n_170), .Y(n_181) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g159 ( .A(n_146), .B(n_153), .Y(n_159) );
INVx2_ASAP7_75t_L g152 ( .A(n_147), .Y(n_152) );
AND2x6_ASAP7_75t_L g179 ( .A(n_147), .B(n_168), .Y(n_179) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g502 ( .A(n_160), .Y(n_502) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_161), .A2(n_175), .B(n_185), .Y(n_174) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_161), .A2(n_469), .B(n_475), .Y(n_468) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx4f_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx5_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
AND2x4_ASAP7_75t_L g184 ( .A(n_165), .B(n_167), .Y(n_184) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g248 ( .A(n_173), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_173), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g274 ( .A(n_173), .Y(n_274) );
OR2x2_ASAP7_75t_L g279 ( .A(n_173), .B(n_263), .Y(n_279) );
AND2x2_ASAP7_75t_L g292 ( .A(n_173), .B(n_250), .Y(n_292) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_173), .Y(n_295) );
INVx1_ASAP7_75t_L g307 ( .A(n_173), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_173), .B(n_261), .Y(n_372) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_183), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .B(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_179), .B(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_182), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_182), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_182), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_182), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_182), .A2(n_253), .B(n_254), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_182), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_182), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_182), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_182), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_182), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_182), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_182), .A2(n_534), .B(n_535), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_186), .Y(n_197) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_186), .A2(n_251), .B(n_255), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_186), .A2(n_461), .B(n_462), .Y(n_460) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_186), .A2(n_479), .B(n_480), .Y(n_478) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_189), .B(n_199), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g236 ( .A(n_190), .B(n_220), .Y(n_236) );
AND2x4_ASAP7_75t_L g266 ( .A(n_190), .B(n_203), .Y(n_266) );
INVx2_ASAP7_75t_L g300 ( .A(n_190), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_190), .B(n_220), .Y(n_358) );
AND2x2_ASAP7_75t_L g405 ( .A(n_190), .B(n_234), .Y(n_405) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_197), .B(n_198), .Y(n_190) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_191), .A2(n_197), .B(n_198), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_196), .Y(n_191) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_197), .A2(n_221), .B(n_227), .Y(n_220) );
AOI21x1_ASAP7_75t_L g519 ( .A1(n_197), .A2(n_520), .B(n_526), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g393 ( .A1(n_199), .A2(n_265), .B1(n_308), .B2(n_368), .C1(n_394), .C2(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g312 ( .A(n_201), .B(n_232), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_201), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g441 ( .A(n_201), .B(n_281), .Y(n_441) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_202), .A2(n_272), .B(n_276), .Y(n_271) );
AND2x2_ASAP7_75t_L g352 ( .A(n_202), .B(n_235), .Y(n_352) );
OR2x2_ASAP7_75t_L g377 ( .A(n_202), .B(n_236), .Y(n_377) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx5_ASAP7_75t_L g231 ( .A(n_203), .Y(n_231) );
AND2x2_ASAP7_75t_L g318 ( .A(n_203), .B(n_300), .Y(n_318) );
AND2x2_ASAP7_75t_L g344 ( .A(n_203), .B(n_220), .Y(n_344) );
OR2x2_ASAP7_75t_L g347 ( .A(n_203), .B(n_234), .Y(n_347) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_203), .Y(n_365) );
AND2x4_ASAP7_75t_SL g422 ( .A(n_203), .B(n_299), .Y(n_422) );
OR2x2_ASAP7_75t_L g431 ( .A(n_203), .B(n_258), .Y(n_431) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
AOI221xp5_ASAP7_75t_SL g382 ( .A1(n_211), .A2(n_266), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_382) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_220), .Y(n_211) );
OR2x2_ASAP7_75t_L g321 ( .A(n_212), .B(n_291), .Y(n_321) );
OR2x2_ASAP7_75t_L g331 ( .A(n_212), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g357 ( .A(n_212), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g363 ( .A(n_212), .B(n_282), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_212), .B(n_346), .Y(n_375) );
INVx2_ASAP7_75t_L g388 ( .A(n_212), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_212), .B(n_266), .Y(n_409) );
AND2x2_ASAP7_75t_L g413 ( .A(n_212), .B(n_235), .Y(n_413) );
AND2x2_ASAP7_75t_L g421 ( .A(n_212), .B(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
AOI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_216), .B(n_219), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_215), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_215), .A2(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_220), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g265 ( .A(n_220), .B(n_234), .Y(n_265) );
INVx2_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
AND2x4_ASAP7_75t_L g299 ( .A(n_220), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_220), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_232), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g411 ( .A(n_230), .B(n_233), .Y(n_411) );
AND2x4_ASAP7_75t_L g257 ( .A(n_231), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g298 ( .A(n_231), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g325 ( .A(n_231), .B(n_265), .Y(n_325) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g429 ( .A(n_233), .B(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g281 ( .A(n_234), .B(n_282), .Y(n_281) );
OAI21xp5_ASAP7_75t_SL g301 ( .A1(n_235), .A2(n_302), .B(n_308), .Y(n_301) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
INVx1_ASAP7_75t_SL g355 ( .A(n_239), .Y(n_355) );
AND2x2_ASAP7_75t_L g385 ( .A(n_239), .B(n_295), .Y(n_385) );
AND2x4_ASAP7_75t_L g396 ( .A(n_239), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g262 ( .A(n_240), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g269 ( .A(n_240), .Y(n_269) );
AND2x4_ASAP7_75t_L g275 ( .A(n_240), .B(n_261), .Y(n_275) );
INVx2_ASAP7_75t_L g286 ( .A(n_240), .Y(n_286) );
INVx1_ASAP7_75t_L g335 ( .A(n_240), .Y(n_335) );
OR2x2_ASAP7_75t_L g356 ( .A(n_240), .B(n_340), .Y(n_356) );
OR2x2_ASAP7_75t_L g370 ( .A(n_240), .B(n_250), .Y(n_370) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_240), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_240), .B(n_292), .Y(n_442) );
OR2x6_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
INVx1_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
AND2x2_ASAP7_75t_L g420 ( .A(n_248), .B(n_286), .Y(n_420) );
AND2x2_ASAP7_75t_L g445 ( .A(n_248), .B(n_275), .Y(n_445) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g263 ( .A(n_250), .Y(n_263) );
BUFx3_ASAP7_75t_L g305 ( .A(n_250), .Y(n_305) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
INVx1_ASAP7_75t_L g341 ( .A(n_250), .Y(n_341) );
AOI33xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_259), .A3(n_264), .B1(n_265), .B2(n_266), .B3(n_267), .Y(n_256) );
AOI21x1_ASAP7_75t_SL g359 ( .A1(n_257), .A2(n_281), .B(n_343), .Y(n_359) );
INVx2_ASAP7_75t_L g389 ( .A(n_257), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_257), .B(n_388), .Y(n_395) );
AND2x2_ASAP7_75t_L g343 ( .A(n_258), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g306 ( .A(n_261), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g407 ( .A(n_262), .Y(n_407) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
OAI32xp33_ASAP7_75t_L g446 ( .A1(n_264), .A2(n_266), .A3(n_442), .B1(n_447), .B2(n_449), .Y(n_446) );
AND2x2_ASAP7_75t_L g364 ( .A(n_265), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g354 ( .A(n_266), .Y(n_354) );
AND2x2_ASAP7_75t_L g419 ( .A(n_266), .B(n_363), .Y(n_419) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI221xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_280), .B1(n_283), .B2(n_297), .C(n_301), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_274), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_275), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_275), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_275), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g324 ( .A(n_279), .Y(n_324) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR3xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .C(n_293), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_285), .A2(n_347), .B1(n_387), .B2(n_390), .Y(n_386) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g290 ( .A(n_286), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g304 ( .A(n_286), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_286), .Y(n_326) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI322xp33_ASAP7_75t_L g353 ( .A1(n_289), .A2(n_331), .A3(n_354), .B1(n_355), .B2(n_356), .C1(n_357), .C2(n_359), .Y(n_353) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_291), .A2(n_310), .B(n_311), .C(n_313), .Y(n_309) );
OR2x2_ASAP7_75t_L g401 ( .A(n_291), .B(n_355), .Y(n_401) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_296), .Y(n_308) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g314 ( .A(n_298), .B(n_315), .Y(n_314) );
INVx3_ASAP7_75t_SL g346 ( .A(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_303), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g350 ( .A(n_306), .Y(n_350) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_307), .Y(n_392) );
OR2x6_ASAP7_75t_SL g447 ( .A(n_310), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_315), .A2(n_438), .B(n_439), .C(n_446), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_319), .B(n_322), .C(n_326), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g328 ( .A1(n_317), .A2(n_329), .B(n_336), .C(n_360), .Y(n_328) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_373), .C(n_417), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_332), .Y(n_424) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
NOR3xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_349), .C(n_353), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B1(n_345), .B2(n_348), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_341), .Y(n_448) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_SL g434 ( .A(n_347), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OR2x2_ASAP7_75t_L g384 ( .A(n_350), .B(n_370), .Y(n_384) );
OR2x2_ASAP7_75t_L g435 ( .A(n_350), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g433 ( .A(n_358), .Y(n_433) );
OR2x2_ASAP7_75t_L g449 ( .A(n_358), .B(n_388), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_366), .Y(n_360) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_361), .A2(n_375), .A3(n_376), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g406 ( .A(n_371), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND4xp25_ASAP7_75t_SL g373 ( .A(n_374), .B(n_382), .C(n_393), .D(n_398), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_398) );
NAND2xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g443 ( .A(n_402), .Y(n_443) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g438 ( .A(n_412), .Y(n_438) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_418), .B(n_437), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_423), .C(n_427), .Y(n_418) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_432), .B(n_435), .Y(n_427) );
INVxp33_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx4f_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
CKINVDCx11_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_SL g751 ( .A(n_454), .Y(n_751) );
AND2x4_ASAP7_75t_SL g454 ( .A(n_455), .B(n_644), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_553), .C(n_585), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_481), .B1(n_510), .B2(n_527), .C(n_538), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g516 ( .A(n_459), .B(n_468), .Y(n_516) );
INVx4_ASAP7_75t_L g544 ( .A(n_459), .Y(n_544) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_459), .B(n_518), .Y(n_584) );
BUFx2_ASAP7_75t_L g594 ( .A(n_459), .Y(n_594) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_459), .B(n_599), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_459), .B(n_597), .Y(n_669) );
OR2x2_ASAP7_75t_L g677 ( .A(n_459), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g703 ( .A(n_459), .B(n_542), .Y(n_703) );
AND2x4_ASAP7_75t_L g722 ( .A(n_459), .B(n_723), .Y(n_722) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .Y(n_459) );
INVx2_ASAP7_75t_SL g635 ( .A(n_467), .Y(n_635) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_476), .Y(n_467) );
AND2x2_ASAP7_75t_L g542 ( .A(n_468), .B(n_519), .Y(n_542) );
INVx2_ASAP7_75t_L g569 ( .A(n_468), .Y(n_569) );
INVx2_ASAP7_75t_L g599 ( .A(n_468), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_468), .B(n_518), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
AND2x2_ASAP7_75t_L g543 ( .A(n_476), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
BUFx3_ASAP7_75t_L g580 ( .A(n_476), .Y(n_580) );
AND2x2_ASAP7_75t_L g609 ( .A(n_476), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x4_ASAP7_75t_L g514 ( .A(n_477), .B(n_478), .Y(n_514) );
INVx1_ASAP7_75t_L g615 ( .A(n_481), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
OR2x2_ASAP7_75t_L g726 ( .A(n_482), .B(n_527), .Y(n_726) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g582 ( .A(n_483), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_483), .B(n_492), .Y(n_643) );
OR2x2_ASAP7_75t_L g741 ( .A(n_483), .B(n_663), .Y(n_741) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g552 ( .A(n_484), .B(n_528), .Y(n_552) );
OR2x2_ASAP7_75t_SL g562 ( .A(n_484), .B(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_484), .Y(n_624) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_484), .B(n_529), .Y(n_630) );
AND2x2_ASAP7_75t_L g655 ( .A(n_484), .B(n_494), .Y(n_655) );
OR2x2_ASAP7_75t_L g676 ( .A(n_484), .B(n_559), .Y(n_676) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g571 ( .A(n_492), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_492), .A2(n_665), .B(n_668), .C(n_670), .Y(n_664) );
AND2x2_ASAP7_75t_L g737 ( .A(n_492), .B(n_513), .Y(n_737) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
INVx1_ASAP7_75t_L g604 ( .A(n_493), .Y(n_604) );
AND2x2_ASAP7_75t_L g674 ( .A(n_493), .B(n_529), .Y(n_674) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g548 ( .A(n_494), .Y(n_548) );
OR2x2_ASAP7_75t_L g563 ( .A(n_494), .B(n_529), .Y(n_563) );
INVx1_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_494), .B(n_501), .Y(n_591) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_494), .Y(n_697) );
NOR2x1_ASAP7_75t_SL g528 ( .A(n_501), .B(n_529), .Y(n_528) );
AO21x1_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B(n_509), .Y(n_501) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_503), .B(n_509), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_508), .Y(n_503) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
OR2x2_ASAP7_75t_L g661 ( .A(n_512), .B(n_596), .Y(n_661) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_513), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g743 ( .A(n_513), .B(n_640), .Y(n_743) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_569), .Y(n_588) );
AND2x2_ASAP7_75t_L g684 ( .A(n_514), .B(n_597), .Y(n_684) );
INVx1_ASAP7_75t_L g601 ( .A(n_515), .Y(n_601) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g651 ( .A(n_516), .Y(n_651) );
INVx2_ASAP7_75t_L g618 ( .A(n_517), .Y(n_618) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g568 ( .A(n_518), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g598 ( .A(n_518), .Y(n_598) );
INVx1_ASAP7_75t_L g723 ( .A(n_518), .Y(n_723) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_519), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
OR2x2_ASAP7_75t_L g694 ( .A(n_527), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g549 ( .A(n_529), .Y(n_549) );
OR2x2_ASAP7_75t_L g572 ( .A(n_529), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g583 ( .A(n_529), .B(n_559), .Y(n_583) );
AND2x2_ASAP7_75t_L g657 ( .A(n_529), .B(n_573), .Y(n_657) );
BUFx2_ASAP7_75t_L g740 ( .A(n_529), .Y(n_740) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_537), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_545), .B(n_550), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_L g692 ( .A(n_541), .B(n_614), .Y(n_692) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g551 ( .A(n_542), .B(n_544), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_543), .B(n_613), .Y(n_714) );
INVx1_ASAP7_75t_L g744 ( .A(n_543), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_544), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_544), .B(n_680), .Y(n_717) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_547), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_547), .B(n_575), .Y(n_728) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_548), .B(n_630), .Y(n_686) );
AND2x2_ASAP7_75t_L g704 ( .A(n_548), .B(n_657), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_549), .B(n_591), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_549), .A2(n_595), .B(n_637), .C(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_549), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_551), .A2(n_624), .B1(n_732), .B2(n_738), .C(n_742), .Y(n_731) );
INVx1_ASAP7_75t_SL g719 ( .A(n_552), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_564), .B1(n_570), .B2(n_574), .C(n_784), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g629 ( .A(n_558), .Y(n_629) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g603 ( .A(n_559), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g634 ( .A(n_559), .B(n_579), .Y(n_634) );
INVx2_ASAP7_75t_L g667 ( .A(n_559), .Y(n_667) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_562), .A2(n_609), .A3(n_640), .B1(n_719), .B2(n_720), .Y(n_718) );
OR2x2_ASAP7_75t_L g689 ( .A(n_563), .B(n_676), .Y(n_689) );
INVx1_ASAP7_75t_L g699 ( .A(n_564), .Y(n_699) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx2_ASAP7_75t_L g614 ( .A(n_565), .Y(n_614) );
AND2x2_ASAP7_75t_L g685 ( .A(n_565), .B(n_660), .Y(n_685) );
OR2x2_ASAP7_75t_L g716 ( .A(n_565), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_566), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g610 ( .A(n_569), .Y(n_610) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_SL g575 ( .A(n_572), .Y(n_575) );
OR2x2_ASAP7_75t_L g662 ( .A(n_572), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_573), .B(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_573), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g709 ( .A(n_573), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_581), .C(n_584), .Y(n_574) );
AND2x2_ASAP7_75t_L g724 ( .A(n_576), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g650 ( .A(n_580), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_580), .B(n_584), .Y(n_671) );
AND2x2_ASAP7_75t_L g702 ( .A(n_580), .B(n_703), .Y(n_702) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_582), .A2(n_713), .B(n_715), .C(n_718), .Y(n_712) );
AOI222xp33_ASAP7_75t_L g586 ( .A1(n_583), .A2(n_587), .B1(n_589), .B2(n_592), .C1(n_600), .C2(n_602), .Y(n_586) );
AND2x2_ASAP7_75t_L g654 ( .A(n_583), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g587 ( .A(n_584), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_SL g608 ( .A(n_584), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_605), .C(n_626), .D(n_636), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_588), .B(n_594), .Y(n_648) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g656 ( .A(n_591), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_SL g663 ( .A(n_591), .Y(n_663) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_593), .A2(n_627), .B(n_631), .C(n_635), .Y(n_626) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_594), .B(n_609), .Y(n_730) );
OR2x2_ASAP7_75t_L g734 ( .A(n_594), .B(n_620), .Y(n_734) );
INVx1_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_SL g641 ( .A(n_598), .Y(n_641) );
INVx1_ASAP7_75t_L g621 ( .A(n_599), .Y(n_621) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_601), .B(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g625 ( .A(n_603), .Y(n_625) );
AOI322xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .A3(n_609), .B1(n_611), .B2(n_615), .C1(n_616), .C2(n_622), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_SL g687 ( .A1(n_608), .A2(n_688), .B(n_689), .C(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g710 ( .A(n_609), .Y(n_710) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g668 ( .A(n_614), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_620), .Y(n_690) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx3_ASAP7_75t_L g633 ( .A(n_630), .Y(n_633) );
OR2x2_ASAP7_75t_L g701 ( .A(n_630), .B(n_663), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_630), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_SL g733 ( .A(n_634), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_635), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g738 ( .A(n_643), .B(n_739), .C(n_741), .Y(n_738) );
NOR3xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_682), .C(n_711), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_664), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_652), .C(n_658), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g691 ( .A1(n_647), .A2(n_669), .A3(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx2_ASAP7_75t_L g706 ( .A(n_654), .Y(n_706) );
INVx1_ASAP7_75t_L g681 ( .A(n_656), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g708 ( .A(n_666), .B(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g747 ( .A(n_667), .Y(n_747) );
OAI22xp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_672), .B1(n_677), .B2(n_681), .Y(n_670) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_676), .Y(n_688) );
OR2x2_ASAP7_75t_L g739 ( .A(n_676), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_691), .C(n_698), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B(n_686), .C(n_687), .Y(n_683) );
INVx2_ASAP7_75t_L g720 ( .A(n_684), .Y(n_720) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_710), .Y(n_705) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_712), .B(n_721), .C(n_731), .Y(n_711) );
INVxp33_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_727), .B2(n_729), .Y(n_721) );
INVx2_ASAP7_75t_L g735 ( .A(n_722), .Y(n_735) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp33_ASAP7_75t_SL g742 ( .A1(n_741), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_766), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx3_ASAP7_75t_SL g782 ( .A(n_773), .Y(n_782) );
INVx3_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_SL g774 ( .A(n_775), .B(n_776), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
endmodule