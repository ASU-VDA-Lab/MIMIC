module fake_jpeg_11614_n_522 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_522);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_522;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_20),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_2),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_1),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_41),
.Y(n_147)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_101),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_38),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_19),
.B1(n_23),
.B2(n_44),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_121),
.A2(n_49),
.B1(n_8),
.B2(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_128),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_23),
.B1(n_37),
.B2(n_39),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_127),
.A2(n_129),
.B1(n_133),
.B2(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_48),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_51),
.A2(n_23),
.B1(n_39),
.B2(n_27),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_53),
.A2(n_39),
.B1(n_18),
.B2(n_27),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_60),
.A2(n_39),
.B1(n_22),
.B2(n_27),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_137),
.A2(n_49),
.B1(n_4),
.B2(n_6),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_62),
.A2(n_65),
.B1(n_64),
.B2(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_48),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_147),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_54),
.A2(n_28),
.B1(n_61),
.B2(n_58),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_148),
.B1(n_93),
.B2(n_92),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_98),
.A2(n_28),
.B1(n_40),
.B2(n_97),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_72),
.B(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_19),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_47),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_162),
.Y(n_221)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_163),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_165),
.B(n_174),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_166),
.A2(n_169),
.B1(n_172),
.B2(n_213),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_89),
.B(n_82),
.C(n_79),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_170),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_168),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_47),
.B1(n_46),
.B2(n_42),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_176),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_46),
.B1(n_42),
.B2(n_43),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_103),
.B(n_43),
.Y(n_174)
);

AND2x4_ASAP7_75t_SL g175 ( 
.A(n_105),
.B(n_122),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_43),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_183),
.Y(n_228)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_106),
.A2(n_18),
.B(n_4),
.C(n_5),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_119),
.B1(n_100),
.B2(n_135),
.Y(n_254)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_111),
.Y(n_185)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_108),
.B(n_18),
.C(n_49),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_133),
.CI(n_148),
.CON(n_233),
.SN(n_233)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_107),
.B(n_49),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_152),
.Y(n_231)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_197),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_215),
.B1(n_135),
.B2(n_145),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_3),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_209),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_134),
.B(n_3),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_146),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_3),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_129),
.A2(n_49),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_217),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_100),
.B1(n_8),
.B2(n_11),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_255),
.B1(n_169),
.B2(n_172),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_231),
.B(n_266),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_218),
.B(n_206),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_166),
.A2(n_145),
.B1(n_144),
.B2(n_132),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_250),
.B1(n_236),
.B2(n_246),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_260),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_173),
.B(n_190),
.CI(n_160),
.CON(n_242),
.SN(n_242)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_242),
.B(n_245),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_164),
.A2(n_124),
.B(n_104),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_175),
.B(n_124),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_246),
.B(n_254),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_136),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_253),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_167),
.A2(n_130),
.B1(n_144),
.B2(n_119),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_136),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_254),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_7),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_191),
.B(n_7),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_219),
.A2(n_211),
.B1(n_213),
.B2(n_196),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_277),
.B1(n_281),
.B2(n_284),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_278),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_220),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_280),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_220),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_219),
.A2(n_161),
.B1(n_218),
.B2(n_201),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_224),
.A2(n_179),
.B1(n_184),
.B2(n_210),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_182),
.B1(n_186),
.B2(n_181),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_293),
.B1(n_299),
.B2(n_303),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_185),
.B(n_217),
.C(n_199),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_316),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_195),
.B1(n_204),
.B2(n_192),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_230),
.B(n_256),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_188),
.B1(n_200),
.B2(n_202),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_295),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_243),
.B(n_202),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_292),
.B(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_228),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_301),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_234),
.A2(n_15),
.B1(n_233),
.B2(n_226),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_15),
.C(n_242),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_221),
.C(n_228),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_233),
.A2(n_15),
.B1(n_254),
.B2(n_269),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_255),
.A2(n_262),
.B1(n_242),
.B2(n_254),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_221),
.B1(n_263),
.B2(n_232),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_269),
.B(n_241),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_252),
.Y(n_327)
);

OAI22x1_ASAP7_75t_SL g308 ( 
.A1(n_254),
.A2(n_262),
.B1(n_263),
.B2(n_251),
.Y(n_308)
);

AOI22x1_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_252),
.B1(n_225),
.B2(n_229),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_240),
.B(n_260),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_310),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_235),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_311),
.B(n_313),
.Y(n_325)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_235),
.B(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_317),
.A2(n_289),
.B1(n_270),
.B2(n_287),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_320),
.B(n_340),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_303),
.A2(n_244),
.B1(n_256),
.B2(n_251),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_333),
.B1(n_344),
.B2(n_345),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_302),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_222),
.C(n_247),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_342),
.C(n_354),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_331),
.B(n_316),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_282),
.A2(n_299),
.B1(n_272),
.B2(n_291),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_247),
.C(n_237),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_298),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_350),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_282),
.A2(n_230),
.B1(n_263),
.B2(n_229),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_304),
.A2(n_225),
.B1(n_237),
.B2(n_257),
.Y(n_345)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_275),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_304),
.A2(n_259),
.B1(n_223),
.B2(n_258),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_290),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_259),
.C(n_258),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_279),
.B(n_223),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_356),
.B(n_357),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_223),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_359),
.B(n_351),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_311),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_360),
.B(n_367),
.C(n_378),
.Y(n_409)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_313),
.C(n_305),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_369),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_343),
.B(n_294),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_372),
.Y(n_400)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_321),
.A2(n_301),
.B1(n_315),
.B2(n_271),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_376),
.A2(n_380),
.B1(n_384),
.B2(n_391),
.Y(n_402)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_302),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_274),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_390),
.C(n_354),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_353),
.A2(n_270),
.B1(n_281),
.B2(n_278),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_310),
.B(n_288),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_381),
.A2(n_388),
.B(n_348),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_295),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_383),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_338),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_321),
.A2(n_293),
.B1(n_308),
.B2(n_310),
.Y(n_384)
);

XNOR2x2_ASAP7_75t_SL g385 ( 
.A(n_336),
.B(n_276),
.Y(n_385)
);

A2O1A1O1Ixp25_ASAP7_75t_L g411 ( 
.A1(n_385),
.A2(n_320),
.B(n_346),
.C(n_351),
.D(n_323),
.Y(n_411)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_388),
.A2(n_331),
.B(n_355),
.Y(n_407)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_350),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_314),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_353),
.A2(n_284),
.B1(n_312),
.B2(n_286),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_345),
.B(n_283),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_324),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_364),
.A2(n_353),
.B1(n_337),
.B2(n_333),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_349),
.B1(n_296),
.B2(n_258),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g395 ( 
.A1(n_381),
.A2(n_329),
.B1(n_337),
.B2(n_348),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_414),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_319),
.B1(n_348),
.B2(n_352),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_399),
.A2(n_405),
.B1(n_412),
.B2(n_418),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_332),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_417),
.C(n_367),
.Y(n_423)
);

XOR2x1_ASAP7_75t_SL g437 ( 
.A(n_404),
.B(n_374),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_364),
.A2(n_319),
.B1(n_344),
.B2(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_406),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g430 ( 
.A1(n_407),
.A2(n_411),
.B(n_371),
.Y(n_430)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_297),
.C(n_334),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_392),
.B1(n_385),
.B2(n_373),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_378),
.C(n_362),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_358),
.A2(n_323),
.B1(n_339),
.B2(n_347),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_339),
.Y(n_419)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_405),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_360),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_441),
.C(n_395),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_403),
.B(n_359),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_429),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_406),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_430),
.A2(n_411),
.B(n_421),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_366),
.C(n_389),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_433),
.C(n_438),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_434),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_387),
.C(n_386),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_407),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_372),
.C(n_363),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_363),
.C(n_334),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_443),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_416),
.B(n_349),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_394),
.B1(n_421),
.B2(n_404),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_456),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_424),
.B(n_409),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_453),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_424),
.B(n_412),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_455),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_414),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_423),
.B(n_397),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_457),
.B(n_463),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_421),
.B(n_399),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_442),
.B1(n_433),
.B2(n_436),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_466),
.C(n_467),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_440),
.B(n_395),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_408),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_465),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_428),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_474),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_451),
.A2(n_445),
.B1(n_427),
.B2(n_434),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_448),
.B1(n_459),
.B2(n_463),
.Y(n_489)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_468),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_478),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_467),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_441),
.C(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_484),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_452),
.B(n_444),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_482),
.Y(n_492)
);

OA21x2_ASAP7_75t_SL g484 ( 
.A1(n_456),
.A2(n_435),
.B(n_415),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_489),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_470),
.A2(n_458),
.B(n_462),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_490),
.B(n_491),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_478),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_449),
.C(n_455),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_493),
.B(n_496),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_453),
.C(n_413),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_420),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_481),
.Y(n_505)
);

BUFx4f_ASAP7_75t_SL g499 ( 
.A(n_492),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_505),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_482),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_502),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_469),
.C(n_471),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_496),
.A2(n_475),
.B1(n_472),
.B2(n_479),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_474),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_506),
.B(n_486),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_511),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_501),
.A2(n_488),
.B(n_493),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_510),
.A2(n_507),
.B(n_509),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_485),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_512),
.B(n_498),
.C(n_490),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_515),
.Y(n_517)
);

AOI31xp33_ASAP7_75t_L g516 ( 
.A1(n_513),
.A2(n_509),
.A3(n_499),
.B(n_498),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_487),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_517),
.B(n_499),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_497),
.B(n_483),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_483),
.C(n_469),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_489),
.B(n_481),
.Y(n_522)
);


endmodule