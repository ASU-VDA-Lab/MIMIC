module fake_jpeg_22174_n_214 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.C(n_2),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_19),
.B1(n_15),
.B2(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_41),
.B1(n_22),
.B2(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_22),
.B1(n_19),
.B2(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_61),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_22),
.C(n_23),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_29),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_73),
.B1(n_21),
.B2(n_17),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_29),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_31),
.C(n_50),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_2),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_40),
.B1(n_32),
.B2(n_34),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_31),
.B1(n_30),
.B2(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_86),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_30),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_91),
.B(n_18),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_36),
.B1(n_20),
.B2(n_16),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_21),
.B(n_18),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_17),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_95),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_105),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_30),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_24),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_109),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_112),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_37),
.B(n_34),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_90),
.B(n_75),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_122),
.B(n_105),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_27),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_82),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_100),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_75),
.B1(n_90),
.B2(n_61),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_99),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_75),
.B1(n_71),
.B2(n_68),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_87),
.C(n_60),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_26),
.B(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_71),
.B1(n_60),
.B2(n_67),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_55),
.B1(n_92),
.B2(n_71),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_87),
.B1(n_99),
.B2(n_89),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_94),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_138),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_140),
.B(n_141),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_106),
.B(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_125),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_146),
.B1(n_116),
.B2(n_119),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_28),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_14),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_120),
.B(n_27),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_127),
.C(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_89),
.B1(n_37),
.B2(n_34),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_161),
.B(n_25),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_159),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_126),
.C(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_59),
.B(n_23),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_156),
.A2(n_132),
.B1(n_124),
.B2(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_145),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_158),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_92),
.B1(n_22),
.B2(n_66),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_175),
.B1(n_162),
.B2(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_66),
.B1(n_53),
.B2(n_52),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_151),
.B1(n_149),
.B2(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_182),
.B1(n_183),
.B2(n_3),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_175),
.B(n_173),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_49),
.B1(n_11),
.B2(n_13),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_49),
.C(n_37),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_34),
.C(n_23),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_170),
.B1(n_166),
.B2(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_28),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_193),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_184),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_194),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g198 ( 
.A1(n_191),
.A2(n_180),
.B(n_13),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_4),
.B(n_5),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_3),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_205),
.C(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_200),
.C(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_4),
.B(n_7),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_180),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_210)
);

AO21x2_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_211),
.B(n_207),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_212),
.A2(n_7),
.B(n_8),
.C(n_28),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_213),
.Y(n_214)
);


endmodule