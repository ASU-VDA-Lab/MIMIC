module fake_jpeg_14622_n_299 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_5),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_6),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_31),
.B(n_30),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_31),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_27),
.B1(n_18),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_32),
.B1(n_33),
.B2(n_17),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_37),
.B1(n_16),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_62),
.B1(n_67),
.B2(n_74),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_63),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_77),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_37),
.B1(n_16),
.B2(n_18),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_56),
.B(n_42),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_37),
.B1(n_32),
.B2(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_72),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_75),
.B1(n_74),
.B2(n_49),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_30),
.B(n_34),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_34),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_91),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_43),
.B1(n_33),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_27),
.B1(n_49),
.B2(n_19),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_88),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_36),
.C(n_35),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_30),
.A3(n_49),
.B1(n_42),
.B2(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_93),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_23),
.B(n_28),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_17),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_0),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_75),
.B(n_78),
.C(n_15),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_42),
.A3(n_14),
.B1(n_24),
.B2(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_14),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_42),
.Y(n_117)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_43),
.B1(n_23),
.B2(n_28),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_75),
.B1(n_15),
.B2(n_21),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_53),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_117),
.B(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_114),
.B1(n_100),
.B2(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_106),
.A2(n_71),
.B1(n_57),
.B2(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_115),
.B1(n_120),
.B2(n_130),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_124),
.B(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_78),
.B1(n_75),
.B2(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_15),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_131),
.Y(n_150)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_21),
.B1(n_22),
.B2(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_26),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_88),
.C(n_101),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_142),
.C(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_103),
.C(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_94),
.B1(n_100),
.B2(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_109),
.B1(n_10),
.B2(n_12),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_81),
.C(n_14),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_20),
.Y(n_148)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_96),
.B1(n_39),
.B2(n_46),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_96),
.B1(n_46),
.B2(n_28),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_24),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_6),
.B(n_9),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_20),
.C(n_29),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_161),
.C(n_26),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_28),
.A3(n_23),
.B1(n_20),
.B2(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_119),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_127),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_8),
.B1(n_11),
.B2(n_9),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_172),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_171),
.B(n_185),
.Y(n_200)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_175),
.B1(n_188),
.B2(n_2),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_128),
.B(n_2),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_181),
.B(n_187),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_1),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_140),
.B(n_136),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_29),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_1),
.Y(n_187)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_86),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_195),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_29),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_158),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_153),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_156),
.C(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_8),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_199),
.C(n_176),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_141),
.B1(n_149),
.B2(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_142),
.C(n_149),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_138),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_168),
.B(n_194),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_206),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_151),
.B1(n_152),
.B2(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_173),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_201),
.B1(n_194),
.B2(n_181),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_174),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_219),
.C(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_193),
.C(n_186),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_177),
.C(n_176),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_225),
.C(n_234),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_177),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_208),
.B(n_203),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_170),
.C(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_187),
.B1(n_179),
.B2(n_170),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_208),
.B1(n_166),
.B2(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_192),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_226),
.B(n_183),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_198),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_246),
.C(n_225),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_210),
.CI(n_204),
.CON(n_242),
.SN(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_249),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_202),
.C(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_215),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_256),
.C(n_263),
.Y(n_264)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_253),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_231),
.B(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_202),
.C(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_211),
.B(n_191),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_262),
.B(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_224),
.C(n_212),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_261),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_272),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_238),
.B1(n_239),
.B2(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_271),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_165),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_244),
.B1(n_236),
.B2(n_241),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_236),
.B(n_242),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_256),
.B(n_263),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_281),
.B(n_237),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_259),
.B1(n_253),
.B2(n_242),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_165),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_258),
.C(n_178),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_287),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_253),
.B(n_260),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_274),
.A3(n_189),
.B1(n_172),
.B2(n_188),
.C1(n_2),
.C2(n_5),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_197),
.B(n_178),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_3),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_286),
.B1(n_289),
.B2(n_283),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_293),
.B(n_288),
.Y(n_296)
);

OAI221xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_4),
.B1(n_5),
.B2(n_29),
.C(n_286),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_4),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_29),
.Y(n_299)
);


endmodule