module fake_jpeg_22617_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_41),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_50),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_19),
.B1(n_30),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_56),
.B1(n_22),
.B2(n_31),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_59),
.B1(n_33),
.B2(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_19),
.B1(n_30),
.B2(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_39),
.B(n_40),
.C(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_81),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_43),
.B1(n_20),
.B2(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_105),
.B1(n_67),
.B2(n_64),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_89),
.B1(n_103),
.B2(n_12),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_29),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_86),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_47),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_45),
.B1(n_41),
.B2(n_26),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_92),
.B1(n_100),
.B2(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_41),
.B1(n_42),
.B2(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_58),
.B1(n_67),
.B2(n_11),
.Y(n_115)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_0),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_42),
.B1(n_44),
.B2(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_44),
.B1(n_26),
.B2(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_17),
.B1(n_26),
.B2(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_130),
.B1(n_87),
.B2(n_75),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_117),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_92),
.B1(n_88),
.B2(n_70),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_10),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_131),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_127),
.B1(n_78),
.B2(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_85),
.Y(n_136)
);

OAI22x1_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_55),
.B1(n_54),
.B2(n_53),
.Y(n_127)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_57),
.B1(n_55),
.B2(n_54),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_57),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_134),
.B(n_136),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_79),
.B(n_81),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_153),
.B(n_155),
.Y(n_175)
);

AO21x1_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_75),
.B(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_107),
.B(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_86),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_96),
.B1(n_100),
.B2(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_101),
.B1(n_97),
.B2(n_99),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_157),
.B1(n_118),
.B2(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_152),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_104),
.B1(n_90),
.B2(n_72),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_151),
.B1(n_158),
.B2(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_162),
.B(n_4),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_102),
.B1(n_98),
.B2(n_78),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_98),
.B1(n_93),
.B2(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_2),
.B(n_3),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_16),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_14),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_116),
.B(n_16),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_16),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_110),
.B1(n_114),
.B2(n_112),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_168),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_114),
.B1(n_119),
.B2(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_197),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_129),
.B1(n_133),
.B2(n_126),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_111),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_5),
.C(n_6),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_121),
.B(n_111),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_179),
.B(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_129),
.B1(n_126),
.B2(n_118),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_111),
.B(n_124),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_189),
.B1(n_163),
.B2(n_147),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_2),
.B(n_3),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_15),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_136),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_2),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_4),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_141),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_14),
.B1(n_13),
.B2(n_9),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_135),
.B1(n_165),
.B2(n_164),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_210),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_182),
.A2(n_152),
.B1(n_149),
.B2(n_162),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_224),
.C(n_172),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_137),
.B(n_141),
.C(n_147),
.Y(n_210)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_137),
.A3(n_141),
.B1(n_14),
.B2(n_13),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_194),
.B1(n_189),
.B2(n_193),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_173),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_229),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_175),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_175),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_176),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_248),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_183),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_236),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_190),
.B1(n_174),
.B2(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_170),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_217),
.B(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_186),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_169),
.B1(n_168),
.B2(n_172),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_187),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_216),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_250),
.B(n_254),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_265),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_238),
.A2(n_220),
.B(n_225),
.Y(n_254)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_260),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_204),
.CI(n_222),
.CON(n_260),
.SN(n_260)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_208),
.B(n_201),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_241),
.B1(n_256),
.B2(n_257),
.Y(n_269)
);

A2O1A1O1Ixp25_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_213),
.B(n_206),
.C(n_210),
.D(n_215),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_210),
.B(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_232),
.C(n_228),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_271),
.C(n_276),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_241),
.B1(n_214),
.B2(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_230),
.C(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_227),
.B1(n_239),
.B2(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_210),
.B1(n_201),
.B2(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_262),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_281),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_236),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_255),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_248),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_199),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_288),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_270),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_294),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_278),
.B1(n_268),
.B2(n_260),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_267),
.B(n_261),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_271),
.C(n_276),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_287),
.C(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_302),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_265),
.B(n_260),
.C(n_270),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_290),
.B1(n_284),
.B2(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_251),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_210),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_286),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.C(n_8),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_8),
.B(n_306),
.Y(n_315)
);

OAI221xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_297),
.B1(n_304),
.B2(n_301),
.C(n_292),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_304),
.B(n_301),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_299),
.A3(n_292),
.B1(n_13),
.B2(n_8),
.C1(n_6),
.C2(n_5),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_315),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_305),
.B(n_317),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_309),
.Y(n_320)
);


endmodule