module fake_aes_5506_n_27 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVxp67_ASAP7_75t_SL g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_15), .B(n_0), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_14), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_17), .Y(n_21) );
NOR3xp33_ASAP7_75t_SL g22 ( .A(n_21), .B(n_18), .C(n_13), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_1), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_5), .B(n_6), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_24), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
OAI221xp5_ASAP7_75t_R g27 ( .A1(n_26), .A2(n_7), .B1(n_9), .B2(n_11), .C(n_12), .Y(n_27) );
endmodule