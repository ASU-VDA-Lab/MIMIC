module real_jpeg_9278_n_18 (n_17, n_8, n_0, n_2, n_10, n_338, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_338;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_1),
.A2(n_23),
.B1(n_61),
.B2(n_62),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_12),
.B(n_33),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_32),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_9),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_90),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_90),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_85),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_85),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_12),
.A2(n_45),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_12),
.B(n_45),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_12),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_12),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_32),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_12),
.B(n_36),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_110),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_13),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_13),
.A2(n_24),
.B1(n_26),
.B2(n_97),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_14),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_126),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_14),
.A2(n_24),
.B1(n_26),
.B2(n_126),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_24),
.B1(n_26),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_15),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_16),
.A2(n_24),
.B1(n_26),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_16),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_17),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_145),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_145),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_17),
.A2(n_24),
.B1(n_26),
.B2(n_145),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_330),
.B(n_333),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_72),
.B(n_329),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_21),
.B(n_37),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_21),
.B(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_21),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_22),
.A2(n_27),
.B1(n_36),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_24),
.A2(n_29),
.B(n_110),
.C(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_27),
.A2(n_36),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_332)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_31),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_28),
.A2(n_31),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_28),
.A2(n_31),
.B1(n_208),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_28),
.A2(n_31),
.B1(n_233),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_28),
.A2(n_31),
.B1(n_251),
.B2(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_28),
.A2(n_31),
.B1(n_52),
.B2(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_65),
.C(n_67),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_38),
.A2(n_39),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.C(n_56),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_304),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_42),
.A2(n_44),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_42),
.A2(n_44),
.B1(n_136),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_42),
.A2(n_44),
.B1(n_153),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_44),
.B1(n_193),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_42),
.A2(n_44),
.B1(n_204),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_42),
.A2(n_44),
.B1(n_230),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_303),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_43),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_44),
.B(n_110),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_45),
.B(n_47),
.Y(n_140)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_46),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_50),
.A2(n_51),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_56),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_56),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_60),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_57),
.A2(n_60),
.B1(n_96),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_60),
.B1(n_123),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_57),
.A2(n_60),
.B1(n_132),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_57),
.A2(n_60),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_57),
.A2(n_60),
.B1(n_216),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_57),
.A2(n_60),
.B1(n_225),
.B2(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_60),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_64),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_65),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_69),
.A2(n_70),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_322),
.B(n_328),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_295),
.A3(n_315),
.B1(n_320),
.B2(n_321),
.C(n_337),
.Y(n_73)
);

AOI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_241),
.A3(n_283),
.B1(n_289),
.B2(n_294),
.C(n_338),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_198),
.C(n_237),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_168),
.B(n_197),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_147),
.B(n_167),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_128),
.B(n_146),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_117),
.B(n_127),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_103),
.B(n_116),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_87),
.B1(n_144),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_107),
.B1(n_108),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_102),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_111),
.B(n_115),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_108),
.B1(n_125),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_107),
.A2(n_108),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_107),
.A2(n_108),
.B1(n_179),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_107),
.A2(n_108),
.B1(n_213),
.B2(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_107),
.A2(n_108),
.B(n_223),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_130),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.CI(n_137),
.CON(n_130),
.SN(n_130)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_160),
.B2(n_161),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_163),
.C(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_170),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_183),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_182),
.C(n_183),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_191),
.C(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_188),
.A2(n_190),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_199),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_218),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_200),
.B(n_218),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_211),
.C(n_217),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_209),
.C(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_217),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_214),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_235),
.B2(n_236),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_226),
.C(n_236),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_224),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_231),
.C(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_260),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_242),
.B(n_260),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.C(n_259),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_243),
.A2(n_244),
.B1(n_253),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_249),
.C(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_253),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_255),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_276),
.B(n_279),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_256),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_281),
.B2(n_282),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_273),
.C(n_282),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_268),
.B(n_271),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_270),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_271),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_271),
.A2(n_297),
.B1(n_306),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_279),
.B2(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_276),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_290),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_286),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_308),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_306),
.C(n_307),
.Y(n_296)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_299),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_304),
.C(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_310),
.C(n_314),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_302),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_327),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule