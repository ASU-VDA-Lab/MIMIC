module real_aes_9359_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_1404;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_0), .A2(n_237), .B1(n_496), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_0), .A2(n_237), .B1(n_490), .B2(n_539), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_1), .A2(n_20), .B1(n_663), .B2(n_750), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_1), .A2(n_254), .B1(n_387), .B2(n_670), .Y(n_1068) );
INVx1_ASAP7_75t_L g1187 ( .A(n_2), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_3), .A2(n_118), .B1(n_394), .B2(n_395), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_118), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g578 ( .A(n_4), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_5), .A2(n_175), .B1(n_666), .B2(n_670), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_5), .A2(n_175), .B1(n_498), .B2(n_696), .Y(n_700) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_6), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_6), .A2(n_45), .B1(n_812), .B2(n_815), .Y(n_811) );
INVx1_ASAP7_75t_L g835 ( .A(n_7), .Y(n_835) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_8), .Y(n_280) );
INVx1_ASAP7_75t_L g408 ( .A(n_8), .Y(n_408) );
INVxp67_ASAP7_75t_SL g900 ( .A(n_9), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_9), .A2(n_25), .B1(n_394), .B2(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g1401 ( .A(n_10), .Y(n_1401) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_11), .A2(n_217), .B1(n_535), .B2(n_536), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_11), .A2(n_217), .B1(n_545), .B2(n_697), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_12), .A2(n_39), .B1(n_416), .B2(n_420), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_12), .A2(n_39), .B1(n_428), .B2(n_430), .Y(n_427) );
AOI221xp5_ASAP7_75t_SL g1096 ( .A1(n_13), .A2(n_37), .B1(n_1097), .B2(n_1098), .C(n_1100), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_13), .A2(n_37), .B1(n_696), .B2(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g317 ( .A(n_14), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_15), .A2(n_213), .B1(n_351), .B2(n_490), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_15), .A2(n_213), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_16), .A2(n_183), .B1(n_535), .B2(n_536), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_16), .A2(n_183), .B1(n_697), .B2(n_929), .Y(n_928) );
AO22x2_ASAP7_75t_L g565 ( .A1(n_17), .A2(n_566), .B1(n_637), .B2(n_638), .Y(n_565) );
INVx1_ASAP7_75t_L g637 ( .A(n_17), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_18), .Y(n_1015) );
INVx1_ASAP7_75t_L g891 ( .A(n_19), .Y(n_891) );
INVx1_ASAP7_75t_L g1055 ( .A(n_20), .Y(n_1055) );
CKINVDCx16_ASAP7_75t_R g1246 ( .A(n_21), .Y(n_1246) );
INVx1_ASAP7_75t_L g756 ( .A(n_22), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_23), .A2(n_259), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_23), .A2(n_259), .B1(n_430), .B2(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_24), .A2(n_210), .B1(n_658), .B2(n_759), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_24), .A2(n_210), .B1(n_1108), .B2(n_1111), .C(n_1113), .Y(n_1107) );
INVx1_ASAP7_75t_L g899 ( .A(n_25), .Y(n_899) );
INVx1_ASAP7_75t_L g939 ( .A(n_26), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_26), .A2(n_130), .B1(n_538), .B2(n_905), .Y(n_965) );
XNOR2xp5_ASAP7_75t_L g1022 ( .A(n_27), .B(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1167 ( .A(n_27), .Y(n_1167) );
AO221x2_ASAP7_75t_L g1177 ( .A1(n_28), .A2(n_60), .B1(n_1148), .B2(n_1156), .C(n_1178), .Y(n_1177) );
INVx2_ASAP7_75t_L g302 ( .A(n_29), .Y(n_302) );
INVx1_ASAP7_75t_L g886 ( .A(n_30), .Y(n_886) );
INVx1_ASAP7_75t_L g1179 ( .A(n_31), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_32), .A2(n_234), .B1(n_535), .B2(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_32), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_33), .A2(n_194), .B1(n_542), .B2(n_722), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g725 ( .A1(n_33), .A2(n_471), .B(n_726), .C(n_729), .Y(n_725) );
BUFx2_ASAP7_75t_L g347 ( .A(n_34), .Y(n_347) );
BUFx2_ASAP7_75t_L g390 ( .A(n_34), .Y(n_390) );
INVx1_ASAP7_75t_L g406 ( .A(n_34), .Y(n_406) );
INVx1_ASAP7_75t_L g1231 ( .A(n_35), .Y(n_1231) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_36), .A2(n_116), .B1(n_545), .B2(n_546), .Y(n_544) );
INVxp67_ASAP7_75t_L g557 ( .A(n_36), .Y(n_557) );
INVx1_ASAP7_75t_L g327 ( .A(n_38), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_38), .A2(n_106), .B1(n_351), .B2(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g337 ( .A(n_40), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_40), .A2(n_144), .B1(n_363), .B2(n_366), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_41), .A2(n_181), .B1(n_351), .B2(n_538), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_41), .A2(n_181), .B1(n_496), .B2(n_503), .Y(n_714) );
INVxp33_ASAP7_75t_L g476 ( .A(n_42), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_42), .A2(n_156), .B1(n_413), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_43), .A2(n_54), .B1(n_394), .B2(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_43), .A2(n_54), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g1066 ( .A(n_44), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_45), .Y(n_790) );
CKINVDCx16_ASAP7_75t_R g1157 ( .A(n_46), .Y(n_1157) );
INVx1_ASAP7_75t_L g1227 ( .A(n_47), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_48), .A2(n_251), .B1(n_351), .B2(n_538), .Y(n_791) );
AOI221xp5_ASAP7_75t_SL g807 ( .A1(n_48), .A2(n_625), .B1(n_808), .B2(n_809), .C(n_817), .Y(n_807) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_49), .A2(n_340), .B(n_752), .C(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g780 ( .A(n_49), .Y(n_780) );
INVx1_ASAP7_75t_L g942 ( .A(n_50), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_50), .A2(n_248), .B1(n_536), .B2(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g890 ( .A(n_51), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_51), .A2(n_205), .B1(n_399), .B2(n_905), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_52), .A2(n_257), .B1(n_498), .B2(n_697), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_52), .A2(n_184), .B1(n_387), .B2(n_670), .Y(n_1018) );
INVx1_ASAP7_75t_L g572 ( .A(n_53), .Y(n_572) );
INVx1_ASAP7_75t_L g868 ( .A(n_55), .Y(n_868) );
OAI211xp5_ASAP7_75t_L g872 ( .A1(n_55), .A2(n_340), .B(n_873), .C(n_875), .Y(n_872) );
XNOR2xp5_ASAP7_75t_L g644 ( .A(n_56), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g1085 ( .A(n_57), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_57), .A2(n_192), .B1(n_1132), .B2(n_1134), .Y(n_1131) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_58), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_59), .A2(n_65), .B1(n_444), .B2(n_1420), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_59), .A2(n_65), .B1(n_1097), .B2(n_1111), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_61), .A2(n_239), .B1(n_503), .B2(n_542), .Y(n_541) );
INVxp33_ASAP7_75t_L g559 ( .A(n_61), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_62), .A2(n_227), .B1(n_351), .B2(n_490), .Y(n_711) );
INVx1_ASAP7_75t_L g736 ( .A(n_62), .Y(n_736) );
INVxp33_ASAP7_75t_L g469 ( .A(n_63), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_63), .A2(n_100), .B1(n_430), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g994 ( .A(n_64), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_64), .A2(n_184), .B1(n_658), .B2(n_663), .Y(n_1010) );
INVx1_ASAP7_75t_L g1241 ( .A(n_66), .Y(n_1241) );
CKINVDCx16_ASAP7_75t_R g1244 ( .A(n_67), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_68), .A2(n_823), .B1(n_877), .B2(n_878), .Y(n_822) );
INVx1_ASAP7_75t_L g878 ( .A(n_68), .Y(n_878) );
INVx1_ASAP7_75t_L g1065 ( .A(n_69), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_70), .A2(n_76), .B1(n_666), .B2(n_670), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_70), .A2(n_76), .B1(n_498), .B2(n_546), .Y(n_846) );
INVx1_ASAP7_75t_L g653 ( .A(n_71), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_72), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_72), .A2(n_129), .B1(n_394), .B2(n_395), .Y(n_687) );
INVx1_ASAP7_75t_L g1036 ( .A(n_73), .Y(n_1036) );
INVx1_ASAP7_75t_L g461 ( .A(n_74), .Y(n_461) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_75), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_75), .A2(n_143), .B1(n_442), .B2(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g1188 ( .A(n_77), .Y(n_1188) );
INVx1_ASAP7_75t_L g957 ( .A(n_78), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_78), .A2(n_89), .B1(n_531), .B2(n_545), .Y(n_971) );
INVx1_ASAP7_75t_L g988 ( .A(n_79), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_79), .A2(n_170), .B1(n_750), .B2(n_759), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_80), .A2(n_151), .B1(n_538), .B2(n_905), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_80), .A2(n_151), .B1(n_496), .B2(n_533), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_81), .A2(n_111), .B1(n_897), .B2(n_947), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_81), .A2(n_111), .B1(n_366), .B2(n_463), .Y(n_952) );
INVx1_ASAP7_75t_L g909 ( .A(n_82), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_82), .A2(n_105), .B1(n_531), .B2(n_545), .Y(n_933) );
INVx1_ASAP7_75t_L g1041 ( .A(n_83), .Y(n_1041) );
OAI211xp5_ASAP7_75t_SL g1069 ( .A1(n_83), .A2(n_471), .B(n_673), .C(n_1070), .Y(n_1069) );
AO22x2_ASAP7_75t_L g452 ( .A1(n_84), .A2(n_453), .B1(n_506), .B2(n_507), .Y(n_452) );
INVx1_ASAP7_75t_L g506 ( .A(n_84), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_85), .Y(n_1081) );
INVxp33_ASAP7_75t_SL g1408 ( .A(n_86), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_86), .A2(n_250), .B1(n_539), .B2(n_1116), .Y(n_1434) );
INVxp33_ASAP7_75t_SL g310 ( .A(n_87), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_87), .A2(n_166), .B1(n_394), .B2(n_395), .Y(n_393) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_88), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_88), .A2(n_208), .B1(n_601), .B2(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g955 ( .A(n_89), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_90), .A2(n_192), .B1(n_666), .B2(n_670), .Y(n_1078) );
INVx1_ASAP7_75t_L g1130 ( .A(n_90), .Y(n_1130) );
INVx1_ASAP7_75t_L g521 ( .A(n_91), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_91), .A2(n_98), .B1(n_363), .B2(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g744 ( .A(n_92), .Y(n_744) );
INVxp33_ASAP7_75t_SL g587 ( .A(n_93), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_93), .A2(n_198), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g345 ( .A(n_94), .Y(n_345) );
INVx1_ASAP7_75t_L g575 ( .A(n_95), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_95), .A2(n_190), .B1(n_606), .B2(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g731 ( .A(n_96), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_97), .A2(n_202), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_97), .A2(n_202), .B1(n_620), .B2(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g522 ( .A(n_98), .Y(n_522) );
INVx1_ASAP7_75t_L g836 ( .A(n_99), .Y(n_836) );
INVx1_ASAP7_75t_L g459 ( .A(n_100), .Y(n_459) );
INVx1_ASAP7_75t_L g1007 ( .A(n_101), .Y(n_1007) );
OAI211xp5_ASAP7_75t_SL g1019 ( .A1(n_101), .A2(n_471), .B(n_673), .C(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_102), .A2(n_163), .B1(n_1422), .B2(n_1425), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_102), .A2(n_163), .B1(n_1108), .B2(n_1399), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_103), .A2(n_196), .B1(n_896), .B2(n_897), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_103), .A2(n_196), .B1(n_363), .B2(n_366), .Y(n_906) );
INVx1_ASAP7_75t_L g1030 ( .A(n_104), .Y(n_1030) );
INVxp67_ASAP7_75t_L g911 ( .A(n_105), .Y(n_911) );
INVxp33_ASAP7_75t_SL g298 ( .A(n_106), .Y(n_298) );
INVx1_ASAP7_75t_L g1058 ( .A(n_107), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_108), .A2(n_139), .B1(n_434), .B2(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_108), .A2(n_139), .B1(n_666), .B2(n_670), .Y(n_724) );
INVx1_ASAP7_75t_L g866 ( .A(n_109), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_109), .A2(n_149), .B1(n_658), .B2(n_759), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_110), .A2(n_135), .B1(n_1171), .B2(n_1174), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g985 ( .A(n_112), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_112), .A2(n_195), .B1(n_697), .B2(n_720), .Y(n_1000) );
INVx1_ASAP7_75t_L g1164 ( .A(n_113), .Y(n_1164) );
INVxp33_ASAP7_75t_SL g1395 ( .A(n_114), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_114), .A2(n_249), .B1(n_1420), .B2(n_1428), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_115), .A2(n_150), .B1(n_444), .B2(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_115), .Y(n_851) );
INVxp33_ASAP7_75t_L g556 ( .A(n_116), .Y(n_556) );
AO221x2_ASAP7_75t_L g1184 ( .A1(n_117), .A2(n_180), .B1(n_1156), .B2(n_1185), .C(n_1186), .Y(n_1184) );
OAI211xp5_ASAP7_75t_L g762 ( .A1(n_119), .A2(n_471), .B(n_763), .C(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g803 ( .A(n_119), .Y(n_803) );
INVx1_ASAP7_75t_L g1040 ( .A(n_120), .Y(n_1040) );
OAI22xp33_ASAP7_75t_SL g1071 ( .A1(n_120), .A2(n_147), .B1(n_281), .B2(n_666), .Y(n_1071) );
AO22x2_ASAP7_75t_L g511 ( .A1(n_121), .A2(n_512), .B1(n_561), .B2(n_562), .Y(n_511) );
INVx1_ASAP7_75t_L g561 ( .A(n_121), .Y(n_561) );
INVx1_ASAP7_75t_L g272 ( .A(n_122), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_123), .A2(n_182), .B1(n_658), .B2(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g771 ( .A(n_123), .Y(n_771) );
INVx1_ASAP7_75t_L g954 ( .A(n_124), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_124), .A2(n_212), .B1(n_533), .B2(n_932), .Y(n_970) );
OAI211xp5_ASAP7_75t_L g826 ( .A1(n_125), .A2(n_471), .B(n_827), .C(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g845 ( .A(n_125), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_126), .A2(n_194), .B1(n_281), .B2(n_387), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_126), .A2(n_227), .B1(n_658), .B2(n_663), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_127), .A2(n_172), .B1(n_1148), .B2(n_1156), .Y(n_1176) );
INVx1_ASAP7_75t_L g524 ( .A(n_128), .Y(n_524) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_129), .Y(n_655) );
INVx1_ASAP7_75t_L g945 ( .A(n_130), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_131), .A2(n_134), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_131), .A2(n_134), .B1(n_535), .B2(n_536), .Y(n_547) );
INVx1_ASAP7_75t_L g1180 ( .A(n_132), .Y(n_1180) );
XOR2xp5_ASAP7_75t_L g973 ( .A(n_133), .B(n_974), .Y(n_973) );
INVxp33_ASAP7_75t_SL g515 ( .A(n_136), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_136), .A2(n_153), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g470 ( .A(n_137), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_138), .A2(n_146), .B1(n_535), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_138), .A2(n_146), .B1(n_498), .B2(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_140), .A2(n_191), .B1(n_658), .B2(n_663), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_140), .A2(n_226), .B1(n_420), .B2(n_689), .Y(n_688) );
INVxp33_ASAP7_75t_L g457 ( .A(n_141), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_141), .A2(n_155), .B1(n_434), .B2(n_498), .Y(n_505) );
INVx1_ASAP7_75t_L g1033 ( .A(n_142), .Y(n_1033) );
INVxp33_ASAP7_75t_L g377 ( .A(n_143), .Y(n_377) );
INVx1_ASAP7_75t_L g332 ( .A(n_144), .Y(n_332) );
INVx1_ASAP7_75t_L g464 ( .A(n_145), .Y(n_464) );
INVx1_ASAP7_75t_L g1044 ( .A(n_147), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1082 ( .A(n_148), .Y(n_1082) );
INVx1_ASAP7_75t_L g859 ( .A(n_149), .Y(n_859) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_150), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_152), .A2(n_161), .B1(n_1171), .B2(n_1174), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_153), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_154), .Y(n_1101) );
INVxp33_ASAP7_75t_L g456 ( .A(n_155), .Y(n_456) );
INVxp33_ASAP7_75t_L g478 ( .A(n_156), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_157), .A2(n_229), .B1(n_351), .B2(n_399), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_157), .A2(n_229), .B1(n_495), .B2(n_496), .Y(n_494) );
INVxp33_ASAP7_75t_SL g525 ( .A(n_158), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_158), .A2(n_176), .B1(n_535), .B2(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g981 ( .A(n_159), .Y(n_981) );
INVx1_ASAP7_75t_L g1054 ( .A(n_160), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_160), .A2(n_174), .B1(n_658), .B2(n_759), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_162), .A2(n_215), .B1(n_1185), .B2(n_1195), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_164), .Y(n_274) );
AND3x2_ASAP7_75t_L g1149 ( .A(n_164), .B(n_272), .C(n_1150), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_164), .B(n_272), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_165), .A2(n_228), .B1(n_663), .B2(n_750), .Y(n_749) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_165), .A2(n_199), .B1(n_281), .B2(n_387), .Y(n_767) );
INVxp33_ASAP7_75t_SL g321 ( .A(n_166), .Y(n_321) );
INVxp33_ASAP7_75t_SL g384 ( .A(n_167), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_167), .A2(n_233), .B1(n_428), .B2(n_430), .Y(n_440) );
INVxp33_ASAP7_75t_L g479 ( .A(n_168), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_168), .A2(n_173), .B1(n_351), .B2(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g652 ( .A(n_169), .Y(n_652) );
INVx1_ASAP7_75t_L g991 ( .A(n_170), .Y(n_991) );
INVx2_ASAP7_75t_L g285 ( .A(n_171), .Y(n_285) );
INVx1_ASAP7_75t_L g474 ( .A(n_173), .Y(n_474) );
INVx1_ASAP7_75t_L g1057 ( .A(n_174), .Y(n_1057) );
INVxp33_ASAP7_75t_SL g516 ( .A(n_176), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1212 ( .A1(n_177), .A2(n_186), .B1(n_1148), .B2(n_1156), .Y(n_1212) );
INVx1_ASAP7_75t_L g830 ( .A(n_178), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_179), .A2(n_204), .B1(n_487), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_179), .A2(n_204), .B1(n_498), .B2(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g778 ( .A(n_182), .Y(n_778) );
INVx1_ASAP7_75t_L g1150 ( .A(n_185), .Y(n_1150) );
CKINVDCx16_ASAP7_75t_R g1154 ( .A(n_187), .Y(n_1154) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_188), .A2(n_471), .B(n_673), .C(n_677), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_188), .A2(n_264), .B1(n_533), .B2(n_693), .Y(n_699) );
INVx1_ASAP7_75t_L g1229 ( .A(n_189), .Y(n_1229) );
INVxp33_ASAP7_75t_SL g569 ( .A(n_190), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_191), .A2(n_264), .B1(n_281), .B2(n_387), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_193), .A2(n_258), .B1(n_666), .B2(n_670), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_193), .A2(n_258), .B1(n_433), .B2(n_805), .Y(n_804) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_195), .Y(n_983) );
INVx1_ASAP7_75t_L g978 ( .A(n_197), .Y(n_978) );
INVxp33_ASAP7_75t_SL g588 ( .A(n_198), .Y(n_588) );
INVx1_ASAP7_75t_L g799 ( .A(n_199), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_200), .A2(n_265), .B1(n_281), .B2(n_387), .Y(n_825) );
INVx1_ASAP7_75t_L g842 ( .A(n_200), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_201), .Y(n_940) );
INVx1_ASAP7_75t_L g287 ( .A(n_203), .Y(n_287) );
INVx2_ASAP7_75t_L g361 ( .A(n_203), .Y(n_361) );
INVx1_ASAP7_75t_L g894 ( .A(n_205), .Y(n_894) );
INVx1_ASAP7_75t_L g903 ( .A(n_206), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_206), .A2(n_256), .B1(n_692), .B2(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_207), .A2(n_240), .B1(n_399), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_207), .A2(n_240), .B1(n_925), .B2(n_926), .Y(n_924) );
INVxp33_ASAP7_75t_SL g570 ( .A(n_208), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g935 ( .A(n_209), .B(n_936), .Y(n_935) );
INVxp67_ASAP7_75t_SL g1415 ( .A(n_211), .Y(n_1415) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_211), .A2(n_252), .B1(n_1108), .B2(n_1111), .Y(n_1433) );
INVx1_ASAP7_75t_L g950 ( .A(n_212), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_214), .A2(n_242), .B1(n_1171), .B2(n_1174), .Y(n_1211) );
XOR2xp5_ASAP7_75t_L g1442 ( .A(n_216), .B(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g995 ( .A(n_218), .Y(n_995) );
OAI211xp5_ASAP7_75t_L g1089 ( .A1(n_219), .A2(n_340), .B(n_800), .C(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1117 ( .A(n_219), .Y(n_1117) );
INVx1_ASAP7_75t_L g757 ( .A(n_220), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_221), .A2(n_747), .B1(n_819), .B2(n_820), .Y(n_746) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_221), .Y(n_820) );
INVx1_ASAP7_75t_L g1404 ( .A(n_222), .Y(n_1404) );
INVx1_ASAP7_75t_L g1004 ( .A(n_223), .Y(n_1004) );
OAI22xp33_ASAP7_75t_SL g1021 ( .A1(n_223), .A2(n_257), .B1(n_281), .B2(n_666), .Y(n_1021) );
INVx1_ASAP7_75t_L g1398 ( .A(n_224), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_224), .A2(n_245), .B1(n_444), .B2(n_1411), .Y(n_1426) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_225), .Y(n_1083) );
INVx1_ASAP7_75t_L g649 ( .A(n_226), .Y(n_649) );
INVx1_ASAP7_75t_L g775 ( .A(n_228), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_230), .A2(n_246), .B1(n_663), .B2(n_750), .Y(n_1092) );
INVx1_ASAP7_75t_L g1114 ( .A(n_230), .Y(n_1114) );
INVx1_ASAP7_75t_L g829 ( .A(n_231), .Y(n_829) );
INVx1_ASAP7_75t_L g1242 ( .A(n_232), .Y(n_1242) );
AO22x2_ASAP7_75t_L g1391 ( .A1(n_232), .A2(n_1242), .B1(n_1392), .B2(n_1435), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1440 ( .A1(n_232), .A2(n_1441), .B1(n_1445), .B2(n_1447), .Y(n_1440) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_233), .Y(n_356) );
INVx1_ASAP7_75t_L g742 ( .A(n_234), .Y(n_742) );
INVx1_ASAP7_75t_L g1153 ( .A(n_235), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_235), .B(n_1163), .Y(n_1166) );
XOR2x2_ASAP7_75t_L g294 ( .A(n_236), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g581 ( .A(n_238), .Y(n_581) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_239), .Y(n_551) );
INVx1_ASAP7_75t_L g1028 ( .A(n_241), .Y(n_1028) );
INVx1_ASAP7_75t_L g730 ( .A(n_243), .Y(n_730) );
AO22x2_ASAP7_75t_L g1074 ( .A1(n_244), .A2(n_1075), .B1(n_1076), .B2(n_1136), .Y(n_1074) );
INVxp67_ASAP7_75t_L g1136 ( .A(n_244), .Y(n_1136) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_245), .Y(n_1396) );
INVx1_ASAP7_75t_L g1086 ( .A(n_246), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_247), .Y(n_1014) );
INVx1_ASAP7_75t_L g943 ( .A(n_248), .Y(n_943) );
INVxp33_ASAP7_75t_SL g1403 ( .A(n_249), .Y(n_1403) );
INVx1_ASAP7_75t_L g1410 ( .A(n_250), .Y(n_1410) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_251), .Y(n_810) );
INVxp33_ASAP7_75t_SL g1413 ( .A(n_252), .Y(n_1413) );
INVx2_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
INVx1_ASAP7_75t_L g1045 ( .A(n_254), .Y(n_1045) );
INVxp33_ASAP7_75t_SL g597 ( .A(n_255), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_255), .A2(n_266), .B1(n_629), .B2(n_631), .Y(n_628) );
INVxp33_ASAP7_75t_L g908 ( .A(n_256), .Y(n_908) );
INVx1_ASAP7_75t_L g861 ( .A(n_260), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_260), .A2(n_265), .B1(n_663), .B2(n_750), .Y(n_876) );
BUFx3_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
INVx1_ASAP7_75t_L g325 ( .A(n_261), .Y(n_325) );
BUFx3_ASAP7_75t_L g309 ( .A(n_262), .Y(n_309) );
INVx1_ASAP7_75t_L g315 ( .A(n_262), .Y(n_315) );
INVx1_ASAP7_75t_L g1400 ( .A(n_263), .Y(n_1400) );
INVx1_ASAP7_75t_L g593 ( .A(n_266), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_288), .B(n_1139), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_270), .B(n_276), .Y(n_1439) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1446 ( .A(n_271), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_271), .B(n_273), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_273), .B(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g389 ( .A(n_278), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g560 ( .A(n_278), .B(n_390), .Y(n_560) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g425 ( .A(n_279), .B(n_287), .Y(n_425) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g793 ( .A(n_280), .B(n_372), .Y(n_793) );
INVx8_ASAP7_75t_L g385 ( .A(n_281), .Y(n_385) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
OR2x6_ASAP7_75t_L g387 ( .A(n_282), .B(n_371), .Y(n_387) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_282), .Y(n_779) );
INVx1_ASAP7_75t_L g865 ( .A(n_282), .Y(n_865) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_282), .Y(n_993) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_282), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1103 ( .A(n_282), .Y(n_1103) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g354 ( .A(n_284), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_284), .Y(n_368) );
INVx2_ASAP7_75t_L g374 ( .A(n_284), .Y(n_374) );
AND2x4_ASAP7_75t_L g381 ( .A(n_284), .B(n_355), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_284), .B(n_285), .Y(n_402) );
INVx2_ASAP7_75t_L g355 ( .A(n_285), .Y(n_355) );
INVx1_ASAP7_75t_L g365 ( .A(n_285), .Y(n_365) );
INVx1_ASAP7_75t_L g376 ( .A(n_285), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_285), .B(n_374), .Y(n_669) );
INVx1_ASAP7_75t_L g676 ( .A(n_285), .Y(n_676) );
AND2x4_ASAP7_75t_L g364 ( .A(n_286), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g366 ( .A(n_287), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g554 ( .A(n_287), .B(n_367), .Y(n_554) );
XOR2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_640), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_509), .B2(n_510), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_451), .B1(n_452), .B2(n_508), .Y(n_293) );
INVx1_ASAP7_75t_L g508 ( .A(n_294), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_343), .B1(n_348), .B2(n_388), .C(n_391), .Y(n_295) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_297), .B(n_316), .C(n_326), .D(n_340), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_310), .B2(n_311), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_299), .A2(n_311), .B1(n_515), .B2(n_516), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_299), .A2(n_311), .B1(n_569), .B2(n_570), .Y(n_568) );
AOI22xp5_ASAP7_75t_SL g889 ( .A1(n_299), .A2(n_318), .B1(n_890), .B2(n_891), .Y(n_889) );
HB1xp67_ASAP7_75t_L g1414 ( .A(n_299), .Y(n_1414) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
AND2x6_ASAP7_75t_L g322 ( .A(n_300), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g480 ( .A(n_300), .B(n_303), .Y(n_480) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g738 ( .A(n_301), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g313 ( .A(n_302), .Y(n_313) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
AND2x2_ASAP7_75t_L g438 ( .A(n_302), .B(n_345), .Y(n_438) );
INVx2_ASAP7_75t_L g450 ( .A(n_302), .Y(n_450) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_304), .Y(n_429) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_304), .Y(n_630) );
INVx1_ASAP7_75t_L g722 ( .A(n_304), .Y(n_722) );
INVx1_ASAP7_75t_L g925 ( .A(n_304), .Y(n_925) );
INVx2_ASAP7_75t_L g1133 ( .A(n_304), .Y(n_1133) );
INVx2_ASAP7_75t_L g1424 ( .A(n_304), .Y(n_1424) );
INVx6_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g318 ( .A(n_305), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g504 ( .A(n_305), .Y(n_504) );
BUFx2_ASAP7_75t_L g692 ( .A(n_305), .Y(n_692) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g314 ( .A(n_307), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g331 ( .A(n_307), .B(n_309), .Y(n_331) );
INVx1_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g324 ( .A(n_309), .B(n_325), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_311), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_311), .A2(n_322), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_311), .A2(n_322), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx6p67_ASAP7_75t_R g759 ( .A(n_311), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_311), .A2(n_322), .B1(n_899), .B2(n_900), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_311), .A2(n_322), .B1(n_942), .B2(n_943), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_311), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
AND2x6_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
INVx1_ASAP7_75t_L g659 ( .A(n_312), .Y(n_659) );
AND2x2_ASAP7_75t_L g893 ( .A(n_312), .B(n_496), .Y(n_893) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x6_ASAP7_75t_L g338 ( .A(n_313), .B(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g433 ( .A(n_314), .Y(n_433) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_314), .Y(n_443) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_314), .Y(n_498) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_314), .Y(n_530) );
BUFx3_ASAP7_75t_L g545 ( .A(n_314), .Y(n_545) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_314), .Y(n_633) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_314), .Y(n_720) );
INVx2_ASAP7_75t_SL g839 ( .A(n_314), .Y(n_839) );
INVx1_ASAP7_75t_L g662 ( .A(n_315), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_321), .B2(n_322), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_317), .A2(n_384), .B1(n_385), .B2(n_386), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_318), .A2(n_322), .B1(n_341), .B2(n_470), .C(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_318), .A2(n_322), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_318), .A2(n_322), .B1(n_572), .B2(n_573), .Y(n_571) );
INVx4_ASAP7_75t_L g663 ( .A(n_318), .Y(n_663) );
AOI22xp5_ASAP7_75t_SL g938 ( .A1(n_318), .A2(n_480), .B1(n_939), .B2(n_940), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_318), .A2(n_322), .B1(n_1404), .B2(n_1408), .Y(n_1407) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_319), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g580 ( .A(n_319), .B(n_334), .Y(n_580) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g750 ( .A(n_322), .Y(n_750) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_323), .Y(n_434) );
INVx1_ASAP7_75t_L g500 ( .A(n_323), .Y(n_500) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_323), .Y(n_531) );
INVx2_ASAP7_75t_L g623 ( .A(n_323), .Y(n_623) );
INVx1_ASAP7_75t_L g806 ( .A(n_323), .Y(n_806) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g447 ( .A(n_324), .Y(n_447) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_324), .Y(n_697) );
INVx1_ASAP7_75t_L g717 ( .A(n_324), .Y(n_717) );
INVx1_ASAP7_75t_L g661 ( .A(n_325), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_332), .B2(n_333), .C1(n_337), .C2(n_338), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g473 ( .A1(n_328), .A2(n_333), .B1(n_338), .B2(n_461), .C1(n_464), .C2(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g341 ( .A(n_330), .B(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_330), .Y(n_496) );
INVx2_ASAP7_75t_L g543 ( .A(n_330), .Y(n_543) );
INVx1_ASAP7_75t_L g927 ( .A(n_330), .Y(n_927) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_331), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g517 ( .A1(n_333), .A2(n_338), .B1(n_518), .B2(n_519), .C1(n_521), .C2(n_522), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g648 ( .A1(n_333), .A2(n_338), .B1(n_649), .B2(n_650), .C1(n_652), .C2(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g739 ( .A(n_335), .Y(n_739) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g814 ( .A(n_336), .Y(n_814) );
AOI222xp33_ASAP7_75t_L g574 ( .A1(n_338), .A2(n_575), .B1(n_576), .B2(n_578), .C1(n_579), .C2(n_581), .Y(n_574) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_338), .A2(n_730), .B1(n_731), .B2(n_736), .C1(n_737), .C2(n_738), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_338), .A2(n_580), .B1(n_756), .B2(n_757), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_338), .A2(n_580), .B1(n_829), .B2(n_830), .Y(n_875) );
INVx3_ASAP7_75t_L g897 ( .A(n_338), .Y(n_897) );
AOI222xp33_ASAP7_75t_L g1012 ( .A1(n_338), .A2(n_738), .B1(n_995), .B2(n_1013), .C1(n_1014), .C2(n_1015), .Y(n_1012) );
AOI222xp33_ASAP7_75t_L g1063 ( .A1(n_338), .A2(n_738), .B1(n_1058), .B2(n_1064), .C1(n_1065), .C2(n_1066), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_338), .A2(n_579), .B1(n_1081), .B2(n_1083), .Y(n_1090) );
AOI222xp33_ASAP7_75t_L g1409 ( .A1(n_338), .A2(n_579), .B1(n_1400), .B2(n_1401), .C1(n_1410), .C2(n_1411), .Y(n_1409) );
BUFx3_ASAP7_75t_L g816 ( .A(n_339), .Y(n_816) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_340), .B(n_514), .C(n_517), .D(n_523), .Y(n_513) );
NAND3xp33_ASAP7_75t_SL g647 ( .A(n_340), .B(n_648), .C(n_654), .Y(n_647) );
NAND3xp33_ASAP7_75t_SL g734 ( .A(n_340), .B(n_735), .C(n_740), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g1011 ( .A(n_340), .B(n_1012), .Y(n_1011) );
NAND2xp5_ASAP7_75t_SL g1062 ( .A(n_340), .B(n_1063), .Y(n_1062) );
CKINVDCx8_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
INVx5_ASAP7_75t_L g583 ( .A(n_341), .Y(n_583) );
AOI221x1_ASAP7_75t_L g453 ( .A1(n_343), .A2(n_388), .B1(n_454), .B2(n_472), .C(n_481), .Y(n_453) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_343), .Y(n_584) );
AOI221x1_ASAP7_75t_L g1392 ( .A1(n_343), .A2(n_388), .B1(n_1393), .B2(n_1406), .C(n_1416), .Y(n_1392) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AND2x4_ASAP7_75t_L g526 ( .A(n_344), .B(n_346), .Y(n_526) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g449 ( .A(n_345), .B(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
OR2x6_ASAP7_75t_L g792 ( .A(n_347), .B(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_369), .C(n_383), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_356), .B(n_357), .C(n_362), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g357 ( .A(n_353), .B(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_353), .Y(n_422) );
BUFx2_ASAP7_75t_L g460 ( .A(n_353), .Y(n_460) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_353), .Y(n_539) );
BUFx3_ASAP7_75t_L g905 ( .A(n_353), .Y(n_905) );
INVx1_ASAP7_75t_L g917 ( .A(n_353), .Y(n_917) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
CKINVDCx11_ASAP7_75t_R g471 ( .A(n_357), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_357), .A2(n_551), .B(n_552), .C(n_553), .Y(n_550) );
AOI211xp5_ASAP7_75t_L g902 ( .A1(n_357), .A2(n_903), .B(n_904), .C(n_906), .Y(n_902) );
AOI211xp5_ASAP7_75t_L g949 ( .A1(n_357), .A2(n_950), .B(n_951), .C(n_952), .Y(n_949) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g467 ( .A(n_359), .Y(n_467) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_360), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_361), .Y(n_372) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g463 ( .A(n_364), .Y(n_463) );
INVx2_ASAP7_75t_L g591 ( .A(n_364), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_364), .A2(n_592), .B1(n_730), .B2(n_731), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_364), .A2(n_592), .B1(n_1014), .B2(n_1015), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_364), .A2(n_592), .B1(n_1065), .B2(n_1066), .Y(n_1070) );
AOI222xp33_ASAP7_75t_L g1080 ( .A1(n_364), .A2(n_539), .B1(n_592), .B2(n_1081), .C1(n_1082), .C2(n_1083), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g1397 ( .A1(n_364), .A2(n_592), .B1(n_1398), .B2(n_1399), .C1(n_1400), .C2(n_1401), .Y(n_1397) );
INVx1_ASAP7_75t_L g466 ( .A(n_367), .Y(n_466) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g675 ( .A(n_368), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_368), .B(n_676), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_377), .B1(n_378), .B2(n_382), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_370), .A2(n_378), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_370), .A2(n_378), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_370), .A2(n_378), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_370), .A2(n_385), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_370), .A2(n_385), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_370), .A2(n_671), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x4_ASAP7_75t_L g378 ( .A(n_371), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g667 ( .A(n_371), .Y(n_667) );
AND2x4_ASAP7_75t_L g671 ( .A(n_371), .B(n_379), .Y(n_671) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
INVx1_ASAP7_75t_L g488 ( .A(n_373), .Y(n_488) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_373), .Y(n_535) );
BUFx2_ASAP7_75t_L g601 ( .A(n_373), .Y(n_601) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_373), .Y(n_964) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_373), .Y(n_1099) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_380), .Y(n_921) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_381), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_385), .A2(n_386), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_385), .A2(n_386), .B1(n_524), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_385), .A2(n_386), .B1(n_572), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_385), .A2(n_386), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_385), .A2(n_1403), .B1(n_1404), .B2(n_1405), .Y(n_1402) );
AOI22xp33_ASAP7_75t_SL g910 ( .A1(n_386), .A2(n_671), .B1(n_891), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_386), .A2(n_671), .B1(n_940), .B2(n_957), .Y(n_956) );
INVx5_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx4_ASAP7_75t_L g1405 ( .A(n_387), .Y(n_1405) );
AOI221x1_ASAP7_75t_L g566 ( .A1(n_388), .A2(n_567), .B1(n_584), .B2(n_585), .C(n_598), .Y(n_566) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_388), .A2(n_665), .A3(n_672), .B(n_678), .Y(n_664) );
OAI31xp33_ASAP7_75t_SL g723 ( .A1(n_388), .A2(n_724), .A3(n_725), .B(n_732), .Y(n_723) );
OAI31xp33_ASAP7_75t_L g760 ( .A1(n_388), .A2(n_761), .A3(n_762), .B(n_767), .Y(n_760) );
OAI31xp33_ASAP7_75t_L g824 ( .A1(n_388), .A2(n_825), .A3(n_826), .B(n_831), .Y(n_824) );
OAI31xp33_ASAP7_75t_SL g1017 ( .A1(n_388), .A2(n_1018), .A3(n_1019), .B(n_1021), .Y(n_1017) );
OAI31xp33_ASAP7_75t_SL g1067 ( .A1(n_388), .A2(n_1068), .A3(n_1069), .B(n_1071), .Y(n_1067) );
O2A1O1Ixp33_ASAP7_75t_L g1077 ( .A1(n_388), .A2(n_1078), .B(n_1079), .C(n_1087), .Y(n_1077) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g448 ( .A(n_390), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g636 ( .A(n_390), .B(n_449), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g391 ( .A(n_392), .B(n_409), .C(n_426), .D(n_439), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_398), .C(n_403), .Y(n_392) );
INVx1_ASAP7_75t_L g862 ( .A(n_395), .Y(n_862) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g706 ( .A(n_396), .Y(n_706) );
INVx2_ASAP7_75t_L g710 ( .A(n_396), .Y(n_710) );
INVx2_ASAP7_75t_L g789 ( .A(n_396), .Y(n_789) );
INVx3_ASAP7_75t_L g857 ( .A(n_396), .Y(n_857) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g684 ( .A(n_397), .Y(n_684) );
INVx3_ASAP7_75t_L g990 ( .A(n_397), .Y(n_990) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g490 ( .A(n_400), .Y(n_490) );
INVx2_ASAP7_75t_L g538 ( .A(n_400), .Y(n_538) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g689 ( .A(n_401), .Y(n_689) );
BUFx6f_ASAP7_75t_L g1110 ( .A(n_401), .Y(n_1110) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g419 ( .A(n_402), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_403), .B(n_610), .C(n_613), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_403), .B(n_687), .C(n_688), .Y(n_686) );
CKINVDCx8_ASAP7_75t_R g1121 ( .A(n_403), .Y(n_1121) );
INVx5_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx6_ASAP7_75t_L g712 ( .A(n_404), .Y(n_712) );
OR2x6_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g492 ( .A(n_407), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_415), .C(n_423), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g615 ( .A(n_418), .Y(n_615) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g605 ( .A(n_419), .Y(n_605) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g951 ( .A(n_421), .Y(n_951) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_423), .B(n_483), .C(n_484), .Y(n_482) );
AOI33xp33_ASAP7_75t_L g540 ( .A1(n_423), .A2(n_448), .A3(n_541), .B1(n_544), .B2(n_547), .B3(n_548), .Y(n_540) );
INVx2_ASAP7_75t_L g608 ( .A(n_423), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_423), .B(n_681), .C(n_685), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_423), .B(n_705), .C(n_707), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g913 ( .A(n_423), .B(n_914), .C(n_915), .Y(n_913) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_423), .B(n_960), .C(n_961), .Y(n_959) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OR2x2_ASAP7_75t_L g436 ( .A(n_424), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g491 ( .A(n_424), .B(n_492), .Y(n_491) );
OR2x6_ASAP7_75t_L g625 ( .A(n_424), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_424), .B(n_626), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .C(n_435), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
INVx4_ASAP7_75t_L g618 ( .A(n_429), .Y(n_618) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_430), .Y(n_1411) );
BUFx4f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g520 ( .A(n_431), .Y(n_520) );
BUFx3_ASAP7_75t_L g631 ( .A(n_431), .Y(n_631) );
INVx1_ASAP7_75t_L g651 ( .A(n_431), .Y(n_651) );
INVx2_ASAP7_75t_SL g694 ( .A(n_431), .Y(n_694) );
BUFx6f_ASAP7_75t_L g932 ( .A(n_431), .Y(n_932) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_435), .B(n_494), .C(n_497), .Y(n_493) );
AOI33xp33_ASAP7_75t_L g528 ( .A1(n_435), .A2(n_491), .A3(n_529), .B1(n_532), .B2(n_534), .B3(n_537), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_435), .B(n_691), .C(n_695), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_435), .B(n_714), .C(n_715), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_435), .B(n_924), .C(n_928), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_435), .B(n_967), .C(n_968), .Y(n_966) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g997 ( .A1(n_436), .A2(n_998), .B1(n_1001), .B2(n_1002), .Y(n_997) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g626 ( .A(n_438), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .C(n_448), .Y(n_439) );
BUFx4f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g1029 ( .A(n_443), .Y(n_1029) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g546 ( .A(n_446), .Y(n_546) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_448), .B(n_502), .C(n_505), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_448), .B(n_699), .C(n_700), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_448), .B(n_719), .C(n_721), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_448), .B(n_931), .C(n_933), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_448), .B(n_970), .C(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g1046 ( .A(n_448), .Y(n_1046) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g507 ( .A(n_453), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .C(n_468), .D(n_471), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_461), .B2(n_462), .C1(n_464), .C2(n_465), .Y(n_458) );
INVx1_ASAP7_75t_L g595 ( .A(n_460), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_462), .A2(n_592), .B1(n_652), .B2(n_653), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_462), .A2(n_592), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x4_ASAP7_75t_L g592 ( .A(n_466), .B(n_467), .Y(n_592) );
NAND4xp25_ASAP7_75t_SL g585 ( .A(n_471), .B(n_586), .C(n_589), .D(n_596), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g1079 ( .A(n_471), .B(n_1080), .C(n_1084), .Y(n_1079) );
NAND4xp25_ASAP7_75t_L g1393 ( .A(n_471), .B(n_1394), .C(n_1397), .D(n_1402), .Y(n_1393) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .C(n_477), .Y(n_472) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .C(n_493), .D(n_501), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .C(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_491), .B(n_919), .C(n_922), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g962 ( .A(n_491), .B(n_963), .C(n_965), .Y(n_962) );
INVx1_ASAP7_75t_L g996 ( .A(n_491), .Y(n_996) );
INVx2_ASAP7_75t_L g621 ( .A(n_498), .Y(n_621) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g1428 ( .A(n_503), .Y(n_1428) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g533 ( .A(n_504), .Y(n_533) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_563), .B1(n_564), .B2(n_639), .Y(n_510) );
INVx2_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
INVx1_ASAP7_75t_L g562 ( .A(n_512), .Y(n_562) );
AOI211x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_526), .B(n_527), .C(n_549), .Y(n_512) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_526), .A2(n_647), .B(n_657), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_526), .A2(n_734), .B(n_743), .Y(n_733) );
OAI31xp33_ASAP7_75t_SL g870 ( .A1(n_526), .A2(n_871), .A3(n_872), .B(n_876), .Y(n_870) );
AOI211xp5_ASAP7_75t_L g887 ( .A1(n_526), .A2(n_888), .B(n_901), .C(n_912), .Y(n_887) );
AOI211xp5_ASAP7_75t_L g936 ( .A1(n_526), .A2(n_937), .B(n_948), .C(n_958), .Y(n_936) );
OAI31xp33_ASAP7_75t_SL g1009 ( .A1(n_526), .A2(n_1010), .A3(n_1011), .B(n_1016), .Y(n_1009) );
OAI31xp33_ASAP7_75t_L g1059 ( .A1(n_526), .A2(n_1060), .A3(n_1061), .B(n_1062), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_540), .Y(n_527) );
INVx1_ASAP7_75t_L g1043 ( .A(n_530), .Y(n_1043) );
BUFx3_ASAP7_75t_L g1126 ( .A(n_530), .Y(n_1126) );
INVx2_ASAP7_75t_SL g603 ( .A(n_536), .Y(n_603) );
INVx4_ASAP7_75t_L g612 ( .A(n_536), .Y(n_612) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_536), .Y(n_1116) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_539), .Y(n_552) );
INVx1_ASAP7_75t_L g577 ( .A(n_542), .Y(n_577) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g1064 ( .A(n_543), .Y(n_1064) );
AOI31xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_555), .A3(n_558), .B(n_560), .Y(n_549) );
AOI31xp33_ASAP7_75t_L g901 ( .A1(n_560), .A2(n_902), .A3(n_907), .B(n_910), .Y(n_901) );
AOI31xp33_ASAP7_75t_L g948 ( .A1(n_560), .A2(n_949), .A3(n_953), .B(n_956), .Y(n_948) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g638 ( .A(n_566), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .C(n_574), .D(n_582), .Y(n_567) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g589 ( .A1(n_578), .A2(n_581), .B1(n_590), .B2(n_592), .C1(n_593), .C2(n_594), .Y(n_589) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND4xp25_ASAP7_75t_SL g1406 ( .A(n_582), .B(n_1407), .C(n_1409), .D(n_1412), .Y(n_1406) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND4xp25_ASAP7_75t_L g888 ( .A(n_583), .B(n_889), .C(n_892), .D(n_898), .Y(n_888) );
NAND4xp25_ASAP7_75t_L g937 ( .A(n_583), .B(n_938), .C(n_941), .D(n_944), .Y(n_937) );
OAI31xp33_ASAP7_75t_L g748 ( .A1(n_584), .A2(n_749), .A3(n_751), .B(n_758), .Y(n_748) );
INVx1_ASAP7_75t_L g1094 ( .A(n_584), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_590), .A2(n_592), .B1(n_756), .B2(n_757), .Y(n_766) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g606 ( .A(n_595), .Y(n_606) );
INVx1_ASAP7_75t_L g1399 ( .A(n_595), .Y(n_1399) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_609), .C(n_616), .D(n_627), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .C(n_607), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_607), .A2(n_1096), .B1(n_1107), .B2(n_1120), .C(n_1122), .Y(n_1095) );
AOI33xp33_ASAP7_75t_L g1430 ( .A1(n_607), .A2(n_1120), .A3(n_1431), .B1(n_1432), .B2(n_1433), .B3(n_1434), .Y(n_1430) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .C(n_624), .Y(n_616) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g634 ( .A(n_623), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_623), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_625), .A2(n_794), .B1(n_834), .B2(n_840), .Y(n_833) );
OAI22xp5_ASAP7_75t_SL g1122 ( .A1(n_625), .A2(n_1001), .B1(n_1123), .B2(n_1127), .Y(n_1122) );
INVx2_ASAP7_75t_L g1418 ( .A(n_625), .Y(n_1418) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .C(n_635), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx4f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx4f_ASAP7_75t_L g795 ( .A(n_636), .Y(n_795) );
INVx4_ASAP7_75t_L g1001 ( .A(n_636), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_637), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
AO22x2_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_1074), .B1(n_1137), .B2(n_1138), .Y(n_640) );
INVx1_ASAP7_75t_L g1137 ( .A(n_641), .Y(n_1137) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_882), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_745), .B1(n_880), .B2(n_881), .Y(n_642) );
INVx2_ASAP7_75t_L g880 ( .A(n_643), .Y(n_880) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_701), .Y(n_643) );
NAND3x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_664), .C(n_679), .Y(n_645) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g737 ( .A(n_651), .Y(n_737) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g798 ( .A(n_660), .Y(n_798) );
INVx1_ASAP7_75t_L g818 ( .A(n_660), .Y(n_818) );
BUFx2_ASAP7_75t_L g841 ( .A(n_660), .Y(n_841) );
INVx1_ASAP7_75t_L g1035 ( .A(n_660), .Y(n_1035) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g754 ( .A(n_661), .B(n_662), .Y(n_754) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx2_ASAP7_75t_L g786 ( .A(n_668), .Y(n_786) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g774 ( .A(n_669), .Y(n_774) );
INVx1_ASAP7_75t_L g854 ( .A(n_669), .Y(n_854) );
INVx5_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g781 ( .A(n_674), .Y(n_781) );
INVx1_ASAP7_75t_L g849 ( .A(n_674), .Y(n_849) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g728 ( .A(n_675), .Y(n_728) );
INVx3_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
INVx2_ASAP7_75t_L g867 ( .A(n_675), .Y(n_867) );
AND4x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_686), .C(n_690), .D(n_698), .Y(n_679) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g986 ( .A(n_684), .Y(n_986) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_692), .Y(n_808) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g1013 ( .A(n_694), .Y(n_1013) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g1031 ( .A(n_697), .Y(n_1031) );
INVx1_ASAP7_75t_L g1135 ( .A(n_697), .Y(n_1135) );
XOR2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_744), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_723), .C(n_733), .Y(n_702) );
AND4x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_708), .C(n_713), .D(n_718), .Y(n_703) );
INVx1_ASAP7_75t_L g776 ( .A(n_706), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .C(n_712), .Y(n_708) );
INVx2_ASAP7_75t_L g782 ( .A(n_712), .Y(n_782) );
INVx1_ASAP7_75t_L g869 ( .A(n_712), .Y(n_869) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_720), .Y(n_1129) );
BUFx2_ASAP7_75t_L g1420 ( .A(n_720), .Y(n_1420) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g896 ( .A(n_738), .Y(n_896) );
INVx1_ASAP7_75t_L g947 ( .A(n_738), .Y(n_947) );
INVx1_ASAP7_75t_L g881 ( .A(n_745), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_821), .B1(n_822), .B2(n_879), .Y(n_745) );
INVx1_ASAP7_75t_L g879 ( .A(n_746), .Y(n_879) );
INVx1_ASAP7_75t_L g819 ( .A(n_747), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_760), .C(n_768), .Y(n_747) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g802 ( .A(n_754), .Y(n_802) );
INVx1_ASAP7_75t_L g844 ( .A(n_754), .Y(n_844) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_754), .Y(n_1006) );
BUFx4f_ASAP7_75t_L g1038 ( .A(n_754), .Y(n_1038) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g827 ( .A(n_765), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_765), .A2(n_1049), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_783), .C(n_807), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_777), .C(n_782), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_775), .B2(n_776), .Y(n_770) );
BUFx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g984 ( .A(n_774), .Y(n_984) );
INVx1_ASAP7_75t_L g1053 ( .A(n_774), .Y(n_1053) );
OAI22xp33_ASAP7_75t_SL g777 ( .A1(n_778), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_779), .A2(n_835), .B1(n_836), .B2(n_849), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_779), .A2(n_978), .B1(n_979), .B2(n_981), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_792), .B1(n_794), .B2(n_796), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_787), .B1(n_788), .B2(n_790), .C(n_791), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI33xp33_ASAP7_75t_L g847 ( .A1(n_792), .A2(n_848), .A3(n_850), .B1(n_858), .B2(n_863), .B3(n_869), .Y(n_847) );
OAI33xp33_ASAP7_75t_L g976 ( .A1(n_792), .A2(n_977), .A3(n_982), .B1(n_987), .B2(n_992), .B3(n_996), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g1047 ( .A1(n_792), .A2(n_996), .A3(n_1048), .B1(n_1051), .B2(n_1052), .B3(n_1056), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_799), .B1(n_800), .B2(n_803), .C(n_804), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_797), .A2(n_800), .B1(n_835), .B2(n_836), .C(n_837), .Y(n_834) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g999 ( .A(n_798), .Y(n_999) );
INVx2_ASAP7_75t_L g1003 ( .A(n_798), .Y(n_1003) );
OAI21xp33_ASAP7_75t_SL g809 ( .A1(n_800), .A2(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_802), .Y(n_1124) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g877 ( .A(n_823), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_832), .C(n_870), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_847), .Y(n_832) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_SL g929 ( .A(n_839), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_843), .B2(n_845), .C(n_846), .Y(n_840) );
BUFx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g874 ( .A(n_844), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_855), .B2(n_856), .Y(n_850) );
INVx2_ASAP7_75t_SL g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g860 ( .A(n_853), .Y(n_860) );
BUFx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
OAI22xp5_ASAP7_75t_SL g858 ( .A1(n_859), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_867), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
OAI221xp5_ASAP7_75t_L g998 ( .A1(n_873), .A2(n_978), .B1(n_981), .B2(n_999), .C(n_1000), .Y(n_998) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
XOR2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_972), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_934), .B2(n_935), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B(n_895), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g944 ( .A1(n_893), .A2(n_945), .B(n_946), .Y(n_944) );
BUFx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND4xp25_ASAP7_75t_L g912 ( .A(n_913), .B(n_918), .C(n_923), .D(n_930), .Y(n_912) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
HB1xp67_ASAP7_75t_L g1425 ( .A(n_932), .Y(n_1425) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND4xp25_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .C(n_966), .D(n_969), .Y(n_958) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_964), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_1022), .B1(n_1072), .B2(n_1073), .Y(n_972) );
INVx1_ASAP7_75t_L g1072 ( .A(n_973), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_1009), .C(n_1017), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_997), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_979), .A2(n_1033), .B1(n_1036), .B2(n_1049), .Y(n_1048) );
INVx2_ASAP7_75t_L g1106 ( .A(n_979), .Y(n_1106) );
BUFx3_ASAP7_75t_L g1119 ( .A(n_979), .Y(n_1119) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
OAI22xp33_ASAP7_75t_SL g982 ( .A1(n_983), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_984), .A2(n_988), .B1(n_989), .B2(n_991), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_984), .A2(n_989), .B1(n_1028), .B2(n_1030), .Y(n_1051) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_989), .A2(n_1053), .B1(n_1054), .B2(n_1055), .Y(n_1052) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_990), .Y(n_1097) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1001), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1004), .B1(n_1005), .B2(n_1007), .C(n_1008), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_1003), .A2(n_1101), .B1(n_1104), .B2(n_1124), .C(n_1125), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1022), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1059), .C(n_1067), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1047), .Y(n_1024) );
OAI33xp33_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .A3(n_1032), .B1(n_1039), .B2(n_1042), .B3(n_1046), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1029), .B1(n_1030), .B2(n_1031), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .B1(n_1036), .B2(n_1037), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1034), .A2(n_1037), .B1(n_1040), .B2(n_1041), .Y(n_1039) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1074), .Y(n_1138) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1095), .Y(n_1076) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_1082), .A2(n_1124), .B1(n_1128), .B2(n_1130), .C(n_1131), .Y(n_1127) );
AOI21xp5_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1091), .B(n_1094), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
OAI22xp5_ASAP7_75t_SL g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1104), .B2(n_1105), .Y(n_1100) );
INVx3_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx3_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI22xp33_ASAP7_75t_SL g1113 ( .A1(n_1114), .A2(n_1115), .B1(n_1117), .B2(n_1118), .Y(n_1113) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
BUFx3_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
OAI221xp5_ASAP7_75t_L g1139 ( .A1(n_1140), .A2(n_1389), .B1(n_1390), .B2(n_1436), .C(n_1440), .Y(n_1139) );
NOR2x1_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1326), .Y(n_1140) );
NAND3xp33_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1247), .C(n_1286), .Y(n_1141) );
OAI21xp5_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1204), .B(n_1222), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1181), .B1(n_1198), .B2(n_1200), .Y(n_1143) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1144), .B(n_1208), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1168), .Y(n_1144) );
CKINVDCx6p67_ASAP7_75t_R g1197 ( .A(n_1145), .Y(n_1197) );
OAI222xp33_ASAP7_75t_L g1204 ( .A1(n_1145), .A2(n_1205), .B1(n_1208), .B2(n_1213), .C1(n_1217), .C2(n_1221), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1145), .B(n_1169), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1145), .B(n_1220), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1145), .B(n_1202), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1145), .B(n_1219), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1145), .B(n_1266), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1145), .B(n_1220), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1145), .B(n_1190), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1145), .B(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1145), .B(n_1293), .Y(n_1332) );
OR2x6_ASAP7_75t_SL g1145 ( .A(n_1146), .B(n_1158), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1154), .B1(n_1155), .B2(n_1157), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1151), .Y(n_1148) );
AND2x4_ASAP7_75t_L g1156 ( .A(n_1149), .B(n_1152), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1185 ( .A(n_1149), .B(n_1151), .Y(n_1185) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1150), .Y(n_1163) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1153), .B(n_1163), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_1155), .A2(n_1244), .B1(n_1245), .B2(n_1246), .Y(n_1243) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_1156), .Y(n_1155) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1156), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1164), .B1(n_1165), .B2(n_1167), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1186 ( .A1(n_1159), .A2(n_1165), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_1159), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_1159), .A2(n_1234), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
BUFx6f_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_1160), .A2(n_1165), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1161), .B(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1161), .Y(n_1173) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1162), .Y(n_1172) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1165), .Y(n_1235) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1166), .Y(n_1175) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1168), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_1168), .A2(n_1288), .B1(n_1294), .B2(n_1297), .C(n_1299), .Y(n_1287) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1168), .B(n_1203), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1177), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1169), .B(n_1177), .Y(n_1190) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1169), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1169), .B(n_1250), .Y(n_1293) );
NOR2xp33_ASAP7_75t_SL g1364 ( .A(n_1169), .B(n_1365), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1176), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1173), .B(n_1175), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1449 ( .A(n_1175), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1177), .B(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1177), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1177), .B(n_1197), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1189), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1182), .B(n_1330), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1182), .B(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1183), .Y(n_1199) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1183), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1183), .B(n_1304), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1183), .B(n_1290), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1184), .B(n_1210), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_1184), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1184), .B(n_1210), .Y(n_1270) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1185), .Y(n_1228) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1185), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1190), .B(n_1203), .Y(n_1202) );
AOI322xp5_ASAP7_75t_L g1376 ( .A1(n_1190), .A2(n_1237), .A3(n_1250), .B1(n_1276), .B2(n_1353), .C1(n_1377), .C2(n_1378), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1191), .B(n_1219), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1191), .B(n_1266), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1197), .Y(n_1191) );
INVx4_ASAP7_75t_L g1203 ( .A(n_1192), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1192), .B(n_1215), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1192), .B(n_1197), .Y(n_1267) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1192), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1192), .B(n_1216), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1192), .B(n_1332), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1192), .B(n_1239), .Y(n_1353) );
A2O1A1Ixp33_ASAP7_75t_SL g1360 ( .A1(n_1192), .A2(n_1361), .B(n_1362), .C(n_1369), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1192), .B(n_1276), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1192), .B(n_1284), .Y(n_1368) );
AND2x6_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_1196), .A2(n_1227), .B1(n_1228), .B2(n_1229), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1197), .B(n_1202), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1197), .B(n_1219), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1197), .B(n_1293), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1197), .B(n_1250), .Y(n_1304) );
NOR3xp33_ASAP7_75t_SL g1345 ( .A(n_1197), .B(n_1203), .C(n_1346), .Y(n_1345) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1197), .B(n_1250), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1197), .B(n_1220), .Y(n_1374) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1203), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1203), .B(n_1215), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1203), .B(n_1254), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1203), .B(n_1218), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1203), .B(n_1292), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1203), .B(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
OAI211xp5_ASAP7_75t_L g1313 ( .A1(n_1208), .A2(n_1314), .B(n_1317), .C(n_1321), .Y(n_1313) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1210), .B(n_1216), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1210), .B(n_1216), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_1210), .A2(n_1250), .B1(n_1251), .B2(n_1253), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1210), .B(n_1239), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1210), .B(n_1238), .Y(n_1272) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1210), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1210), .B(n_1309), .Y(n_1308) );
OAI21xp5_ASAP7_75t_L g1328 ( .A1(n_1210), .A2(n_1329), .B(n_1331), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1210), .B(n_1238), .Y(n_1339) );
O2A1O1Ixp33_ASAP7_75t_L g1379 ( .A1(n_1210), .A2(n_1323), .B(n_1380), .C(n_1381), .Y(n_1379) );
AND2x4_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1215), .B(n_1257), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1215), .B(n_1332), .Y(n_1331) );
INVx2_ASAP7_75t_SL g1276 ( .A(n_1216), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1216), .B(n_1238), .Y(n_1385) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1218), .B(n_1275), .Y(n_1301) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1219), .Y(n_1350) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1221), .Y(n_1298) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1236), .Y(n_1223) );
OAI21xp5_ASAP7_75t_L g1286 ( .A1(n_1224), .A2(n_1287), .B(n_1313), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1224), .B(n_1296), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1225), .B(n_1237), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_1225), .A2(n_1328), .B1(n_1333), .B2(n_1335), .C(n_1337), .Y(n_1327) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1225), .Y(n_1370) );
OR2x6_ASAP7_75t_SL g1225 ( .A(n_1226), .B(n_1230), .Y(n_1225) );
BUFx2_ASAP7_75t_SL g1389 ( .A(n_1233), .Y(n_1389) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1236), .B(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_SL g1236 ( .A(n_1237), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1367 ( .A(n_1237), .B(n_1315), .C(n_1368), .Y(n_1367) );
INVx3_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1238), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1238), .B(n_1296), .Y(n_1347) );
INVx3_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1239), .B(n_1270), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1243), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1271), .Y(n_1247) );
A2O1A1Ixp33_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1255), .B(n_1259), .C(n_1260), .Y(n_1248) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1253), .A2(n_1261), .B1(n_1262), .B2(n_1268), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1254), .B(n_1306), .Y(n_1305) );
INVxp67_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1261), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1261), .B(n_1276), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1264), .Y(n_1386) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1267), .Y(n_1265) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1267), .Y(n_1316) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1269), .B(n_1350), .Y(n_1361) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1270), .Y(n_1359) );
A2O1A1Ixp33_ASAP7_75t_L g1271 ( .A1(n_1272), .A2(n_1273), .B(n_1278), .C(n_1279), .Y(n_1271) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1272), .Y(n_1300) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_1274), .Y(n_1273) );
OAI21xp5_ASAP7_75t_L g1317 ( .A1(n_1274), .A2(n_1318), .B(n_1320), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1277), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1276), .Y(n_1284) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1276), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1277), .B(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1277), .B(n_1359), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_1278), .A2(n_1385), .B1(n_1386), .B2(n_1387), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1285), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_1282), .B(n_1315), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1283), .B(n_1296), .Y(n_1295) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1283), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1283), .B(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1291), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_1291), .A2(n_1338), .B1(n_1346), .B2(n_1363), .C(n_1366), .Y(n_1362) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
OAI21xp5_ASAP7_75t_SL g1355 ( .A1(n_1292), .A2(n_1356), .B(n_1358), .Y(n_1355) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1293), .Y(n_1315) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1296), .Y(n_1388) );
OAI211xp5_ASAP7_75t_L g1372 ( .A1(n_1297), .A2(n_1373), .B(n_1375), .C(n_1376), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1352 ( .A(n_1298), .B(n_1353), .C(n_1354), .Y(n_1352) );
AOI211xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1301), .B(n_1302), .C(n_1312), .Y(n_1299) );
A2O1A1Ixp33_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1305), .B(n_1307), .C(n_1308), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1310), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1315), .B(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1320), .Y(n_1380) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1324), .Y(n_1322) );
NAND3xp33_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1360), .C(n_1371), .Y(n_1326) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
OAI211xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1340), .B(n_1341), .C(n_1355), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
AOI221xp5_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1343), .B1(n_1345), .B2(n_1348), .C(n_1351), .Y(n_1341) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_SL g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
OAI31xp33_ASAP7_75t_SL g1371 ( .A1(n_1369), .A2(n_1372), .A3(n_1379), .B(n_1384), .Y(n_1371) );
CKINVDCx14_ASAP7_75t_R g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx2_ASAP7_75t_SL g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1392), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g1444 ( .A(n_1392), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1430), .Y(n_1416) );
AOI33xp33_ASAP7_75t_L g1417 ( .A1(n_1418), .A2(n_1419), .A3(n_1421), .B1(n_1426), .B2(n_1427), .B3(n_1429), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
BUFx6f_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx2_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVxp33_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
OAI21xp5_ASAP7_75t_L g1448 ( .A1(n_1446), .A2(n_1449), .B(n_1450), .Y(n_1448) );
BUFx2_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
endmodule