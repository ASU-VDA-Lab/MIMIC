module fake_jpeg_8906_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_11),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx2_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_47),
.B1(n_17),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_30),
.B(n_26),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_25),
.B(n_26),
.C(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_60),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_21),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_67),
.Y(n_89)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_77),
.B1(n_53),
.B2(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_32),
.B(n_40),
.C(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_54),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_41),
.B(n_34),
.C(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_84),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_65),
.B1(n_85),
.B2(n_90),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_43),
.B(n_42),
.C(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_56),
.B(n_69),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_88),
.B(n_92),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_61),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_51),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_19),
.B(n_30),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_83),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_68),
.C(n_42),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_70),
.B1(n_72),
.B2(n_68),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_128),
.B1(n_102),
.B2(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_84),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_53),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_130),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_95),
.B(n_87),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_101),
.B(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_108),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_39),
.CI(n_57),
.CON(n_131),
.SN(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_111),
.C(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_140),
.C(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_147),
.B1(n_123),
.B2(n_122),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_41),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_123),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_98),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_101),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_28),
.B(n_27),
.C(n_16),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_97),
.B1(n_87),
.B2(n_86),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_134),
.C(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_149),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_120),
.B(n_116),
.Y(n_155)
);

AOI31xp67_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_142),
.A3(n_137),
.B(n_144),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_120),
.C(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_134),
.C(n_131),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_131),
.C(n_57),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_164),
.B1(n_28),
.B2(n_163),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_148),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_163),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_141),
.B1(n_15),
.B2(n_45),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_185),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_161),
.B(n_162),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_161),
.B(n_160),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_9),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_170),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_189),
.Y(n_195)
);

NOR4xp25_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_165),
.C(n_169),
.D(n_168),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_1),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_175),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_177),
.B(n_180),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_197),
.C(n_192),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_182),
.B(n_2),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_201),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_188),
.C(n_4),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_199),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);


endmodule