module fake_jpeg_14135_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_50),
.B1(n_55),
.B2(n_63),
.Y(n_101)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_18),
.B1(n_31),
.B2(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_52),
.B(n_33),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_68),
.Y(n_93)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_18),
.B1(n_24),
.B2(n_31),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_26),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_77),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_35),
.CI(n_44),
.CON(n_76),
.SN(n_76)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_89),
.CI(n_49),
.CON(n_116),
.SN(n_116)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_45),
.A3(n_40),
.B1(n_37),
.B2(n_19),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_80),
.A2(n_20),
.B(n_32),
.C(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_81),
.B(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_22),
.B1(n_40),
.B2(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_54),
.B1(n_66),
.B2(n_16),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_29),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_29),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_90),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_45),
.C(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_98),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_16),
.B1(n_33),
.B2(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_22),
.B1(n_32),
.B2(n_19),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_73),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_30),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_16),
.B1(n_28),
.B2(n_20),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_28),
.B(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_10),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_49),
.B1(n_65),
.B2(n_60),
.Y(n_111)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_22),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_113),
.A2(n_128),
.B(n_17),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_56),
.B1(n_54),
.B2(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_118),
.B1(n_135),
.B2(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_117),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_107),
.B1(n_76),
.B2(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_74),
.A2(n_53),
.B1(n_32),
.B2(n_28),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_129),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_75),
.B(n_66),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_105),
.B1(n_99),
.B2(n_97),
.Y(n_166)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_103),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_107),
.C(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_144),
.C(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_76),
.B1(n_80),
.B2(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_146),
.B1(n_166),
.B2(n_135),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_96),
.B(n_88),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_131),
.B(n_133),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_100),
.B1(n_81),
.B2(n_85),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_156),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_88),
.B1(n_87),
.B2(n_78),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_92),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_117),
.B(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_106),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_158),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_79),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_168),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_103),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_94),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_99),
.B1(n_17),
.B2(n_14),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_119),
.B(n_14),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_9),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_137),
.B(n_129),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_110),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_115),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_174),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_115),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_117),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_179),
.C(n_194),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_189),
.B(n_199),
.C(n_170),
.D(n_151),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_168),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_187),
.B1(n_198),
.B2(n_142),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_112),
.B1(n_120),
.B2(n_109),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_131),
.B(n_110),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_112),
.B(n_109),
.C(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_165),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_14),
.C(n_13),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_200),
.C(n_203),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_139),
.A2(n_123),
.B(n_1),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_17),
.B1(n_13),
.B2(n_12),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_13),
.C(n_12),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_200),
.Y(n_213)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_178),
.B(n_190),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_201),
.B1(n_181),
.B2(n_193),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_212),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_188),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_157),
.B1(n_9),
.B2(n_2),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_145),
.B1(n_154),
.B2(n_150),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_166),
.B1(n_140),
.B2(n_153),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_151),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_229),
.C(n_176),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_162),
.C(n_141),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_175),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_140),
.B1(n_163),
.B2(n_161),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_233),
.B1(n_1),
.B2(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_236),
.C(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_174),
.C(n_189),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_227),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_213),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_194),
.C(n_182),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_221),
.B(n_222),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_199),
.B(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_198),
.C(n_149),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_257),
.C(n_212),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_207),
.B(n_195),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_256),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_157),
.B1(n_167),
.B2(n_10),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_249),
.B1(n_219),
.B2(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_221),
.B(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_216),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_231),
.C(n_225),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_264),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_263),
.Y(n_283)
);

XOR2x2_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_209),
.Y(n_261)
);

FAx1_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_244),
.CI(n_256),
.CON(n_284),
.SN(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_254),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_236),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_217),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_267),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_224),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_276),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_275),
.B1(n_234),
.B2(n_248),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_215),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_206),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_279),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_243),
.B(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_280),
.A2(n_4),
.B(n_6),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_240),
.B1(n_247),
.B2(n_253),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_249),
.B(n_253),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_4),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_3),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_292),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_264),
.C(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_266),
.C(n_270),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_266),
.B(n_258),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_295),
.A2(n_288),
.B(n_284),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_300),
.B1(n_282),
.B2(n_7),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_272),
.C(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_305),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_304),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_4),
.C(n_7),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_280),
.B1(n_283),
.B2(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_314),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_279),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_312),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_289),
.B1(n_281),
.B2(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_297),
.B1(n_299),
.B2(n_296),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_7),
.B(n_8),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_298),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_320),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_302),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_313),
.B(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_321),
.B(n_307),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_322),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_322),
.B(n_311),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.C(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_320),
.B(n_316),
.Y(n_328)
);

AOI211xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_317),
.B(n_294),
.C(n_308),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_303),
.A3(n_296),
.B1(n_315),
.B2(n_305),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule