module fake_netlist_6_2999_n_2139 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2139);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2139;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2017;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_135),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_96),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_133),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_81),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_43),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_57),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_173),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_113),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_145),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_30),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_39),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_182),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_102),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_129),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_114),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_18),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_161),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_156),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_228),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_96),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_28),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_84),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_28),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_189),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_82),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_150),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_159),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_36),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_109),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_71),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_127),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_152),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_199),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_101),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_61),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_123),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_57),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_39),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_18),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_56),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_70),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_121),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_65),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_177),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_126),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_196),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_117),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_88),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_81),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_23),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_164),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_207),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_146),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_99),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_42),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_120),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_84),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_37),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_140),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_23),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_29),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_43),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_10),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_169),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_49),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_218),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_50),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_151),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_92),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_167),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_79),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_139),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_94),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_100),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_205),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_67),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_26),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_184),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_37),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_91),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_90),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_24),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_193),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_134),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_178),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_87),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_49),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_53),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_48),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_98),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_44),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_86),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_80),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_70),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_222),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_194),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_13),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_111),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_69),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_163),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_105),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_92),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_71),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_10),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_31),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_131),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_83),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_106),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_76),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_98),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_63),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_148),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_35),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_62),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_26),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_55),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_44),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_154),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_110),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_214),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_51),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_34),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_94),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_180),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_31),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_21),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_38),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_190),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_62),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_55),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_19),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_168),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_153),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_33),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_66),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_51),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_112),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_64),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_13),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_211),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_166),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_93),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_32),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_143),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_32),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_122),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_208),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_224),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_191),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_147),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_12),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_210),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_225),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_78),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_99),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_155),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_11),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_176),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_216),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_78),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_24),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_7),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_5),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_221),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_29),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_5),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_72),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_192),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_137),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_130),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_201),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_170),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_38),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_33),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_217),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_14),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_223),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_213),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_80),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_54),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_0),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_88),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_247),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_231),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_237),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_237),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_286),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_301),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_350),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_236),
.B(n_0),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_233),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_237),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_393),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_241),
.B(n_1),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_234),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_237),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_241),
.B(n_1),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_240),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_237),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_237),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_312),
.Y(n_470)
);

BUFx2_ASAP7_75t_SL g471 ( 
.A(n_236),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_251),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_315),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_293),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_337),
.B(n_2),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_239),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_314),
.B(n_2),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_337),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_293),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_252),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_314),
.B(n_4),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_346),
.B(n_6),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_254),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_255),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_253),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_293),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_259),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_293),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_383),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_293),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_282),
.B(n_6),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_262),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_266),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_267),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_268),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_271),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_265),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_279),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_250),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_231),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_281),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_292),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_346),
.B(n_7),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_283),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_287),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_257),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_296),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_231),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_306),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_307),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_322),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_311),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_313),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_318),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_322),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_322),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_322),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_322),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_326),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_328),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_230),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_257),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_269),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_322),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_250),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_380),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_380),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_270),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_380),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_330),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_249),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_249),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_249),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_230),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_340),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_380),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_380),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_347),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_380),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_242),
.B(n_8),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_321),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_321),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_348),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_321),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_354),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_334),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_382),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_382),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_382),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_360),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_366),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_382),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_385),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_242),
.B(n_8),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_389),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_246),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_402),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_246),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_406),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_334),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_246),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_278),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_409),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_250),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_272),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_278),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_297),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_411),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_452),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_523),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_490),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_453),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_500),
.A2(n_304),
.B1(n_339),
.B2(n_336),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_523),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_523),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_509),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_500),
.B(n_250),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_565),
.B(n_341),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_471),
.B(n_444),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_509),
.B(n_334),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_565),
.B(n_341),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_501),
.B(n_292),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_412),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_503),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_467),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_468),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_542),
.B(n_413),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_414),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_416),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_469),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_479),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_277),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_507),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_479),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_454),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_450),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_486),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

CKINVDCx9p33_ASAP7_75t_R g620 ( 
.A(n_462),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_545),
.B(n_422),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_488),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_533),
.B(n_292),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_491),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_493),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_491),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_545),
.B(n_425),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_516),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_516),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_543),
.B(n_434),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_518),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_451),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_503),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_519),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_547),
.B(n_435),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_525),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_527),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_528),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

AND2x2_ASAP7_75t_R g649 ( 
.A(n_526),
.B(n_232),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_465),
.A2(n_374),
.B1(n_394),
.B2(n_358),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_492),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_537),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_538),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_561),
.B(n_370),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_538),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_540),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_458),
.A2(n_290),
.B(n_261),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_540),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_548),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_451),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_451),
.B(n_370),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_549),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_549),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_532),
.B(n_436),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_458),
.B(n_282),
.Y(n_667)
);

CKINVDCx8_ASAP7_75t_R g668 ( 
.A(n_625),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_634),
.B(n_485),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_661),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_581),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_581),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_583),
.A2(n_478),
.B1(n_495),
.B2(n_494),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_581),
.Y(n_675)
);

AND2x6_ASAP7_75t_L g676 ( 
.A(n_610),
.B(n_611),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_588),
.A2(n_475),
.B1(n_482),
.B2(n_481),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_582),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_629),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_637),
.B(n_459),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_634),
.B(n_566),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_582),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_590),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_640),
.B(n_463),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_640),
.B(n_466),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_615),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_578),
.B(n_461),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_590),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_615),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_615),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_615),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_661),
.B(n_532),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_637),
.B(n_472),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_667),
.B(n_504),
.C(n_498),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_580),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_661),
.B(n_483),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_590),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_577),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_593),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_604),
.B(n_484),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_666),
.B(n_487),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_577),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_588),
.A2(n_555),
.B1(n_541),
.B2(n_454),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_609),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_590),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_496),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_597),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_604),
.B(n_461),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_591),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_610),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_651),
.B(n_499),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_597),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_591),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_588),
.A2(n_477),
.B1(n_457),
.B2(n_492),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_625),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_595),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_623),
.B(n_532),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_617),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_595),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_600),
.B(n_502),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_583),
.A2(n_477),
.B1(n_342),
.B2(n_369),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_584),
.A2(n_497),
.B1(n_511),
.B2(n_510),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_505),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_610),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_584),
.B(n_440),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_585),
.B(n_506),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_580),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_597),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_585),
.B(n_508),
.Y(n_735)
);

INVx4_ASAP7_75t_SL g736 ( 
.A(n_610),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_663),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_587),
.B(n_520),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_596),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_SL g740 ( 
.A(n_650),
.B(n_514),
.C(n_513),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_597),
.Y(n_741)
);

INVx6_ASAP7_75t_L g742 ( 
.A(n_610),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_587),
.B(n_521),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_593),
.B(n_531),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_596),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_612),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_650),
.A2(n_638),
.B1(n_395),
.B2(n_319),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_580),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_599),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_610),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_623),
.B(n_536),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_638),
.B(n_539),
.Y(n_752)
);

INVx11_ASAP7_75t_L g753 ( 
.A(n_614),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_599),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_580),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_580),
.Y(n_757)
);

OAI21xp33_ASAP7_75t_SL g758 ( 
.A1(n_658),
.A2(n_440),
.B(n_245),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_612),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_614),
.A2(n_455),
.B1(n_470),
.B2(n_456),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_605),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_667),
.B(n_261),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_601),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_612),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_601),
.B(n_544),
.Y(n_765)
);

BUFx6f_ASAP7_75t_SL g766 ( 
.A(n_586),
.Y(n_766)
);

AND3x2_ASAP7_75t_L g767 ( 
.A(n_575),
.B(n_363),
.C(n_290),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_575),
.Y(n_769)
);

BUFx8_ASAP7_75t_SL g770 ( 
.A(n_617),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_SL g771 ( 
.A(n_655),
.B(n_274),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_598),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_616),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_602),
.B(n_480),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_606),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_624),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_624),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_602),
.B(n_546),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_616),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_616),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_616),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_618),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_586),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_621),
.A2(n_551),
.B1(n_552),
.B2(n_515),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_554),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_610),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_626),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_618),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_257),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_628),
.B(n_556),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_611),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_627),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_598),
.B(n_569),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_586),
.A2(n_355),
.B1(n_428),
.B2(n_297),
.Y(n_796)
);

BUFx6f_ASAP7_75t_SL g797 ( 
.A(n_586),
.Y(n_797)
);

BUFx6f_ASAP7_75t_SL g798 ( 
.A(n_586),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_586),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_631),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_618),
.Y(n_801)
);

INVx5_ASAP7_75t_L g802 ( 
.A(n_611),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_631),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_614),
.B(n_558),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_632),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_622),
.Y(n_806)
);

INVx5_ASAP7_75t_L g807 ( 
.A(n_611),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_622),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_622),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_598),
.B(n_534),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_632),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_598),
.B(n_560),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_658),
.A2(n_428),
.B1(n_355),
.B2(n_426),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_658),
.A2(n_426),
.B1(n_370),
.B2(n_534),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_575),
.B(n_524),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_614),
.B(n_529),
.C(n_522),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_622),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_676),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_799),
.Y(n_820)
);

AND2x2_ASAP7_75t_SL g821 ( 
.A(n_762),
.B(n_363),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_735),
.B(n_669),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_683),
.B(n_614),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_708),
.A2(n_564),
.B1(n_473),
.B2(n_489),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_738),
.A2(n_285),
.B1(n_614),
.B2(n_439),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_686),
.B(n_578),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_670),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_672),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_676),
.B(n_790),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_770),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_727),
.B(n_620),
.C(n_276),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_672),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_687),
.B(n_535),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_703),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_799),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_688),
.B(n_244),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_763),
.B(n_786),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_791),
.A2(n_437),
.B1(n_245),
.B2(n_248),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_795),
.B(n_613),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_737),
.A2(n_248),
.B1(n_256),
.B2(n_244),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_677),
.A2(n_258),
.B1(n_260),
.B2(n_256),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_707),
.B(n_284),
.C(n_275),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_723),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_812),
.B(n_611),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_673),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_702),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_770),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_762),
.A2(n_263),
.B1(n_280),
.B2(n_264),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_673),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_696),
.B(n_264),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_688),
.A2(n_280),
.B1(n_299),
.B2(n_288),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_675),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_729),
.B(n_613),
.Y(n_853)
);

INVxp33_ASAP7_75t_L g854 ( 
.A(n_744),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_711),
.B(n_298),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_SL g856 ( 
.A(n_774),
.B(n_288),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_675),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_726),
.B(n_635),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_815),
.B(n_235),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_765),
.B(n_645),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_815),
.B(n_235),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_690),
.B(n_257),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_706),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_774),
.B(n_341),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_778),
.A2(n_299),
.B1(n_332),
.B2(n_305),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_704),
.B(n_341),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_784),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_710),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_705),
.B(n_300),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_752),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_723),
.B(n_257),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_724),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_758),
.A2(n_692),
.B(n_694),
.C(n_689),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_676),
.B(n_415),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_715),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_696),
.B(n_305),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_715),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_784),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_769),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_689),
.A2(n_361),
.B1(n_365),
.B2(n_332),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_720),
.B(n_361),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_692),
.B(n_645),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_784),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_694),
.B(n_646),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_695),
.B(n_646),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_674),
.B(n_415),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_695),
.B(n_696),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_731),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_719),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_671),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_732),
.B(n_415),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_719),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_671),
.Y(n_894)
);

AND2x6_ASAP7_75t_SL g895 ( 
.A(n_731),
.B(n_238),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_772),
.B(n_648),
.Y(n_896)
);

OAI22xp33_ASAP7_75t_L g897 ( 
.A1(n_731),
.A2(n_373),
.B1(n_377),
.B2(n_371),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_693),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_722),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_813),
.A2(n_384),
.B1(n_397),
.B2(n_377),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_785),
.B(n_415),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_731),
.A2(n_397),
.B1(n_398),
.B2(n_384),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_751),
.B(n_303),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_740),
.B(n_620),
.C(n_310),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_722),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_771),
.A2(n_405),
.B1(n_418),
.B2(n_398),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_713),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_771),
.A2(n_418),
.B1(n_419),
.B2(n_405),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_725),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_682),
.B(n_415),
.Y(n_910)
);

NOR2x1p5_ASAP7_75t_L g911 ( 
.A(n_816),
.B(n_698),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_697),
.B(n_424),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_725),
.B(n_557),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_739),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_745),
.B(n_749),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_721),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_743),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_745),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_700),
.B(n_430),
.Y(n_919)
);

INVx8_ASAP7_75t_L g920 ( 
.A(n_766),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_693),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_754),
.B(n_557),
.Y(n_922)
);

AND2x2_ASAP7_75t_SL g923 ( 
.A(n_814),
.B(n_438),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_754),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_756),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_L g926 ( 
.A(n_676),
.B(n_438),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_761),
.B(n_652),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_761),
.B(n_559),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_728),
.B(n_442),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_747),
.B(n_309),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_721),
.B(n_238),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_775),
.B(n_654),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_776),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_777),
.B(n_654),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_777),
.B(n_571),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_788),
.B(n_571),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_788),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_716),
.B(n_442),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_793),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_794),
.B(n_572),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_699),
.Y(n_941)
);

AO22x2_ASAP7_75t_L g942 ( 
.A1(n_804),
.A2(n_445),
.B1(n_338),
.B2(n_335),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_716),
.B(n_317),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_668),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_800),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_803),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_805),
.Y(n_947)
);

CKINVDCx6p67_ASAP7_75t_R g948 ( 
.A(n_668),
.Y(n_948)
);

NAND3xp33_ASAP7_75t_L g949 ( 
.A(n_796),
.B(n_767),
.C(n_818),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_716),
.B(n_323),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_805),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_811),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_811),
.B(n_572),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_766),
.A2(n_797),
.B1(n_798),
.B2(n_818),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_699),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_678),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_678),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_810),
.B(n_594),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_730),
.B(n_594),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_730),
.B(n_594),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_730),
.B(n_603),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_797),
.A2(n_426),
.B1(n_664),
.B2(n_603),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_797),
.A2(n_798),
.B1(n_790),
.B2(n_679),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_760),
.B(n_243),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_787),
.B(n_607),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_837),
.B(n_680),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_874),
.A2(n_681),
.B(n_680),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_822),
.A2(n_681),
.B(n_792),
.C(n_787),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_864),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_833),
.B(n_680),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_853),
.B(n_733),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_858),
.B(n_733),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_860),
.B(n_733),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_L g974 ( 
.A(n_879),
.B(n_676),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_826),
.A2(n_273),
.B(n_289),
.C(n_243),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_855),
.B(n_748),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_870),
.B(n_748),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_888),
.A2(n_681),
.B(n_748),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_839),
.A2(n_802),
.B(n_750),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_824),
.B(n_325),
.C(n_324),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_819),
.B(n_736),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_854),
.B(n_753),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_871),
.B(n_563),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_894),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_854),
.B(n_753),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_923),
.B(n_757),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_923),
.B(n_699),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_894),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_841),
.A2(n_685),
.B(n_691),
.C(n_684),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_862),
.A2(n_289),
.B(n_291),
.C(n_273),
.Y(n_990)
);

OAI321xp33_ASAP7_75t_L g991 ( 
.A1(n_930),
.A2(n_908),
.A3(n_929),
.B1(n_906),
.B2(n_897),
.C(n_866),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_875),
.A2(n_807),
.B(n_736),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_875),
.A2(n_807),
.B(n_736),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_862),
.B(n_798),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_882),
.A2(n_294),
.B(n_291),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_821),
.A2(n_691),
.B(n_685),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_924),
.B(n_699),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_819),
.A2(n_807),
.B(n_714),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_894),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_903),
.A2(n_329),
.B(n_327),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_887),
.A2(n_709),
.B(n_712),
.C(n_701),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_829),
.A2(n_714),
.B(n_699),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_829),
.A2(n_755),
.B(n_714),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_843),
.B(n_333),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_821),
.B(n_714),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_864),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_882),
.A2(n_917),
.B(n_856),
.C(n_848),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_836),
.A2(n_709),
.B(n_701),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_955),
.A2(n_868),
.B(n_959),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_901),
.A2(n_718),
.B(n_734),
.C(n_712),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_924),
.B(n_755),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_838),
.B(n_345),
.C(n_344),
.Y(n_1012)
);

CKINVDCx6p67_ASAP7_75t_R g1013 ( 
.A(n_948),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_960),
.A2(n_734),
.B(n_718),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_894),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_879),
.B(n_755),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_846),
.B(n_755),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_846),
.B(n_741),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_863),
.B(n_741),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_859),
.B(n_563),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_842),
.A2(n_353),
.B(n_351),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_868),
.A2(n_576),
.B(n_742),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_856),
.A2(n_294),
.B(n_295),
.C(n_302),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_907),
.B(n_356),
.Y(n_1024)
);

AND2x2_ASAP7_75t_SL g1025 ( 
.A(n_831),
.B(n_825),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_867),
.B(n_359),
.C(n_357),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_863),
.B(n_746),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_961),
.A2(n_576),
.B(n_742),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_869),
.B(n_746),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_827),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_931),
.B(n_964),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_869),
.B(n_817),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_876),
.B(n_817),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_876),
.B(n_759),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_965),
.A2(n_576),
.B(n_742),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_836),
.A2(n_764),
.B(n_759),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_890),
.B(n_809),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_900),
.A2(n_742),
.B1(n_808),
.B2(n_806),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_958),
.A2(n_576),
.B(n_580),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_859),
.B(n_567),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_931),
.B(n_362),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_883),
.A2(n_576),
.B(n_764),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_885),
.A2(n_773),
.B(n_768),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_894),
.Y(n_1044)
);

INVx11_ASAP7_75t_L g1045 ( 
.A(n_948),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_890),
.B(n_779),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_886),
.A2(n_780),
.B(n_779),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_920),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_899),
.B(n_809),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_911),
.A2(n_820),
.B1(n_835),
.B2(n_904),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_879),
.B(n_780),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_844),
.A2(n_782),
.B(n_781),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_893),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_899),
.B(n_808),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_873),
.B(n_364),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_893),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_964),
.B(n_367),
.Y(n_1057)
);

NOR2x1p5_ASAP7_75t_L g1058 ( 
.A(n_830),
.B(n_649),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_914),
.B(n_781),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_891),
.B(n_295),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_879),
.Y(n_1061)
);

BUFx8_ASAP7_75t_SL g1062 ( 
.A(n_830),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_865),
.B(n_372),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_919),
.A2(n_790),
.B1(n_801),
.B2(n_806),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_914),
.A2(n_801),
.B1(n_789),
.B2(n_783),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_920),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_789),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_933),
.A2(n_308),
.B(n_316),
.C(n_320),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_828),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_L g1070 ( 
.A(n_880),
.B(n_379),
.C(n_378),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_L g1071 ( 
.A(n_920),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_850),
.A2(n_790),
.B1(n_607),
.B2(n_608),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_920),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_884),
.A2(n_898),
.B(n_891),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_834),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_945),
.B(n_608),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_884),
.A2(n_573),
.B(n_570),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_573),
.B(n_570),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_916),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_884),
.B(n_629),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_884),
.B(n_629),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_951),
.A2(n_579),
.B(n_574),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_850),
.A2(n_608),
.B1(n_619),
.B2(n_657),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_861),
.B(n_944),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_861),
.B(n_381),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_905),
.B(n_629),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_951),
.A2(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_921),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_896),
.A2(n_579),
.B(n_574),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_828),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_832),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_579),
.B(n_574),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_878),
.B(n_619),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_925),
.B(n_391),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_926),
.A2(n_642),
.B(n_636),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_832),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_937),
.B(n_619),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_946),
.B(n_630),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_916),
.B(n_567),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_926),
.A2(n_642),
.B(n_636),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_845),
.A2(n_642),
.B(n_636),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_845),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_905),
.B(n_630),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_849),
.A2(n_647),
.B(n_643),
.Y(n_1104)
);

AO21x1_ASAP7_75t_L g1105 ( 
.A1(n_823),
.A2(n_331),
.B(n_320),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_954),
.A2(n_433),
.B1(n_392),
.B2(n_396),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_849),
.A2(n_857),
.B(n_852),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_889),
.B(n_399),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_909),
.B(n_629),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_909),
.B(n_630),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_872),
.A2(n_432),
.B(n_335),
.C(n_338),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_941),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_939),
.B(n_630),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_939),
.A2(n_639),
.B(n_630),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_947),
.B(n_639),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_941),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_850),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_963),
.A2(n_952),
.B1(n_902),
.B2(n_962),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_938),
.A2(n_656),
.B(n_662),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_913),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_949),
.B(n_943),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_950),
.A2(n_656),
.B(n_662),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_935),
.A2(n_656),
.B(n_662),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_936),
.A2(n_643),
.B(n_647),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_913),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_940),
.A2(n_653),
.B(n_659),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_922),
.B(n_928),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_912),
.A2(n_331),
.B(n_343),
.C(n_432),
.Y(n_1128)
);

BUFx8_ASAP7_75t_L g1129 ( 
.A(n_1075),
.Y(n_1129)
);

INVx6_ASAP7_75t_L g1130 ( 
.A(n_1066),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_SL g1131 ( 
.A(n_1031),
.B(n_847),
.C(n_401),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1008),
.A2(n_892),
.B(n_877),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1031),
.B(n_895),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1053),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1106),
.B(n_847),
.C(n_403),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_969),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1127),
.B(n_1025),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1025),
.A2(n_400),
.B1(n_404),
.B2(n_408),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1084),
.B(n_877),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1006),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1056),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1099),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1057),
.A2(n_840),
.B(n_927),
.C(n_934),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_988),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1066),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1066),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1036),
.A2(n_953),
.B(n_932),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1120),
.B(n_922),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1062),
.B(n_928),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1053),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1041),
.B(n_910),
.C(n_420),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1125),
.B(n_942),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1041),
.B(n_956),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_987),
.A2(n_942),
.B1(n_881),
.B2(n_851),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_994),
.A2(n_942),
.B1(n_956),
.B2(n_957),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_983),
.B(n_942),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1024),
.B(n_957),
.Y(n_1157)
);

BUFx8_ASAP7_75t_SL g1158 ( 
.A(n_1079),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_994),
.A2(n_1061),
.B1(n_986),
.B2(n_1005),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1066),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1013),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_L g1162 ( 
.A(n_991),
.B(n_443),
.C(n_410),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1048),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1085),
.B(n_568),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1085),
.B(n_639),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1050),
.B(n_649),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1024),
.B(n_423),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_988),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1061),
.A2(n_427),
.B1(n_429),
.B2(n_431),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1020),
.B(n_568),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_970),
.B(n_641),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_967),
.A2(n_665),
.B(n_659),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1048),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1117),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_980),
.A2(n_448),
.B1(n_349),
.B2(n_352),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1040),
.B(n_641),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1121),
.A2(n_985),
.B1(n_982),
.B2(n_1026),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_988),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_966),
.A2(n_665),
.B(n_659),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_976),
.A2(n_641),
.B(n_657),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_977),
.A2(n_641),
.B(n_657),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_985),
.A2(n_449),
.B1(n_343),
.B2(n_446),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_974),
.A2(n_971),
.B(n_1009),
.Y(n_1183)
);

INVx3_ASAP7_75t_SL g1184 ( 
.A(n_1055),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1060),
.B(n_641),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1000),
.B(n_349),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1088),
.B(n_559),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1060),
.B(n_1094),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_R g1189 ( 
.A(n_1071),
.B(n_107),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1016),
.A2(n_550),
.B(n_553),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1005),
.A2(n_446),
.B1(n_368),
.B2(n_375),
.Y(n_1191)
);

INVx6_ASAP7_75t_L g1192 ( 
.A(n_1088),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_972),
.A2(n_657),
.B(n_660),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_973),
.A2(n_657),
.B(n_660),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1045),
.Y(n_1195)
);

OAI22x1_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_407),
.B1(n_448),
.B2(n_447),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1094),
.B(n_352),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1063),
.A2(n_990),
.B(n_1004),
.C(n_1118),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1030),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_1071),
.B(n_108),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1004),
.B(n_368),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_975),
.A2(n_417),
.B(n_376),
.C(n_447),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1088),
.B(n_562),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1051),
.A2(n_553),
.B(n_562),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_975),
.A2(n_441),
.B(n_421),
.C(n_417),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_990),
.B(n_375),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_988),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1088),
.B(n_376),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1063),
.B(n_1093),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_SL g1210 ( 
.A1(n_1070),
.A2(n_441),
.B(n_421),
.C(n_407),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_999),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1108),
.B(n_386),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_978),
.A2(n_660),
.B(n_644),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1069),
.Y(n_1214)
);

XNOR2xp5_ASAP7_75t_L g1215 ( 
.A(n_1012),
.B(n_115),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1090),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_999),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_999),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1108),
.A2(n_644),
.B(n_633),
.C(n_629),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1021),
.A2(n_644),
.B(n_633),
.C(n_629),
.Y(n_1220)
);

CKINVDCx8_ASAP7_75t_R g1221 ( 
.A(n_999),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1087),
.B(n_9),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_995),
.A2(n_660),
.B1(n_644),
.B2(n_633),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_L g1224 ( 
.A1(n_1105),
.A2(n_229),
.B(n_206),
.C(n_202),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1097),
.B(n_629),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1091),
.B(n_633),
.Y(n_1226)
);

HAxp5_ASAP7_75t_L g1227 ( 
.A(n_1023),
.B(n_9),
.CON(n_1227),
.SN(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1044),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_968),
.A2(n_660),
.B(n_644),
.Y(n_1229)
);

NOR3xp33_ASAP7_75t_SL g1230 ( 
.A(n_1023),
.B(n_11),
.C(n_14),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1096),
.Y(n_1231)
);

AO32x1_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1102),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_SL g1234 ( 
.A(n_1068),
.B(n_15),
.C(n_16),
.Y(n_1234)
);

CKINVDCx6p67_ASAP7_75t_R g1235 ( 
.A(n_1044),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1076),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1018),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_984),
.B(n_17),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1074),
.A2(n_633),
.B(n_21),
.C(n_22),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1051),
.A2(n_633),
.B(n_197),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_997),
.B(n_633),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1011),
.B(n_20),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1073),
.B(n_633),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1073),
.B(n_195),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1044),
.B(n_188),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1078),
.A2(n_186),
.B(n_183),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1068),
.A2(n_22),
.B(n_25),
.C(n_27),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1044),
.Y(n_1248)
);

O2A1O1Ixp5_ASAP7_75t_SL g1249 ( 
.A1(n_1086),
.A2(n_25),
.B(n_35),
.C(n_40),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1017),
.A2(n_1015),
.B1(n_984),
.B2(n_1067),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1082),
.A2(n_181),
.B(n_174),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1015),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1092),
.A2(n_171),
.B(n_165),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1019),
.A2(n_160),
.B1(n_157),
.B2(n_144),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1112),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1027),
.A2(n_142),
.B1(n_138),
.B2(n_136),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_996),
.A2(n_128),
.B(n_124),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1029),
.Y(n_1258)
);

AO21x1_ASAP7_75t_L g1259 ( 
.A1(n_1080),
.A2(n_40),
.B(n_41),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1039),
.A2(n_118),
.B(n_119),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1098),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_992),
.A2(n_100),
.B(n_46),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_1112),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_45),
.B(n_47),
.C(n_50),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1112),
.B(n_1116),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_981),
.A2(n_47),
.B(n_52),
.C(n_53),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1083),
.A2(n_52),
.B(n_54),
.C(n_56),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_R g1268 ( 
.A(n_1112),
.B(n_58),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1116),
.B(n_58),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1116),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1002),
.A2(n_59),
.B(n_60),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1032),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1003),
.A2(n_63),
.B(n_65),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1022),
.A2(n_66),
.B(n_67),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1033),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_SL g1276 ( 
.A1(n_1111),
.A2(n_1114),
.B(n_1010),
.C(n_1128),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1014),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1080),
.A2(n_68),
.B(n_72),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1042),
.A2(n_68),
.B(n_73),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1198),
.A2(n_1047),
.B(n_1043),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1164),
.B(n_1059),
.Y(n_1281)
);

AO22x2_ASAP7_75t_L g1282 ( 
.A1(n_1166),
.A2(n_1081),
.B1(n_1054),
.B2(n_1049),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1188),
.A2(n_1034),
.B1(n_1046),
.B2(n_1037),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1147),
.A2(n_1052),
.B(n_1107),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1129),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1143),
.A2(n_1089),
.B(n_1081),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1214),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1219),
.A2(n_1038),
.A3(n_979),
.B(n_1122),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1257),
.A2(n_1086),
.B(n_1109),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1167),
.A2(n_1109),
.B(n_1103),
.C(n_1110),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1136),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_SL g1292 ( 
.A(n_1212),
.B(n_1072),
.C(n_1064),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1186),
.A2(n_1001),
.B(n_1035),
.C(n_1028),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1209),
.B(n_1113),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_L g1295 ( 
.A(n_1222),
.B(n_1126),
.C(n_1124),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1153),
.A2(n_993),
.B1(n_1115),
.B2(n_998),
.Y(n_1296)
);

AO22x1_ASAP7_75t_L g1297 ( 
.A1(n_1133),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1142),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_1195),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1177),
.B(n_1077),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1140),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1163),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1184),
.A2(n_1095),
.B1(n_1100),
.B2(n_1123),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1141),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1149),
.B(n_1119),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1139),
.B(n_1104),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1129),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1137),
.A2(n_1101),
.B1(n_75),
.B2(n_76),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1132),
.A2(n_74),
.B(n_77),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1201),
.B(n_1170),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1216),
.Y(n_1311)
);

OAI22x1_ASAP7_75t_L g1312 ( 
.A1(n_1182),
.A2(n_77),
.B1(n_79),
.B2(n_82),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1163),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1263),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1174),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1236),
.B(n_97),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1255),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1162),
.B(n_85),
.C(n_86),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1229),
.A2(n_85),
.B(n_87),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1197),
.A2(n_89),
.B(n_91),
.C(n_95),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1172),
.A2(n_1213),
.B(n_1220),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1161),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1275),
.B(n_1237),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1157),
.B(n_1138),
.Y(n_1324)
);

OAI22x1_ASAP7_75t_L g1325 ( 
.A1(n_1215),
.A2(n_1269),
.B1(n_1156),
.B2(n_1242),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1175),
.B(n_1151),
.C(n_1261),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1199),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1165),
.A2(n_1159),
.B(n_1171),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1158),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1264),
.A2(n_1267),
.B(n_1239),
.C(n_1245),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1148),
.B(n_1169),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1228),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1258),
.B(n_1208),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1213),
.A2(n_1253),
.A3(n_1259),
.B(n_1250),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1176),
.B(n_1152),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1225),
.A2(n_1241),
.B(n_1246),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1231),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1251),
.A2(n_1180),
.B(n_1181),
.Y(n_1338)
);

AO32x2_ASAP7_75t_L g1339 ( 
.A1(n_1191),
.A2(n_1154),
.A3(n_1272),
.B1(n_1254),
.B2(n_1256),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1185),
.B(n_1233),
.Y(n_1340)
);

AOI211x1_ASAP7_75t_L g1341 ( 
.A1(n_1271),
.A2(n_1273),
.B(n_1279),
.C(n_1274),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1192),
.A2(n_1221),
.B1(n_1207),
.B2(n_1134),
.Y(n_1342)
);

AOI31xp67_ASAP7_75t_L g1343 ( 
.A1(n_1206),
.A2(n_1243),
.A3(n_1226),
.B(n_1150),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1276),
.A2(n_1260),
.B(n_1181),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1238),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1146),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1268),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1260),
.A2(n_1180),
.B(n_1277),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1252),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1196),
.A2(n_1230),
.B1(n_1234),
.B2(n_1131),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1274),
.A2(n_1279),
.B(n_1271),
.C(n_1273),
.Y(n_1351)
);

BUFx2_ASAP7_75t_R g1352 ( 
.A(n_1244),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1135),
.Y(n_1353)
);

AO21x1_ASAP7_75t_L g1354 ( 
.A1(n_1262),
.A2(n_1247),
.B(n_1205),
.Y(n_1354)
);

INVx5_ASAP7_75t_SL g1355 ( 
.A(n_1235),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1270),
.B(n_1163),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1210),
.A2(n_1203),
.B(n_1187),
.C(n_1265),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1278),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1202),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_SL g1360 ( 
.A1(n_1144),
.A2(n_1178),
.B(n_1168),
.C(n_1277),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1146),
.B(n_1145),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1193),
.A2(n_1194),
.B(n_1179),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1193),
.A2(n_1194),
.B(n_1179),
.Y(n_1363)
);

OR2x4_ASAP7_75t_L g1364 ( 
.A(n_1173),
.B(n_1145),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1144),
.Y(n_1365)
);

INVxp67_ASAP7_75t_SL g1366 ( 
.A(n_1217),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1224),
.A2(n_1240),
.B(n_1190),
.C(n_1204),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1211),
.A2(n_1248),
.B(n_1178),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1173),
.B(n_1145),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1211),
.A2(n_1248),
.B(n_1218),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1223),
.A2(n_1249),
.B(n_1192),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1217),
.A2(n_1218),
.B(n_1160),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1217),
.B(n_1218),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1227),
.A2(n_1160),
.B(n_1189),
.C(n_1200),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1160),
.A2(n_1266),
.B(n_1232),
.C(n_1130),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_730),
.B(n_716),
.Y(n_1376)
);

NOR2xp67_ASAP7_75t_L g1377 ( 
.A(n_1130),
.B(n_1232),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1130),
.B(n_822),
.Y(n_1378)
);

BUFx2_ASAP7_75t_R g1379 ( 
.A(n_1158),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1142),
.B(n_1031),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1142),
.B(n_724),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1198),
.A2(n_822),
.B(n_826),
.C(n_837),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1129),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1167),
.B(n_822),
.C(n_826),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1164),
.B(n_822),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1167),
.B(n_822),
.C(n_826),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1183),
.A2(n_730),
.B(n_716),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1164),
.B(n_822),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1219),
.A2(n_1155),
.A3(n_1198),
.B(n_1183),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1198),
.A2(n_822),
.B(n_826),
.C(n_837),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1142),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1167),
.B(n_822),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1136),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1142),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1164),
.B(n_822),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1164),
.B(n_822),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1129),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1142),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1198),
.A2(n_822),
.B(n_826),
.C(n_837),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1198),
.A2(n_822),
.B(n_826),
.C(n_837),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1163),
.B(n_1048),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1195),
.B(n_880),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1214),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1214),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1164),
.B(n_822),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_SL g1406 ( 
.A1(n_1198),
.A2(n_1007),
.B(n_823),
.C(n_990),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1136),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1198),
.A2(n_822),
.B(n_837),
.Y(n_1408)
);

OAI21xp33_ASAP7_75t_L g1409 ( 
.A1(n_1212),
.A2(n_822),
.B(n_826),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1219),
.A2(n_1155),
.A3(n_1198),
.B(n_1183),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1219),
.A2(n_1155),
.A3(n_1198),
.B(n_1183),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1164),
.B(n_822),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1129),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1137),
.A2(n_822),
.B1(n_826),
.B2(n_833),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1198),
.A2(n_822),
.B(n_837),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1163),
.B(n_1048),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1136),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1184),
.Y(n_1418)
);

AO32x2_ASAP7_75t_L g1419 ( 
.A1(n_1155),
.A2(n_841),
.A3(n_1159),
.B1(n_1191),
.B2(n_1154),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1158),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1255),
.B(n_1066),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1167),
.B(n_822),
.C(n_826),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1136),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1164),
.B(n_822),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1164),
.B(n_822),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1163),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1129),
.Y(n_1427)
);

CKINVDCx12_ASAP7_75t_R g1428 ( 
.A(n_1139),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1212),
.A2(n_826),
.B1(n_822),
.B2(n_747),
.C(n_727),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_SL g1430 ( 
.A(n_1167),
.B(n_822),
.C(n_826),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1164),
.B(n_822),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1155),
.A2(n_841),
.A3(n_1159),
.B1(n_1191),
.B2(n_1154),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1198),
.A2(n_822),
.B(n_826),
.C(n_837),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1291),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1392),
.A2(n_1409),
.B1(n_1422),
.B2(n_1384),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1329),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1304),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1393),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1324),
.A2(n_1386),
.B1(n_1422),
.B2(n_1384),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1302),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1299),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1409),
.A2(n_1430),
.B1(n_1386),
.B2(n_1429),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1407),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1417),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1364),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1418),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1414),
.A2(n_1326),
.B(n_1350),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1420),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1364),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1423),
.Y(n_1452)
);

CKINVDCx14_ASAP7_75t_R g1453 ( 
.A(n_1314),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1414),
.A2(n_1425),
.B1(n_1405),
.B2(n_1431),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1401),
.Y(n_1455)
);

BUFx2_ASAP7_75t_SL g1456 ( 
.A(n_1402),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1408),
.A2(n_1415),
.B1(n_1318),
.B2(n_1326),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1353),
.A2(n_1412),
.B1(n_1424),
.B2(n_1395),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1385),
.A2(n_1396),
.B1(n_1388),
.B2(n_1350),
.Y(n_1459)
);

CKINVDCx6p67_ASAP7_75t_R g1460 ( 
.A(n_1427),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1382),
.A2(n_1433),
.B1(n_1400),
.B2(n_1399),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1318),
.A2(n_1312),
.B1(n_1325),
.B2(n_1331),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1292),
.A2(n_1308),
.B1(n_1333),
.B2(n_1354),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1379),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1390),
.B(n_1323),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1308),
.A2(n_1359),
.B1(n_1281),
.B2(n_1309),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1322),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1316),
.A2(n_1345),
.B1(n_1378),
.B2(n_1294),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1374),
.A2(n_1391),
.B1(n_1298),
.B2(n_1398),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1327),
.Y(n_1470)
);

BUFx8_ASAP7_75t_SL g1471 ( 
.A(n_1285),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1298),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1287),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1391),
.Y(n_1474)
);

INVx8_ASAP7_75t_L g1475 ( 
.A(n_1421),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1421),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1428),
.A2(n_1347),
.B1(n_1305),
.B2(n_1398),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_SL g1478 ( 
.A(n_1307),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1381),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1305),
.A2(n_1394),
.B1(n_1315),
.B2(n_1413),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1332),
.Y(n_1481)
);

BUFx8_ASAP7_75t_L g1482 ( 
.A(n_1383),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1311),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1282),
.A2(n_1335),
.B1(n_1283),
.B2(n_1295),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1352),
.A2(n_1282),
.B1(n_1351),
.B2(n_1356),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1295),
.A2(n_1404),
.B1(n_1403),
.B2(n_1337),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1299),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1302),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1313),
.Y(n_1489)
);

BUFx4_ASAP7_75t_R g1490 ( 
.A(n_1365),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1340),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1300),
.A2(n_1306),
.B1(n_1280),
.B2(n_1286),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1280),
.A2(n_1344),
.B1(n_1328),
.B2(n_1358),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1313),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1397),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1349),
.Y(n_1496)
);

BUFx4f_ASAP7_75t_SL g1497 ( 
.A(n_1313),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1426),
.Y(n_1498)
);

BUFx8_ASAP7_75t_SL g1499 ( 
.A(n_1317),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1421),
.A2(n_1341),
.B1(n_1416),
.B2(n_1317),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1297),
.A2(n_1377),
.B1(n_1426),
.B2(n_1321),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1426),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1346),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1366),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1321),
.A2(n_1338),
.B1(n_1289),
.B2(n_1319),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1373),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1355),
.B(n_1361),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1361),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1360),
.Y(n_1509)
);

CKINVDCx6p67_ASAP7_75t_R g1510 ( 
.A(n_1355),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1338),
.A2(n_1303),
.B1(n_1284),
.B2(n_1419),
.Y(n_1511)
);

BUFx2_ASAP7_75t_SL g1512 ( 
.A(n_1346),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1320),
.B(n_1406),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1284),
.A2(n_1432),
.B1(n_1419),
.B2(n_1363),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1342),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1343),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1290),
.A2(n_1375),
.B(n_1293),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1372),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1355),
.B(n_1432),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1419),
.A2(n_1432),
.B1(n_1362),
.B2(n_1348),
.Y(n_1520)
);

NAND2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1370),
.B(n_1368),
.Y(n_1521)
);

INVx6_ASAP7_75t_L g1522 ( 
.A(n_1357),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1296),
.B(n_1336),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1339),
.A2(n_1330),
.B1(n_1371),
.B2(n_1376),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1389),
.B(n_1411),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1387),
.Y(n_1526)
);

BUFx10_ASAP7_75t_L g1527 ( 
.A(n_1339),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1339),
.A2(n_1334),
.B1(n_1411),
.B2(n_1410),
.Y(n_1528)
);

CKINVDCx6p67_ASAP7_75t_R g1529 ( 
.A(n_1367),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1389),
.A2(n_1410),
.B1(n_1411),
.B2(n_1334),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1410),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1334),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1288),
.B(n_1310),
.Y(n_1533)
);

BUFx8_ASAP7_75t_SL g1534 ( 
.A(n_1288),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1288),
.A2(n_1409),
.B1(n_1392),
.B2(n_1430),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1298),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1291),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1324),
.B2(n_1384),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1379),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1302),
.Y(n_1542)
);

BUFx8_ASAP7_75t_L g1543 ( 
.A(n_1285),
.Y(n_1543)
);

BUFx2_ASAP7_75t_R g1544 ( 
.A(n_1427),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1545)
);

CKINVDCx11_ASAP7_75t_R g1546 ( 
.A(n_1329),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1369),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1548)
);

BUFx8_ASAP7_75t_L g1549 ( 
.A(n_1285),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1299),
.Y(n_1550)
);

INVx5_ASAP7_75t_L g1551 ( 
.A(n_1421),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1324),
.B2(n_1384),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1291),
.Y(n_1555)
);

CKINVDCx6p67_ASAP7_75t_R g1556 ( 
.A(n_1418),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1430),
.B2(n_1409),
.Y(n_1557)
);

CKINVDCx6p67_ASAP7_75t_R g1558 ( 
.A(n_1418),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1364),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1409),
.B2(n_1386),
.Y(n_1562)
);

CKINVDCx11_ASAP7_75t_R g1563 ( 
.A(n_1329),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1364),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1291),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1384),
.A2(n_1386),
.B1(n_1422),
.B2(n_1392),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_1329),
.Y(n_1570)
);

CKINVDCx6p67_ASAP7_75t_R g1571 ( 
.A(n_1418),
.Y(n_1571)
);

INVx4_ASAP7_75t_SL g1572 ( 
.A(n_1364),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1346),
.B(n_1146),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1299),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1364),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1291),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1329),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1302),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1409),
.B2(n_1386),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1291),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1421),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1324),
.B2(n_1384),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1291),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1291),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1291),
.Y(n_1588)
);

CKINVDCx6p67_ASAP7_75t_R g1589 ( 
.A(n_1418),
.Y(n_1589)
);

BUFx8_ASAP7_75t_L g1590 ( 
.A(n_1285),
.Y(n_1590)
);

INVx8_ASAP7_75t_L g1591 ( 
.A(n_1364),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1291),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1291),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1302),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1291),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1364),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1392),
.A2(n_822),
.B1(n_1324),
.B2(n_1384),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1430),
.B2(n_1386),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1302),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1379),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1291),
.Y(n_1602)
);

CKINVDCx11_ASAP7_75t_R g1603 ( 
.A(n_1329),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1454),
.B(n_1557),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1454),
.B(n_1539),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1437),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1531),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1525),
.Y(n_1608)
);

INVx5_ASAP7_75t_SL g1609 ( 
.A(n_1529),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1540),
.A2(n_1585),
.B1(n_1597),
.B2(n_1552),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1527),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1527),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1441),
.A2(n_1559),
.B1(n_1567),
.B2(n_1537),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1528),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1532),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1533),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1452),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1565),
.B(n_1600),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1546),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1516),
.A2(n_1461),
.A3(n_1435),
.B(n_1579),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1551),
.Y(n_1622)
);

AOI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1523),
.A2(n_1513),
.B(n_1509),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1562),
.A2(n_1444),
.B1(n_1568),
.B2(n_1545),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1458),
.B(n_1438),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1443),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1568),
.A2(n_1459),
.B1(n_1462),
.B2(n_1554),
.C(n_1553),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1475),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1475),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1561),
.B(n_1569),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1534),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1505),
.A2(n_1493),
.B(n_1492),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1434),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_L g1635 ( 
.A(n_1537),
.B(n_1545),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1519),
.B(n_1535),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1439),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1515),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1535),
.B(n_1530),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1518),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1472),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1475),
.Y(n_1642)
);

BUFx12f_ASAP7_75t_L g1643 ( 
.A(n_1448),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1440),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1517),
.A2(n_1501),
.B(n_1449),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1445),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1446),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1538),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1522),
.Y(n_1649)
);

AOI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1465),
.A2(n_1500),
.B(n_1485),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1474),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1501),
.A2(n_1459),
.B(n_1588),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1555),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1480),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1548),
.B(n_1553),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1566),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1443),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_SL g1658 ( 
.A1(n_1457),
.A2(n_1444),
.B(n_1514),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1530),
.B(n_1484),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1503),
.B(n_1476),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1576),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1493),
.A2(n_1492),
.B(n_1511),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1581),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1522),
.A2(n_1469),
.B1(n_1591),
.B2(n_1456),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1511),
.B(n_1514),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1536),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_SL g1667 ( 
.A(n_1543),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1551),
.B(n_1587),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1443),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1520),
.A2(n_1486),
.B(n_1463),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1580),
.B(n_1583),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1551),
.Y(n_1673)
);

AO31x2_ASAP7_75t_L g1674 ( 
.A1(n_1524),
.A2(n_1602),
.A3(n_1595),
.B(n_1593),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1592),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1520),
.A2(n_1463),
.B(n_1466),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1548),
.A2(n_1567),
.B1(n_1598),
.B2(n_1554),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1551),
.B(n_1476),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1466),
.A2(n_1598),
.B(n_1526),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1470),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1591),
.Y(n_1682)
);

BUFx5_ASAP7_75t_L g1683 ( 
.A(n_1508),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1483),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1491),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1550),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1496),
.B(n_1473),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1462),
.A2(n_1486),
.B(n_1468),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1504),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1506),
.Y(n_1690)
);

AO21x1_ASAP7_75t_SL g1691 ( 
.A1(n_1477),
.A2(n_1490),
.B(n_1572),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1481),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1479),
.Y(n_1693)
);

AOI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1451),
.A2(n_1560),
.B(n_1507),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1512),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1573),
.A2(n_1547),
.B(n_1489),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1489),
.A2(n_1572),
.B(n_1582),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1490),
.Y(n_1698)
);

BUFx8_ASAP7_75t_L g1699 ( 
.A(n_1508),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1455),
.B(n_1596),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1447),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1447),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1564),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1564),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1510),
.A2(n_1596),
.B(n_1575),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1575),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1497),
.A2(n_1502),
.B(n_1442),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1478),
.A2(n_1453),
.B1(n_1590),
.B2(n_1543),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1494),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1453),
.B(n_1542),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1542),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1578),
.Y(n_1712)
);

AO21x1_ASAP7_75t_L g1713 ( 
.A1(n_1502),
.A2(n_1599),
.B(n_1594),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1488),
.B(n_1498),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1550),
.B(n_1574),
.Y(n_1715)
);

BUFx2_ASAP7_75t_SL g1716 ( 
.A(n_1436),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1574),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1574),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1487),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1570),
.B(n_1590),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1460),
.B(n_1495),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1482),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1482),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1478),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1499),
.Y(n_1725)
);

BUFx12f_ASAP7_75t_L g1726 ( 
.A(n_1643),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1618),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1610),
.A2(n_1464),
.B(n_1601),
.C(n_1541),
.Y(n_1728)
);

AND2x4_ASAP7_75t_SL g1729 ( 
.A(n_1679),
.B(n_1556),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1644),
.Y(n_1730)
);

AND2x2_ASAP7_75t_SL g1731 ( 
.A(n_1680),
.B(n_1544),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1635),
.A2(n_1577),
.B(n_1450),
.C(n_1549),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1678),
.B(n_1558),
.Y(n_1733)
);

BUFx4f_ASAP7_75t_L g1734 ( 
.A(n_1643),
.Y(n_1734)
);

INVxp33_ASAP7_75t_L g1735 ( 
.A(n_1693),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1672),
.B(n_1571),
.Y(n_1737)
);

AND2x4_ASAP7_75t_SL g1738 ( 
.A(n_1679),
.B(n_1448),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1644),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1613),
.A2(n_1549),
.B(n_1471),
.C(n_1467),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1617),
.B(n_1563),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1628),
.A2(n_1467),
.B(n_1563),
.C(n_1603),
.Y(n_1742)
);

AO21x1_ASAP7_75t_L g1743 ( 
.A1(n_1655),
.A2(n_1603),
.B(n_1604),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1669),
.B(n_1646),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1658),
.A2(n_1624),
.B(n_1677),
.C(n_1668),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1636),
.B(n_1631),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_SL g1747 ( 
.A1(n_1664),
.A2(n_1708),
.B1(n_1620),
.B2(n_1632),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1640),
.B(n_1671),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1658),
.A2(n_1605),
.B(n_1668),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1619),
.A2(n_1654),
.B(n_1645),
.C(n_1680),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1662),
.A2(n_1671),
.B(n_1633),
.C(n_1659),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1716),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1669),
.B(n_1647),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1662),
.A2(n_1633),
.B(n_1659),
.C(n_1614),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1698),
.B(n_1692),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1641),
.B(n_1651),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1666),
.B(n_1685),
.Y(n_1758)
);

NOR2xp67_ASAP7_75t_SL g1759 ( 
.A(n_1721),
.B(n_1725),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1680),
.A2(n_1650),
.B(n_1688),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1614),
.A2(n_1665),
.B(n_1640),
.C(n_1626),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1645),
.A2(n_1639),
.B1(n_1638),
.B2(n_1652),
.C(n_1690),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1648),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1615),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1688),
.A2(n_1705),
.B(n_1660),
.Y(n_1766)
);

A2O1A1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1665),
.A2(n_1639),
.B(n_1649),
.C(n_1638),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1623),
.A2(n_1607),
.B(n_1612),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1653),
.B(n_1656),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1653),
.B(n_1656),
.Y(n_1770)
);

A2O1A1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1649),
.A2(n_1705),
.B(n_1690),
.C(n_1611),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1661),
.B(n_1663),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1689),
.B(n_1691),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_L g1774 ( 
.A(n_1642),
.B(n_1683),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1689),
.B(n_1687),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1687),
.B(n_1606),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1688),
.A2(n_1676),
.B1(n_1700),
.B2(n_1724),
.Y(n_1777)
);

AO22x2_ASAP7_75t_L g1778 ( 
.A1(n_1615),
.A2(n_1612),
.B1(n_1611),
.B2(n_1608),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1709),
.A2(n_1724),
.B(n_1720),
.C(n_1706),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1649),
.A2(n_1630),
.B(n_1629),
.C(n_1676),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1688),
.B(n_1649),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1694),
.B(n_1652),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1701),
.A2(n_1702),
.B1(n_1704),
.B2(n_1703),
.C(n_1706),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_SL g1784 ( 
.A(n_1725),
.B(n_1721),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1676),
.A2(n_1700),
.B1(n_1716),
.B2(n_1719),
.Y(n_1785)
);

BUFx12f_ASAP7_75t_L g1786 ( 
.A(n_1723),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1629),
.A2(n_1630),
.B(n_1676),
.C(n_1608),
.Y(n_1787)
);

AO32x2_ASAP7_75t_L g1788 ( 
.A1(n_1622),
.A2(n_1673),
.A3(n_1670),
.B1(n_1686),
.B2(n_1657),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1704),
.A2(n_1695),
.B(n_1718),
.C(n_1710),
.Y(n_1789)
);

CKINVDCx14_ASAP7_75t_R g1790 ( 
.A(n_1714),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1629),
.A2(n_1630),
.B(n_1697),
.C(n_1707),
.Y(n_1791)
);

OA21x2_ASAP7_75t_L g1792 ( 
.A1(n_1607),
.A2(n_1681),
.B(n_1675),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1660),
.A2(n_1697),
.B(n_1696),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1667),
.A2(n_1609),
.B1(n_1723),
.B2(n_1722),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1731),
.A2(n_1609),
.B1(n_1714),
.B2(n_1699),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1775),
.B(n_1621),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1769),
.B(n_1621),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1731),
.A2(n_1749),
.B1(n_1790),
.B2(n_1760),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1792),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1792),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1792),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1769),
.B(n_1621),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1744),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1769),
.B(n_1621),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1788),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1753),
.B(n_1674),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1753),
.B(n_1621),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1727),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1730),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1739),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1747),
.A2(n_1722),
.B1(n_1609),
.B2(n_1699),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1765),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1748),
.B(n_1751),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1765),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1771),
.B(n_1616),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1770),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1616),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1781),
.B(n_1625),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1779),
.B(n_1712),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1743),
.A2(n_1609),
.B1(n_1699),
.B2(n_1700),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1770),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1791),
.B(n_1793),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1754),
.B(n_1616),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1738),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1764),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1764),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1754),
.B(n_1684),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1746),
.B(n_1711),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1756),
.B(n_1757),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1780),
.B(n_1673),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1816),
.B(n_1785),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1787),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1787),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1816),
.B(n_1788),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1812),
.Y(n_1836)
);

AOI222xp33_ASAP7_75t_L g1837 ( 
.A1(n_1811),
.A2(n_1745),
.B1(n_1742),
.B2(n_1763),
.C1(n_1761),
.C2(n_1760),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1798),
.A2(n_1745),
.B1(n_1742),
.B2(n_1784),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1826),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1808),
.Y(n_1840)
);

INVxp67_ASAP7_75t_SL g1841 ( 
.A(n_1819),
.Y(n_1841)
);

INVxp67_ASAP7_75t_SL g1842 ( 
.A(n_1819),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1798),
.A2(n_1750),
.B1(n_1762),
.B2(n_1782),
.C(n_1789),
.Y(n_1843)
);

OAI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1811),
.A2(n_1732),
.B1(n_1728),
.B2(n_1740),
.C(n_1762),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1803),
.B(n_1788),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1825),
.A2(n_1780),
.B(n_1767),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1795),
.A2(n_1790),
.B1(n_1726),
.B2(n_1752),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1831),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1795),
.A2(n_1728),
.B(n_1732),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1830),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1812),
.Y(n_1851)
);

OR2x6_ASAP7_75t_L g1852 ( 
.A(n_1815),
.B(n_1766),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1830),
.B(n_1735),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1820),
.A2(n_1771),
.B(n_1782),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1820),
.A2(n_1759),
.B1(n_1777),
.B2(n_1794),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1814),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1824),
.B(n_1783),
.C(n_1779),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1814),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1809),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1809),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1821),
.B(n_1778),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1800),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1817),
.B(n_1776),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1807),
.B(n_1778),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1810),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1825),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1810),
.Y(n_1867)
);

INVx5_ASAP7_75t_L g1868 ( 
.A(n_1831),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1823),
.A2(n_1735),
.B1(n_1767),
.B2(n_1758),
.C(n_1755),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1800),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1800),
.Y(n_1871)
);

INVxp67_ASAP7_75t_SL g1872 ( 
.A(n_1827),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1807),
.B(n_1778),
.Y(n_1873)
);

INVx4_ASAP7_75t_L g1874 ( 
.A(n_1825),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_SL g1875 ( 
.A(n_1824),
.B(n_1773),
.Y(n_1875)
);

INVx5_ASAP7_75t_SL g1876 ( 
.A(n_1831),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1802),
.B(n_1768),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1845),
.B(n_1805),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1859),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1860),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1838),
.A2(n_1815),
.B(n_1823),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1862),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1841),
.B(n_1842),
.Y(n_1883)
);

NAND2xp67_ASAP7_75t_L g1884 ( 
.A(n_1832),
.B(n_1738),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1805),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1835),
.B(n_1823),
.Y(n_1886)
);

INVx3_ASAP7_75t_SL g1887 ( 
.A(n_1852),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1835),
.B(n_1823),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1877),
.B(n_1799),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1865),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1868),
.B(n_1817),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1839),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1868),
.B(n_1817),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1868),
.B(n_1813),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1867),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1866),
.Y(n_1896)
);

OR2x6_ASAP7_75t_L g1897 ( 
.A(n_1846),
.B(n_1852),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1862),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1877),
.B(n_1799),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1836),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1847),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1857),
.Y(n_1902)
);

NAND2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1868),
.B(n_1831),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1875),
.B(n_1806),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1850),
.B(n_1818),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1875),
.B(n_1806),
.Y(n_1906)
);

INVx6_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1848),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1866),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1864),
.B(n_1873),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1851),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1870),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1870),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1848),
.B(n_1817),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1856),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1858),
.B(n_1818),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1833),
.B(n_1801),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1864),
.B(n_1813),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_L g1919 ( 
.A(n_1846),
.B(n_1825),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1873),
.B(n_1822),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1840),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_L g1922 ( 
.A(n_1843),
.B(n_1854),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1840),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1871),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1917),
.B(n_1833),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1883),
.B(n_1905),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1879),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1883),
.B(n_1853),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1902),
.B(n_1869),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1902),
.B(n_1834),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1905),
.B(n_1834),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1879),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1894),
.B(n_1848),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1880),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1892),
.B(n_1802),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1922),
.B(n_1863),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1881),
.B(n_1863),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1892),
.B(n_1804),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1880),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1881),
.B(n_1863),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1890),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_L g1942 ( 
.A(n_1901),
.B(n_1844),
.C(n_1849),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1897),
.A2(n_1837),
.B1(n_1852),
.B2(n_1855),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1890),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1907),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1895),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1897),
.A2(n_1852),
.B1(n_1828),
.B2(n_1741),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1916),
.B(n_1910),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1916),
.B(n_1861),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1900),
.B(n_1861),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1897),
.B(n_1876),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1882),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1895),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1900),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1896),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1897),
.A2(n_1848),
.B1(n_1876),
.B2(n_1832),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1911),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1882),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1911),
.B(n_1915),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1915),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1918),
.B(n_1829),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1921),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1897),
.B(n_1876),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1910),
.B(n_1804),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1882),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1910),
.B(n_1796),
.Y(n_1966)
);

NOR2x1_ASAP7_75t_L g1967 ( 
.A(n_1919),
.B(n_1874),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1898),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1921),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1917),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1918),
.B(n_1829),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1898),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1918),
.B(n_1822),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1919),
.B(n_1848),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1923),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1898),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1951),
.B(n_1897),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1925),
.B(n_1917),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1929),
.B(n_1886),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1951),
.B(n_1887),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1930),
.B(n_1955),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1970),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1970),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1952),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1942),
.A2(n_1887),
.B1(n_1914),
.B2(n_1891),
.Y(n_1985)
);

NOR2xp67_ASAP7_75t_SL g1986 ( 
.A(n_1974),
.B(n_1726),
.Y(n_1986)
);

AND2x2_ASAP7_75t_SL g1987 ( 
.A(n_1942),
.B(n_1734),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1927),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1932),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1963),
.B(n_1887),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1952),
.Y(n_1991)
);

INVx1_ASAP7_75t_SL g1992 ( 
.A(n_1936),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1925),
.B(n_1889),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1958),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1955),
.B(n_1886),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1948),
.B(n_1889),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1943),
.B(n_1886),
.Y(n_1997)
);

OAI21xp33_ASAP7_75t_L g1998 ( 
.A1(n_1947),
.A2(n_1884),
.B(n_1903),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1931),
.B(n_1889),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1963),
.B(n_1887),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1934),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1933),
.B(n_1904),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1947),
.B(n_1894),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1939),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1933),
.B(n_1904),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1941),
.Y(n_2006)
);

CKINVDCx16_ASAP7_75t_R g2007 ( 
.A(n_1967),
.Y(n_2007)
);

NAND3xp33_ASAP7_75t_L g2008 ( 
.A(n_1974),
.B(n_1899),
.C(n_1736),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1944),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1933),
.B(n_1904),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1928),
.B(n_1888),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1926),
.B(n_1899),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1937),
.B(n_1734),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1958),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1946),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1940),
.B(n_1884),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1945),
.B(n_1906),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1953),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_SL g2019 ( 
.A1(n_1985),
.A2(n_1956),
.B(n_1903),
.Y(n_2019)
);

OAI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_2007),
.A2(n_1903),
.B1(n_1907),
.B2(n_1945),
.Y(n_2020)
);

NAND4xp25_ASAP7_75t_L g2021 ( 
.A(n_1981),
.B(n_1733),
.C(n_1909),
.D(n_1896),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1998),
.A2(n_1907),
.B1(n_1891),
.B2(n_1893),
.Y(n_2022)
);

OAI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_2007),
.A2(n_1903),
.B1(n_1907),
.B2(n_1896),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1982),
.Y(n_2024)
);

AOI21xp33_ASAP7_75t_SL g2025 ( 
.A1(n_1987),
.A2(n_1908),
.B(n_1893),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_SL g2026 ( 
.A(n_2003),
.B(n_1884),
.Y(n_2026)
);

OAI322xp33_ASAP7_75t_SL g2027 ( 
.A1(n_1997),
.A2(n_1979),
.A3(n_1995),
.B1(n_1983),
.B2(n_1982),
.C1(n_2011),
.C2(n_2018),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1983),
.Y(n_2028)
);

OAI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1992),
.A2(n_2008),
.B1(n_1907),
.B2(n_2012),
.Y(n_2029)
);

A2O1A1Ixp33_ASAP7_75t_L g2030 ( 
.A1(n_1998),
.A2(n_1891),
.B(n_1893),
.C(n_1914),
.Y(n_2030)
);

CKINVDCx14_ASAP7_75t_R g2031 ( 
.A(n_2013),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1988),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1987),
.B(n_1786),
.Y(n_2033)
);

AOI211xp5_ASAP7_75t_L g2034 ( 
.A1(n_1986),
.A2(n_1891),
.B(n_1893),
.C(n_1909),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1987),
.A2(n_1907),
.B1(n_1891),
.B2(n_1893),
.Y(n_2035)
);

A2O1A1Ixp33_ASAP7_75t_SL g2036 ( 
.A1(n_1986),
.A2(n_1968),
.B(n_1972),
.C(n_1965),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_2016),
.A2(n_2008),
.B1(n_1977),
.B2(n_1990),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1988),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2002),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1989),
.B(n_1961),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1989),
.Y(n_2041)
);

OAI31xp33_ASAP7_75t_L g2042 ( 
.A1(n_1977),
.A2(n_1908),
.A3(n_1909),
.B(n_1914),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2001),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1980),
.A2(n_1876),
.B1(n_1906),
.B2(n_1914),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1980),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2001),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2004),
.Y(n_2047)
);

INVx1_ASAP7_75t_SL g2048 ( 
.A(n_1990),
.Y(n_2048)
);

A2O1A1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_2037),
.A2(n_2000),
.B(n_2012),
.C(n_2006),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2026),
.A2(n_2000),
.B1(n_2005),
.B2(n_2002),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2048),
.B(n_2004),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2024),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2029),
.B(n_1978),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2045),
.B(n_2005),
.Y(n_2054)
);

OAI32xp33_ASAP7_75t_L g2055 ( 
.A1(n_2037),
.A2(n_1978),
.A3(n_1999),
.B1(n_1993),
.B2(n_2017),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2039),
.B(n_2006),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_2028),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_2033),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2032),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2034),
.A2(n_1906),
.B1(n_1914),
.B2(n_2010),
.Y(n_2060)
);

INVxp67_ASAP7_75t_L g2061 ( 
.A(n_2021),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2029),
.A2(n_2009),
.B1(n_2018),
.B2(n_2015),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2038),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2031),
.B(n_2010),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2041),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2043),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2040),
.B(n_1999),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2046),
.Y(n_2068)
);

AND4x1_ASAP7_75t_L g2069 ( 
.A(n_2042),
.B(n_2017),
.C(n_2009),
.D(n_2015),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2047),
.B(n_1993),
.Y(n_2070)
);

INVxp67_ASAP7_75t_SL g2071 ( 
.A(n_2020),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2036),
.A2(n_1957),
.B(n_1954),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2064),
.B(n_2025),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2064),
.B(n_2019),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2057),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2057),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2054),
.B(n_2035),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2054),
.B(n_2022),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_2053),
.Y(n_2079)
);

OAI22xp33_ASAP7_75t_SL g2080 ( 
.A1(n_2053),
.A2(n_2071),
.B1(n_2061),
.B2(n_2050),
.Y(n_2080)
);

OAI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2062),
.A2(n_2030),
.B(n_2023),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2049),
.A2(n_2044),
.B1(n_2027),
.B2(n_1996),
.C(n_1908),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2062),
.A2(n_2049),
.B1(n_2058),
.B2(n_2060),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2051),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2055),
.A2(n_2023),
.B1(n_2020),
.B2(n_2014),
.C(n_1994),
.Y(n_2085)
);

O2A1O1Ixp33_ASAP7_75t_SL g2086 ( 
.A1(n_2072),
.A2(n_1996),
.B(n_1991),
.C(n_1994),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2070),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2079),
.B(n_2067),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2080),
.B(n_2052),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2083),
.A2(n_2056),
.B1(n_2063),
.B2(n_2059),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2081),
.A2(n_2068),
.B(n_2065),
.C(n_2066),
.Y(n_2091)
);

OAI21xp33_ASAP7_75t_SL g2092 ( 
.A1(n_2085),
.A2(n_2069),
.B(n_2014),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_2073),
.Y(n_2093)
);

NAND3xp33_ASAP7_75t_L g2094 ( 
.A(n_2086),
.B(n_2076),
.C(n_2075),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_2073),
.B(n_1984),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2078),
.B(n_2077),
.Y(n_2096)
);

NOR2x1_ASAP7_75t_L g2097 ( 
.A(n_2084),
.B(n_1991),
.Y(n_2097)
);

NOR3xp33_ASAP7_75t_L g2098 ( 
.A(n_2074),
.B(n_1984),
.C(n_1991),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2086),
.A2(n_1959),
.B(n_1960),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2092),
.A2(n_2082),
.B(n_2087),
.Y(n_2100)
);

NOR3xp33_ASAP7_75t_SL g2101 ( 
.A(n_2091),
.B(n_2076),
.C(n_1950),
.Y(n_2101)
);

OAI21xp33_ASAP7_75t_L g2102 ( 
.A1(n_2088),
.A2(n_1949),
.B(n_1965),
.Y(n_2102)
);

AOI221x1_ASAP7_75t_L g2103 ( 
.A1(n_2094),
.A2(n_1969),
.B1(n_1975),
.B2(n_1962),
.C(n_1976),
.Y(n_2103)
);

NOR4xp25_ASAP7_75t_L g2104 ( 
.A(n_2089),
.B(n_1976),
.C(n_1972),
.D(n_1968),
.Y(n_2104)
);

AOI211xp5_ASAP7_75t_L g2105 ( 
.A1(n_2093),
.A2(n_1715),
.B(n_1737),
.C(n_1686),
.Y(n_2105)
);

AND4x1_ASAP7_75t_L g2106 ( 
.A(n_2096),
.B(n_1715),
.C(n_1888),
.D(n_1699),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2090),
.A2(n_1938),
.B(n_1935),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2097),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_2101),
.B(n_2099),
.Y(n_2109)
);

OA211x2_ASAP7_75t_L g2110 ( 
.A1(n_2100),
.A2(n_2095),
.B(n_2098),
.C(n_1973),
.Y(n_2110)
);

NAND3xp33_ASAP7_75t_L g2111 ( 
.A(n_2103),
.B(n_1657),
.C(n_1627),
.Y(n_2111)
);

OAI211xp5_ASAP7_75t_SL g2112 ( 
.A1(n_2108),
.A2(n_1971),
.B(n_1627),
.C(n_1670),
.Y(n_2112)
);

OAI211xp5_ASAP7_75t_SL g2113 ( 
.A1(n_2102),
.A2(n_1964),
.B(n_1966),
.C(n_1786),
.Y(n_2113)
);

BUFx4f_ASAP7_75t_SL g2114 ( 
.A(n_2106),
.Y(n_2114)
);

OAI211xp5_ASAP7_75t_SL g2115 ( 
.A1(n_2105),
.A2(n_1774),
.B(n_1899),
.C(n_1923),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2107),
.Y(n_2116)
);

NAND4xp75_ASAP7_75t_L g2117 ( 
.A(n_2110),
.B(n_2109),
.C(n_2116),
.D(n_2114),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_2111),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2112),
.B(n_2104),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2113),
.Y(n_2120)
);

NOR3xp33_ASAP7_75t_L g2121 ( 
.A(n_2115),
.B(n_1874),
.C(n_1717),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_2109),
.B(n_1729),
.Y(n_2122)
);

AND3x4_ASAP7_75t_L g2123 ( 
.A(n_2121),
.B(n_1717),
.C(n_1700),
.Y(n_2123)
);

OAI221xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2118),
.A2(n_1888),
.B1(n_1717),
.B2(n_1878),
.C(n_1885),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2122),
.B(n_1920),
.Y(n_2125)
);

NAND4xp25_ASAP7_75t_L g2126 ( 
.A(n_2120),
.B(n_1874),
.C(n_1885),
.D(n_1878),
.Y(n_2126)
);

AOI321xp33_ASAP7_75t_L g2127 ( 
.A1(n_2124),
.A2(n_2119),
.A3(n_2117),
.B1(n_1878),
.B2(n_1885),
.C(n_1872),
.Y(n_2127)
);

OAI22x1_ASAP7_75t_L g2128 ( 
.A1(n_2127),
.A2(n_2123),
.B1(n_2125),
.B2(n_2126),
.Y(n_2128)
);

OAI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2128),
.A2(n_1920),
.B(n_1913),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2128),
.B(n_1729),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_2130),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_SL g2132 ( 
.A1(n_2129),
.A2(n_1682),
.B(n_1642),
.Y(n_2132)
);

AOI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_2131),
.A2(n_1913),
.B(n_1912),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_1912),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_2134),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2135),
.B(n_2133),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_2136),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2137),
.A2(n_1924),
.B1(n_1913),
.B2(n_1912),
.C(n_1920),
.Y(n_2138)
);

AOI211xp5_ASAP7_75t_L g2139 ( 
.A1(n_2138),
.A2(n_1682),
.B(n_1713),
.C(n_1774),
.Y(n_2139)
);


endmodule