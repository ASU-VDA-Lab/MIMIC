module fake_jpeg_22023_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_19),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx2_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_15),
.Y(n_69)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_36),
.B1(n_34),
.B2(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_67),
.B1(n_68),
.B2(n_16),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_73),
.B1(n_51),
.B2(n_39),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_55),
.B1(n_51),
.B2(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_36),
.B1(n_34),
.B2(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_25),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_90),
.B1(n_66),
.B2(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_47),
.A3(n_39),
.B1(n_40),
.B2(n_28),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_41),
.B(n_25),
.C(n_37),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_75),
.B1(n_71),
.B2(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_110),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_16),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_60),
.B1(n_56),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_114),
.B1(n_77),
.B2(n_58),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_94),
.A3(n_78),
.B1(n_72),
.B2(n_81),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_24),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_48),
.C(n_75),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_92),
.C(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_85),
.Y(n_109)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_57),
.B1(n_58),
.B2(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_69),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_120),
.B(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_135),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_141),
.B(n_142),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_130),
.C(n_107),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_131),
.B1(n_111),
.B2(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_79),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_79),
.C(n_86),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_86),
.B1(n_76),
.B2(n_67),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_24),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_141),
.B(n_142),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_105),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_84),
.B(n_87),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_112),
.B1(n_145),
.B2(n_110),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_166),
.B1(n_128),
.B2(n_134),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_106),
.B(n_116),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_120),
.B1(n_102),
.B2(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_165),
.B1(n_131),
.B2(n_124),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_169),
.C(n_41),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_120),
.C(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_111),
.B1(n_101),
.B2(n_115),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_171),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_63),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_83),
.C(n_71),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_63),
.A3(n_20),
.B1(n_24),
.B2(n_41),
.C1(n_43),
.C2(n_45),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_181),
.B1(n_192),
.B2(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_127),
.B1(n_130),
.B2(n_135),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_136),
.B1(n_126),
.B2(n_121),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_67),
.B1(n_83),
.B2(n_119),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_112),
.B1(n_84),
.B2(n_71),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_18),
.B1(n_14),
.B2(n_41),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_193),
.B1(n_154),
.B2(n_147),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_169),
.C(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_18),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_54),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_65),
.B1(n_14),
.B2(n_45),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_14),
.B1(n_65),
.B2(n_45),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_150),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_217),
.C(n_216),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_176),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_215),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_158),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_153),
.B1(n_167),
.B2(n_151),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_195),
.B1(n_177),
.B2(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_146),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_212),
.B(n_219),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_148),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_148),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_146),
.C(n_168),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_193),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_20),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_196),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_182),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_214),
.B1(n_175),
.B2(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_233),
.B1(n_22),
.B2(n_21),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_177),
.C(n_191),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_192),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_230),
.B(n_239),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_198),
.B1(n_194),
.B2(n_182),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_168),
.B1(n_27),
.B2(n_22),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_25),
.C(n_35),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_0),
.B(n_1),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_241),
.B(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_12),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_12),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_0),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_12),
.B(n_1),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_208),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_246),
.B(n_258),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_200),
.B(n_204),
.C(n_207),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_238),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_207),
.CI(n_25),
.CON(n_254),
.SN(n_254)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_0),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_221),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_25),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_229),
.B(n_226),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_270),
.B(n_2),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_232),
.C(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_25),
.C(n_3),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_266),
.Y(n_287)
);

NAND2x1_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_231),
.CI(n_21),
.CON(n_266),
.SN(n_266)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_0),
.B(n_2),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_245),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_247),
.B1(n_258),
.B2(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_243),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_276),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_253),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_288),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_267),
.C(n_262),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_2),
.B(n_3),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_269),
.B(n_264),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_287),
.B1(n_7),
.B2(n_9),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_300),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_294),
.B(n_296),
.Y(n_307)
);

AOI31xp67_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_266),
.A3(n_4),
.B(n_5),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_285),
.C(n_279),
.Y(n_296)
);

AOI31xp67_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_3),
.A3(n_5),
.B(n_6),
.Y(n_298)
);

AO22x1_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_5),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_6),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_6),
.B(n_7),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_297),
.B1(n_299),
.B2(n_10),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_7),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_311),
.A3(n_304),
.B1(n_11),
.B2(n_9),
.C1(n_35),
.C2(n_37),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_310),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_304),
.A3(n_11),
.B1(n_9),
.B2(n_35),
.C1(n_37),
.C2(n_31),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_11),
.B(n_31),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_11),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_31),
.B(n_283),
.Y(n_318)
);


endmodule