module fake_jpeg_27815_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_59),
.B1(n_60),
.B2(n_35),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_43),
.A2(n_19),
.B1(n_23),
.B2(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_17),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_27),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_16),
.B1(n_31),
.B2(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_70),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_72),
.B1(n_65),
.B2(n_76),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_38),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_82),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_79),
.Y(n_89)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_85),
.B1(n_87),
.B2(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_48),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_36),
.B1(n_34),
.B2(n_40),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_101),
.B(n_82),
.Y(n_118)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_57),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_103),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_37),
.B(n_1),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_108),
.B1(n_72),
.B2(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_51),
.B1(n_36),
.B2(n_34),
.Y(n_108)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_32),
.B1(n_61),
.B2(n_31),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_126),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_106),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_86),
.C(n_65),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_138),
.C(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_103),
.B1(n_98),
.B2(n_111),
.Y(n_162)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_87),
.B1(n_74),
.B2(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_132),
.B1(n_134),
.B2(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_37),
.B(n_74),
.C(n_56),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_127),
.B(n_121),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_75),
.B1(n_68),
.B2(n_79),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_28),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_95),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_69),
.B1(n_80),
.B2(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_136),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_89),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_81),
.C(n_49),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_91),
.B(n_108),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_49),
.C(n_58),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_44),
.B1(n_40),
.B2(n_61),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_101),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_145),
.B(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_153),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_155),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_125),
.B1(n_122),
.B2(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_125),
.B1(n_115),
.B2(n_129),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_92),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_98),
.B1(n_106),
.B2(n_105),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_114),
.B(n_106),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_105),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_164),
.B1(n_116),
.B2(n_23),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_11),
.C(n_13),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_13),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_23),
.B1(n_19),
.B2(n_111),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_28),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_168),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_112),
.B1(n_96),
.B2(n_91),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_28),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_137),
.B(n_126),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_96),
.B1(n_44),
.B2(n_61),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_22),
.B1(n_30),
.B2(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_24),
.B1(n_26),
.B2(n_168),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_177),
.B(n_193),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_58),
.C(n_38),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_39),
.C(n_26),
.Y(n_221)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_44),
.B1(n_26),
.B2(n_24),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_194),
.B1(n_197),
.B2(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_184),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_21),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_58),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_150),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_191),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_143),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_33),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_147),
.A2(n_154),
.B1(n_145),
.B2(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_165),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_216),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_218),
.B1(n_219),
.B2(n_222),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_154),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_223),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_28),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_181),
.C(n_188),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_227),
.C(n_241),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_193),
.C(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_197),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_186),
.B1(n_191),
.B2(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_200),
.B1(n_219),
.B2(n_199),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_174),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_184),
.C(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_198),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_189),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_239),
.CI(n_188),
.CON(n_249),
.SN(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_190),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_257),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_221),
.C(n_204),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_256),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_224),
.B1(n_226),
.B2(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_210),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_177),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_262),
.B1(n_268),
.B2(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_238),
.C(n_228),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_234),
.B1(n_218),
.B2(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_194),
.C(n_39),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_39),
.C(n_20),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_8),
.B(n_15),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_5),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_270),
.A2(n_251),
.B1(n_257),
.B2(n_247),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_12),
.B1(n_7),
.B2(n_2),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_276),
.B1(n_267),
.B2(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_245),
.C(n_39),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_264),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_282),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_6),
.B1(n_11),
.B2(n_9),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_5),
.C(n_11),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_279),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_4),
.C(n_6),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_4),
.C(n_7),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_12),
.B(n_1),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_289),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_2),
.B(n_291),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_280),
.C(n_281),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_2),
.C(n_0),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_1),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_299),
.B(n_292),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_304),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_298),
.B(n_300),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_307)
);


endmodule