module fake_jpeg_6948_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_46),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_9),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_27),
.B(n_32),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_72),
.Y(n_89)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_70),
.B1(n_31),
.B2(n_26),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_23),
.B1(n_17),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_28),
.B1(n_31),
.B2(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_62),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_24),
.B1(n_29),
.B2(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_81),
.B1(n_87),
.B2(n_19),
.Y(n_108)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_83),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_62),
.B1(n_47),
.B2(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_90),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_34),
.C(n_25),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_98),
.Y(n_124)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_60),
.B(n_61),
.Y(n_104)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_79),
.B1(n_31),
.B2(n_90),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_109),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_88),
.B1(n_87),
.B2(n_84),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_114),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_64),
.B(n_53),
.C(n_52),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_117),
.B1(n_47),
.B2(n_43),
.Y(n_137)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx2_ASAP7_75t_SL g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_61),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_97),
.B(n_84),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_49),
.B1(n_64),
.B2(n_68),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_59),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_122),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_63),
.A3(n_73),
.B1(n_20),
.B2(n_18),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_32),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_125),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_43),
.B1(n_37),
.B2(n_53),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_104),
.B1(n_128),
.B2(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_126),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_93),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_130),
.A2(n_148),
.B(n_25),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_143),
.B1(n_146),
.B2(n_151),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_134),
.B(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_91),
.B(n_25),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_140),
.B(n_122),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_54),
.B1(n_67),
.B2(n_47),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_80),
.B1(n_86),
.B2(n_103),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_123),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_152),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_40),
.B1(n_69),
.B2(n_74),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_71),
.B1(n_51),
.B2(n_79),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_156),
.B1(n_112),
.B2(n_118),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_20),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_80),
.C(n_75),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_125),
.C(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_112),
.B1(n_128),
.B2(n_119),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_141),
.B1(n_69),
.B2(n_27),
.Y(n_205)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_178),
.B1(n_129),
.B2(n_134),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_118),
.B(n_110),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_168),
.B(n_183),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_115),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_142),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_75),
.C(n_79),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_74),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_140),
.B1(n_143),
.B2(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_138),
.B(n_139),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_113),
.B1(n_69),
.B2(n_34),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_22),
.B1(n_27),
.B2(n_32),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_200),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_202),
.B(n_168),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_152),
.B1(n_133),
.B2(n_147),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_175),
.B1(n_176),
.B2(n_163),
.Y(n_223)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_203),
.C(n_182),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_129),
.B1(n_140),
.B2(n_142),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_162),
.B1(n_160),
.B2(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_22),
.A3(n_32),
.B1(n_27),
.B2(n_74),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_166),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_218),
.CI(n_213),
.CON(n_243),
.SN(n_243)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_172),
.B1(n_167),
.B2(n_181),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_217),
.A2(n_223),
.B1(n_235),
.B2(n_216),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_196),
.B1(n_200),
.B2(n_204),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_170),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_236),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_169),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_180),
.B(n_161),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_233),
.B(n_207),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_179),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_149),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_194),
.A2(n_185),
.B1(n_106),
.B2(n_22),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_27),
.C(n_149),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_185),
.C(n_153),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_153),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_202),
.C(n_199),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_194),
.B1(n_210),
.B2(n_197),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_221),
.B1(n_235),
.B2(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_234),
.B1(n_241),
.B2(n_4),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_197),
.B(n_209),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_250),
.B1(n_261),
.B2(n_1),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_199),
.C(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_196),
.C(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_1),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_8),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_215),
.A2(n_1),
.B(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_265),
.C(n_239),
.D(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_249),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_228),
.B(n_236),
.C(n_218),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_270),
.B1(n_282),
.B2(n_8),
.Y(n_299)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_252),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_3),
.C(n_4),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_283),
.C(n_251),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_281),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_259),
.B1(n_263),
.B2(n_244),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_253),
.Y(n_283)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_5),
.B(n_6),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_258),
.B1(n_6),
.B2(n_7),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_254),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_290),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_254),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_242),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_299),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_298),
.C(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_243),
.C(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_10),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_271),
.B1(n_284),
.B2(n_280),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_292),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_304),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_310),
.C(n_311),
.Y(n_324)
);

XOR2x1_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_269),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_283),
.C(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_270),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_269),
.B1(n_297),
.B2(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_316),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_290),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_269),
.B(n_11),
.C(n_12),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_320),
.B(n_14),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_10),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_11),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_12),
.B(n_13),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_305),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_306),
.B(n_301),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_326),
.C(n_317),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_318),
.B(n_329),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_305),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_330),
.B(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_15),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_333),
.A2(n_335),
.B(n_336),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_319),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_334),
.C(n_338),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_15),
.B(n_16),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_15),
.Y(n_344)
);


endmodule