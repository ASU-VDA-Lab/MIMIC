module fake_jpeg_24643_n_167 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_8),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_16),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_52),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_31),
.C(n_23),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_32),
.B2(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_68),
.B1(n_28),
.B2(n_25),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_26),
.B1(n_28),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_81),
.B1(n_83),
.B2(n_49),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_87),
.C(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_56),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_21),
.B1(n_36),
.B2(n_19),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_46),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_82),
.C(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_24),
.B1(n_27),
.B2(n_23),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_34),
.CI(n_19),
.CON(n_82),
.SN(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_29),
.B1(n_19),
.B2(n_5),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_64),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_99),
.B(n_100),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_47),
.B(n_52),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_110),
.B1(n_76),
.B2(n_96),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_88),
.B1(n_90),
.B2(n_84),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_57),
.C(n_51),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.C(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_51),
.C(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_79),
.B1(n_78),
.B2(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_116),
.B1(n_125),
.B2(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_79),
.B1(n_78),
.B2(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_120),
.C(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_69),
.C(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_19),
.Y(n_136)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_54),
.B1(n_89),
.B2(n_88),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_96),
.B1(n_95),
.B2(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_116),
.B1(n_125),
.B2(n_123),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_96),
.B(n_100),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_132),
.B(n_135),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_107),
.B(n_94),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_93),
.B(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_120),
.B1(n_123),
.B2(n_115),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_72),
.B(n_67),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_124),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_67),
.B(n_72),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_119),
.CI(n_118),
.CON(n_146),
.SN(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_148),
.C(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_115),
.C(n_118),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_134),
.A3(n_130),
.B1(n_139),
.B2(n_135),
.C1(n_132),
.C2(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_138),
.B1(n_145),
.B2(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_72),
.C(n_13),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_143),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_142),
.B1(n_4),
.B2(n_6),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_155),
.A3(n_159),
.B1(n_7),
.B2(n_8),
.C1(n_2),
.C2(n_12),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_2),
.B(n_4),
.C(n_9),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_2),
.A3(n_4),
.B1(n_7),
.B2(n_9),
.C1(n_12),
.C2(n_161),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_12),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_165),
.Y(n_167)
);


endmodule