module fake_jpeg_2736_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_44),
.B1(n_56),
.B2(n_53),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_54),
.B1(n_52),
.B2(n_43),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_44),
.B1(n_51),
.B2(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_56),
.B1(n_53),
.B2(n_48),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_57),
.C(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_58),
.B1(n_68),
.B2(n_51),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_74),
.C(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_8),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_87),
.B1(n_22),
.B2(n_23),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_68),
.B(n_61),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_47),
.B1(n_46),
.B2(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_104),
.B1(n_0),
.B2(n_1),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_85),
.C(n_78),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_28),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_46),
.C(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_29),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_108),
.B1(n_117),
.B2(n_123),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_121),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_105),
.B(n_11),
.Y(n_138)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_118),
.B(n_9),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_32),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_31),
.B1(n_38),
.B2(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_27),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_16),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_33),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_10),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_138),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_123),
.B(n_17),
.C(n_34),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_136),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_10),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_135),
.C(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_35),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_125),
.C(n_134),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_141),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_152),
.B1(n_140),
.B2(n_145),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_143),
.B(n_133),
.Y(n_158)
);

NAND4xp25_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_147),
.C(n_141),
.D(n_153),
.Y(n_157)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_158),
.B1(n_156),
.B2(n_36),
.C(n_39),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_11),
.C(n_12),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_14),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_14),
.Y(n_165)
);


endmodule