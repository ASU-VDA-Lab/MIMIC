module fake_ariane_394_n_107 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_107);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_107;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_R g38 ( 
.A(n_25),
.B(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_R g47 ( 
.A(n_28),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_R g48 ( 
.A(n_28),
.B(n_8),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_35),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_33),
.B1(n_20),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_56)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

BUFx4_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_45),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_50),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_48),
.C(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_55),
.B1(n_57),
.B2(n_63),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_68),
.B(n_65),
.Y(n_75)
);

AO31x2_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_64),
.A3(n_59),
.B(n_45),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_56),
.B1(n_55),
.B2(n_69),
.C(n_44),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_65),
.B(n_64),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_67),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_67),
.Y(n_84)
);

AO21x2_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_47),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_42),
.B(n_2),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_84),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_97),
.B(n_94),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_42),
.B1(n_85),
.B2(n_88),
.C(n_1),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_85),
.B1(n_49),
.B2(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI22x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_99),
.B1(n_7),
.B2(n_3),
.Y(n_104)
);

OAI211xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_7),
.C(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_49),
.B1(n_50),
.B2(n_73),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_49),
.B1(n_50),
.B2(n_9),
.C(n_73),
.Y(n_107)
);


endmodule