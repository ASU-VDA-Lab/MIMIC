module real_jpeg_724_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_1),
.B(n_62),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_164),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_1),
.A2(n_28),
.B(n_29),
.C(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_34),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_48),
.C(n_51),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_1),
.B(n_91),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_80),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_43),
.B1(n_62),
.B2(n_63),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_43),
.B1(n_51),
.B2(n_53),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_4),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_123),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_123),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_51),
.B1(n_53),
.B2(n_123),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_10),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_11),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_163),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_11),
.A2(n_51),
.B1(n_53),
.B2(n_163),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_65),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_13),
.A2(n_51),
.B1(n_53),
.B2(n_65),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_14),
.A2(n_40),
.B1(n_51),
.B2(n_53),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_15),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_101),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_15),
.A2(n_51),
.B1(n_53),
.B2(n_101),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_327),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_314),
.B(n_326),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_139),
.B(n_311),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_126),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_22),
.B(n_102),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_58),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_24),
.A2(n_25),
.B(n_44),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_24),
.B(n_58),
.C(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_44),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_26),
.A2(n_41),
.B1(n_42),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_26),
.A2(n_39),
.B1(n_41),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_26),
.A2(n_41),
.B1(n_77),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_26),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_26),
.A2(n_182),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_27),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_34),
.B1(n_181),
.B2(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_27),
.A2(n_34),
.B(n_318),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_30),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_29),
.A2(n_63),
.A3(n_69),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_30),
.B(n_71),
.Y(n_186)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_34),
.B(n_160),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_35),
.A2(n_38),
.B(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_36),
.B(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_41),
.A2(n_119),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_41),
.A2(n_159),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_50),
.B1(n_54),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_45),
.A2(n_50),
.B1(n_207),
.B2(n_241),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_45),
.A2(n_209),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_46),
.A2(n_80),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_46),
.A2(n_80),
.B1(n_117),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_46),
.A2(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_46),
.B(n_210),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_50),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_50),
.A2(n_230),
.B(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_51),
.B(n_270),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_82),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_60),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_60),
.B(n_75),
.C(n_79),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_60),
.B(n_130),
.C(n_137),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_68),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_66),
.B(n_214),
.C(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_66),
.A2(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_66),
.A2(n_68),
.B1(n_73),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_67),
.A2(n_122),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_67),
.A2(n_164),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_67),
.A2(n_164),
.B1(n_321),
.B2(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_68),
.A2(n_98),
.B(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_79),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_79),
.B(n_131),
.C(n_135),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_80),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_97),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_85),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_87),
.B1(n_97),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_88),
.A2(n_91),
.B1(n_114),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_88),
.A2(n_214),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_89),
.A2(n_90),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_89),
.A2(n_90),
.B1(n_189),
.B2(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_89),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_89),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_89),
.A2(n_90),
.B1(n_245),
.B2(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_90),
.A2(n_204),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_90),
.B(n_218),
.Y(n_247)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_91),
.A2(n_217),
.B(n_274),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_109),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.C(n_120),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_111),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_120),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_125),
.B(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_126),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_127),
.B(n_138),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_132),
.Y(n_320)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_136),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_165),
.B(n_310),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_141),
.B(n_144),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.C(n_161),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_152),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_153),
.B(n_155),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_191),
.B(n_309),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_167),
.B(n_169),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.C(n_176),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_170),
.B(n_174),
.Y(n_294)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_176),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_183),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_177),
.B(n_179),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_183),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI31xp33_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_291),
.A3(n_301),
.B(n_306),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_235),
.B(n_290),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_219),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_194),
.B(n_219),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.C(n_211),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_195),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_200),
.C(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_205),
.B(n_211),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_215),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_231),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_220),
.B(n_232),
.C(n_234),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_226),
.C(n_227),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_285),
.B(n_289),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_254),
.B(n_284),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_248),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_248),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_244),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_266),
.B(n_283),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_277),
.B(n_282),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B(n_276),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_280),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);


endmodule