module fake_netlist_1_12757_n_530 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_530);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_530;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_305;
wire n_100;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_59), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_7), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_9), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_68), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_8), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_39), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_69), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_47), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_48), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_32), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_56), .Y(n_88) );
BUFx2_ASAP7_75t_L g89 ( .A(n_42), .Y(n_89) );
NOR2xp33_ASAP7_75t_L g90 ( .A(n_52), .B(n_15), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_18), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_54), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_29), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_14), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_30), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_50), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_41), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_9), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_2), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_21), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_63), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
AND2x6_ASAP7_75t_L g117 ( .A(n_77), .B(n_37), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_89), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_89), .B(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_116), .Y(n_121) );
NAND2x1_ASAP7_75t_L g122 ( .A(n_81), .B(n_3), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_115), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_82), .B(n_4), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_84), .B(n_44), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
NAND2xp33_ASAP7_75t_SL g134 ( .A(n_107), .B(n_5), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
NAND2xp33_ASAP7_75t_L g139 ( .A(n_117), .B(n_88), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_124), .B(n_94), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_137), .B(n_83), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
NOR2xp67_ASAP7_75t_L g144 ( .A(n_120), .B(n_96), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_117), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_124), .B(n_94), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_123), .B(n_99), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_130), .B(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_130), .B(n_101), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_131), .B(n_113), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_121), .B(n_81), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_125), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_134), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_131), .B(n_101), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_133), .B(n_114), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_133), .B(n_104), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_138), .B(n_112), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_138), .B(n_111), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_161), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NAND3xp33_ASAP7_75t_L g165 ( .A(n_139), .B(n_127), .C(n_122), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_153), .B(n_117), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_155), .B(n_122), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_155), .B(n_117), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_145), .B(n_132), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_142), .B(n_119), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_158), .B(n_129), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_160), .B(n_128), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
CKINVDCx14_ASAP7_75t_R g177 ( .A(n_156), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g178 ( .A(n_154), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_154), .B(n_117), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_161), .B(n_118), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_148), .B(n_117), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_143), .Y(n_186) );
AND3x1_ASAP7_75t_SL g187 ( .A(n_144), .B(n_111), .C(n_98), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_150), .B(n_135), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_144), .B(n_135), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_149), .B(n_135), .Y(n_190) );
BUFx8_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_145), .B(n_102), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_149), .B(n_78), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_163), .B(n_185), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_163), .B(n_151), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_167), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_193), .B(n_151), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_181), .A2(n_157), .B1(n_150), .B2(n_140), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_164), .B(n_162), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_193), .B(n_146), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_193), .B(n_188), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_181), .A2(n_146), .B1(n_159), .B2(n_162), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_191), .B(n_162), .Y(n_208) );
BUFx4_ASAP7_75t_SL g209 ( .A(n_168), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_184), .A2(n_145), .B(n_162), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_168), .B(n_193), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_188), .B(n_145), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_173), .B(n_162), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_179), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_166), .A2(n_145), .B(n_162), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_174), .B(n_110), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_175), .B(n_98), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_181), .B(n_126), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_178), .B(n_95), .C(n_90), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_191), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_182), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_170), .A2(n_109), .B(n_108), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_223), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_207), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_207), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_199), .B(n_181), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_198), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_198), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_198), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_215), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_215), .Y(n_236) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_216), .A2(n_182), .B(n_172), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_218), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_199), .B(n_186), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_218), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_204), .B(n_186), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_214), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_224), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_214), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_210), .A2(n_180), .B(n_165), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_204), .B(n_194), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_224), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_205), .B(n_194), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_198), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_229), .B(n_211), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_239), .A2(n_196), .B1(n_202), .B2(n_249), .Y(n_255) );
AO21x1_ASAP7_75t_SL g256 ( .A1(n_248), .A2(n_206), .B(n_86), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_227), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_228), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_239), .B(n_200), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_229), .B(n_211), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_211), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_241), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_229), .B(n_221), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_236), .B(n_221), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_246), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_234), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_260), .Y(n_274) );
OR2x6_ASAP7_75t_L g275 ( .A(n_266), .B(n_223), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_259), .B(n_221), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_222), .B1(n_189), .B2(n_226), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_257), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_252), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_189), .B1(n_226), .B2(n_165), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_265), .A2(n_202), .B1(n_247), .B2(n_236), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_260), .B(n_231), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_273), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_273), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_271), .B(n_246), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_263), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_293), .B(n_258), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_281), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
AOI32xp33_ASAP7_75t_L g306 ( .A1(n_280), .A2(n_95), .A3(n_105), .B1(n_92), .B2(n_109), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_281), .B(n_233), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_291), .B(n_258), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_295), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_264), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_274), .B(n_264), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_274), .B(n_267), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_293), .B(n_267), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_289), .B(n_268), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_278), .B(n_268), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_289), .B(n_234), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_281), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_301), .B(n_294), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_302), .B(n_281), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_305), .B(n_275), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_317), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_310), .B(n_288), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_303), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_302), .B(n_284), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_299), .B(n_286), .Y(n_338) );
NAND3xp33_ASAP7_75t_SL g339 ( .A(n_306), .B(n_87), .C(n_92), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_304), .B(n_292), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_323), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_304), .B(n_292), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_318), .B(n_288), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_324), .B(n_288), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_319), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_320), .B(n_284), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_315), .B(n_284), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_310), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_322), .B(n_284), .Y(n_358) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_302), .B(n_284), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
NAND2xp33_ASAP7_75t_L g361 ( .A(n_323), .B(n_270), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_314), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_321), .B(n_87), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_307), .B(n_97), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_307), .B(n_275), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_307), .B(n_275), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_275), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_327), .B(n_6), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_357), .B(n_97), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_366), .A2(n_285), .B(n_100), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_350), .B(n_100), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_355), .B(n_270), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_351), .B(n_102), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_352), .B(n_103), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_358), .B(n_103), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_330), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_361), .A2(n_208), .B(n_244), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_327), .B(n_6), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_356), .B(n_105), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_360), .B(n_108), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_331), .B(n_8), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_338), .B(n_10), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_362), .B(n_189), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_366), .A2(n_272), .B(n_206), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_358), .B(n_10), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_343), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_340), .B(n_245), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_11), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_348), .B(n_217), .C(n_219), .D(n_189), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_364), .B(n_11), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_336), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_359), .B(n_226), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_329), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_340), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_364), .B(n_12), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_347), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_326), .B(n_226), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_344), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_332), .B(n_12), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_363), .B(n_325), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_325), .B(n_13), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_346), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_365), .B(n_243), .C(n_238), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_353), .A2(n_231), .B(n_250), .Y(n_411) );
OAI21xp33_ASAP7_75t_SL g412 ( .A1(n_344), .A2(n_232), .B(n_231), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_346), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_361), .B(n_233), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_349), .B(n_14), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_335), .B(n_16), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_354), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_333), .B(n_245), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_386), .B(n_339), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_371), .A2(n_337), .B(n_326), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_405), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_395), .A2(n_337), .B(n_326), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_386), .B(n_367), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_SL g426 ( .A1(n_406), .A2(n_177), .B(n_233), .C(n_238), .Y(n_426) );
NAND4xp75_ASAP7_75t_L g427 ( .A(n_412), .B(n_269), .C(n_262), .D(n_232), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_369), .B(n_337), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_379), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_385), .A2(n_253), .B(n_240), .C(n_243), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
NAND5xp2_ASAP7_75t_L g432 ( .A(n_369), .B(n_262), .C(n_209), .D(n_240), .E(n_247), .Y(n_432) );
NAND3xp33_ASAP7_75t_SL g433 ( .A(n_416), .B(n_248), .C(n_251), .Y(n_433) );
NOR2xp67_ASAP7_75t_L g434 ( .A(n_410), .B(n_16), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_377), .B(n_17), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_385), .B(n_244), .C(n_251), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_416), .B(n_244), .C(n_251), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_381), .B(n_17), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_406), .A2(n_225), .B1(n_190), .B2(n_187), .C(n_250), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g440 ( .A1(n_381), .A2(n_250), .B(n_232), .C(n_233), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_407), .B(n_245), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_400), .B(n_251), .Y(n_442) );
AND3x1_ASAP7_75t_L g443 ( .A(n_394), .B(n_233), .C(n_244), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_382), .A2(n_242), .B1(n_230), .B2(n_249), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_384), .A2(n_201), .B(n_230), .C(n_242), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_400), .B(n_19), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_408), .B(n_396), .C(n_402), .D(n_368), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_409), .B(n_242), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_417), .B(n_20), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_390), .B(n_22), .Y(n_450) );
AOI221x1_ASAP7_75t_L g451 ( .A1(n_372), .A2(n_230), .B1(n_213), .B2(n_195), .C(n_176), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_392), .Y(n_452) );
OA22x2_ASAP7_75t_L g453 ( .A1(n_404), .A2(n_212), .B1(n_25), .B2(n_27), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
OAI21xp33_ASAP7_75t_SL g455 ( .A1(n_404), .A2(n_212), .B(n_194), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_413), .B(n_237), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_415), .B(n_192), .C(n_176), .D(n_183), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_375), .B(n_198), .C(n_195), .Y(n_459) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_398), .B(n_23), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_376), .B(n_198), .C(n_195), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_383), .B(n_237), .C(n_176), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_425), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_443), .B(n_414), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_434), .A2(n_391), .B(n_380), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_421), .A2(n_417), .B1(n_374), .B2(n_398), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_422), .B(n_418), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_445), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_453), .A2(n_411), .B(n_370), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_453), .A2(n_389), .B(n_387), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_455), .A2(n_373), .B(n_397), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_447), .B(n_399), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_424), .B(n_418), .C(n_397), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_432), .A2(n_393), .B(n_195), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_422), .B(n_393), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
AND3x2_ASAP7_75t_L g478 ( .A(n_438), .B(n_419), .C(n_428), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_432), .A2(n_195), .B(n_183), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_440), .B(n_203), .C(n_183), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_420), .Y(n_481) );
NOR4xp75_ASAP7_75t_L g482 ( .A(n_427), .B(n_237), .C(n_33), .D(n_40), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_452), .B(n_31), .Y(n_483) );
XOR2xp5_ASAP7_75t_L g484 ( .A(n_437), .B(n_43), .Y(n_484) );
OAI322xp33_ASAP7_75t_L g485 ( .A1(n_454), .A2(n_171), .A3(n_203), .B1(n_51), .B2(n_53), .C1(n_57), .C2(n_58), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_457), .B(n_45), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_436), .B(n_191), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_423), .B(n_191), .C(n_171), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_441), .B(n_46), .Y(n_489) );
XOR2xp5_ASAP7_75t_L g490 ( .A(n_435), .B(n_60), .Y(n_490) );
NOR3xp33_ASAP7_75t_SL g491 ( .A(n_433), .B(n_61), .C(n_62), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_426), .A2(n_430), .B(n_461), .C(n_459), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_467), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_473), .B(n_449), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_466), .B(n_460), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_476), .B(n_442), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_468), .B(n_448), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_468), .A2(n_439), .B1(n_458), .B2(n_444), .C(n_450), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_473), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_474), .B(n_446), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
NOR2xp33_ASAP7_75t_R g502 ( .A(n_478), .B(n_64), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_469), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_471), .A2(n_462), .B1(n_456), .B2(n_451), .C(n_203), .Y(n_504) );
NAND3x1_ASAP7_75t_L g505 ( .A(n_465), .B(n_65), .C(n_66), .Y(n_505) );
AOI31xp33_ASAP7_75t_L g506 ( .A1(n_488), .A2(n_67), .A3(n_70), .B(n_71), .Y(n_506) );
XOR2xp5_ASAP7_75t_L g507 ( .A(n_490), .B(n_73), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_481), .B(n_74), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_464), .B(n_75), .Y(n_509) );
OAI321xp33_ASAP7_75t_L g510 ( .A1(n_495), .A2(n_470), .A3(n_480), .B1(n_472), .B2(n_478), .C(n_487), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_497), .B(n_477), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_499), .A2(n_491), .B1(n_484), .B2(n_475), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_507), .Y(n_513) );
NAND2x1_ASAP7_75t_L g514 ( .A(n_493), .B(n_491), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g515 ( .A1(n_502), .A2(n_492), .B(n_485), .C(n_489), .Y(n_515) );
NOR2xp67_ASAP7_75t_SL g516 ( .A(n_504), .B(n_479), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_497), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_501), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_517), .B(n_498), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_516), .A2(n_498), .B1(n_504), .B2(n_503), .C(n_506), .Y(n_520) );
OAI211xp5_ASAP7_75t_SL g521 ( .A1(n_515), .A2(n_508), .B(n_486), .C(n_496), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_514), .A2(n_494), .B1(n_500), .B2(n_505), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_512), .A2(n_509), .B1(n_483), .B2(n_482), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_522), .A2(n_517), .B1(n_511), .B2(n_518), .Y(n_524) );
NOR3xp33_ASAP7_75t_L g525 ( .A(n_520), .B(n_510), .C(n_509), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_519), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_526), .B(n_523), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_525), .A2(n_521), .B1(n_513), .B2(n_76), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_527), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_529), .A2(n_524), .B(n_528), .Y(n_530) );
endmodule