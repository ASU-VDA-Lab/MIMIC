module real_jpeg_2940_n_6 (n_5, n_4, n_36, n_0, n_39, n_37, n_1, n_2, n_35, n_38, n_3, n_6);

input n_5;
input n_4;
input n_36;
input n_0;
input n_39;
input n_37;
input n_1;
input n_2;
input n_35;
input n_38;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_1),
.A2(n_21),
.B(n_25),
.Y(n_20)
);

AO22x1_ASAP7_75t_L g16 ( 
.A1(n_2),
.A2(n_17),
.B1(n_19),
.B2(n_30),
.Y(n_16)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_16),
.C(n_31),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_4),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_14),
.Y(n_6)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_18),
.Y(n_17)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.C(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_35),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_36),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_37),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_38),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_39),
.Y(n_32)
);


endmodule