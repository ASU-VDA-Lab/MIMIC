module fake_jpeg_374_n_225 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_225);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_24),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_66),
.B1(n_63),
.B2(n_73),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_98),
.B1(n_76),
.B2(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_72),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_66),
.B1(n_80),
.B2(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_77),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_70),
.B1(n_77),
.B2(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_88),
.B1(n_86),
.B2(n_59),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_74),
.B1(n_64),
.B2(n_76),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_116),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_120),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_131),
.B1(n_142),
.B2(n_134),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_81),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_127),
.B(n_9),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_136),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_61),
.B(n_81),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_64),
.B1(n_74),
.B2(n_61),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_68),
.B1(n_58),
.B2(n_54),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_65),
.B1(n_25),
.B2(n_27),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_0),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_0),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_28),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_1),
.C(n_2),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_9),
.C(n_10),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_79),
.B1(n_65),
.B2(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_2),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_3),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_4),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_65),
.B1(n_30),
.B2(n_31),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_19),
.B(n_50),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_53),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_163),
.B(n_165),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_8),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_160),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_138),
.C(n_34),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_175),
.C(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_16),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_35),
.B(n_45),
.Y(n_178)
);

OA21x2_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_41),
.B(n_48),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_32),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_152),
.C(n_154),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_44),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_36),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_198),
.C(n_184),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_17),
.B1(n_21),
.B2(n_39),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_173),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_175),
.B(n_168),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_205),
.C(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_180),
.B1(n_172),
.B2(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_213),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_181),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_198),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_218),
.C(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_206),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_221),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_214),
.A3(n_186),
.B1(n_212),
.B2(n_200),
.C(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_190),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_170),
.C(n_199),
.Y(n_225)
);


endmodule