module fake_jpeg_7900_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_1),
.B(n_4),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_30),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_14),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_12),
.B1(n_22),
.B2(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_30),
.B1(n_18),
.B2(n_21),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_16),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_26),
.C(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_25),
.Y(n_47)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_28),
.B1(n_24),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_42),
.B1(n_28),
.B2(n_52),
.Y(n_56)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_1),
.Y(n_45)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_5),
.Y(n_57)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_11),
.B1(n_30),
.B2(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_57),
.B1(n_62),
.B2(n_11),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_38),
.B1(n_23),
.B2(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_49),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_73),
.B(n_74),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_34),
.C(n_31),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_39),
.B(n_38),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_45),
.B(n_34),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_64),
.B1(n_46),
.B2(n_17),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_57),
.C(n_58),
.Y(n_76)
);

OAI322xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_82),
.A3(n_17),
.B1(n_29),
.B2(n_8),
.C1(n_9),
.C2(n_6),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_61),
.B(n_63),
.C(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_60),
.B(n_14),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_75),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_27),
.B(n_29),
.C(n_23),
.D(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_16),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_74),
.C(n_73),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_93),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_81),
.Y(n_98)
);

NOR4xp25_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_3),
.C(n_29),
.D(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_89),
.C(n_91),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_90),
.B(n_9),
.C(n_3),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_98),
.B(n_102),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);


endmodule