module real_aes_1154_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_758, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_759, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_758;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_759;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g163 ( .A(n_0), .B(n_137), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_1), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_2), .B(n_121), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_3), .B(n_139), .Y(n_450) );
INVx1_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_5), .B(n_121), .Y(n_190) );
NAND2xp33_ASAP7_75t_SL g233 ( .A(n_6), .B(n_127), .Y(n_233) );
INVx1_ASAP7_75t_L g225 ( .A(n_7), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_8), .Y(n_732) );
AND2x2_ASAP7_75t_L g188 ( .A(n_9), .B(n_145), .Y(n_188) );
AND2x2_ASAP7_75t_L g452 ( .A(n_10), .B(n_141), .Y(n_452) );
AND2x2_ASAP7_75t_L g462 ( .A(n_11), .B(n_231), .Y(n_462) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_13), .B(n_139), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
AOI221x1_ASAP7_75t_L g228 ( .A1(n_15), .A2(n_130), .B1(n_229), .B2(n_231), .C(n_232), .Y(n_228) );
AOI22xp5_ASAP7_75t_SL g715 ( .A1(n_16), .A2(n_73), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_16), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_17), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_18), .B(n_121), .Y(n_507) );
INVx1_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_20), .A2(n_89), .B1(n_121), .B2(n_174), .Y(n_466) );
AOI221xp5_ASAP7_75t_SL g152 ( .A1(n_21), .A2(n_37), .B1(n_121), .B2(n_130), .C(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_22), .A2(n_130), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_23), .B(n_137), .Y(n_193) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_24), .A2(n_88), .B(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g146 ( .A(n_24), .B(n_88), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_25), .B(n_139), .Y(n_138) );
INVxp67_ASAP7_75t_L g227 ( .A(n_26), .Y(n_227) );
AND2x2_ASAP7_75t_L g214 ( .A(n_27), .B(n_151), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_28), .A2(n_130), .B(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_29), .A2(n_231), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_30), .B(n_139), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_31), .A2(n_70), .B1(n_742), .B2(n_743), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_31), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_32), .B(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_33), .A2(n_130), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_34), .B(n_139), .Y(n_522) );
AND2x2_ASAP7_75t_L g127 ( .A(n_35), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g131 ( .A(n_35), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g182 ( .A(n_35), .Y(n_182) );
OR2x6_ASAP7_75t_L g109 ( .A(n_36), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_38), .B(n_121), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_39), .A2(n_81), .B1(n_130), .B2(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_40), .B(n_139), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_41), .B(n_121), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_42), .B(n_137), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_43), .A2(n_130), .B(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_44), .A2(n_715), .B1(n_719), .B2(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g166 ( .A(n_45), .B(n_151), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_46), .B(n_137), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_47), .B(n_151), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_48), .B(n_121), .Y(n_499) );
INVx1_ASAP7_75t_L g124 ( .A(n_49), .Y(n_124) );
INVx1_ASAP7_75t_L g134 ( .A(n_49), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_50), .B(n_139), .Y(n_460) );
AND2x2_ASAP7_75t_L g489 ( .A(n_51), .B(n_151), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_52), .B(n_121), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_53), .B(n_137), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_54), .B(n_137), .Y(n_521) );
AND2x2_ASAP7_75t_L g205 ( .A(n_55), .B(n_151), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_56), .B(n_121), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_57), .B(n_139), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_58), .B(n_121), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_59), .A2(n_130), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_60), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_61), .B(n_137), .Y(n_202) );
AND2x2_ASAP7_75t_L g513 ( .A(n_62), .B(n_145), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_63), .A2(n_130), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_64), .B(n_139), .Y(n_194) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_65), .B(n_141), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_66), .B(n_137), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_67), .B(n_137), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_68), .A2(n_91), .B1(n_130), .B2(n_180), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_69), .B(n_139), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_70), .A2(n_101), .B1(n_725), .B2(n_736), .C1(n_746), .C2(n_750), .Y(n_100) );
INVx1_ASAP7_75t_L g742 ( .A(n_70), .Y(n_742) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_71), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_72), .B(n_137), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_73), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_74), .A2(n_130), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_75), .A2(n_130), .B(n_440), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_76), .A2(n_130), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g524 ( .A(n_77), .B(n_145), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_78), .B(n_151), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_79), .A2(n_83), .B1(n_121), .B2(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_80), .B(n_121), .Y(n_203) );
INVx1_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_84), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_85), .B(n_137), .Y(n_155) );
AND2x2_ASAP7_75t_L g443 ( .A(n_86), .B(n_141), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_87), .A2(n_130), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_90), .B(n_139), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_92), .A2(n_130), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_93), .B(n_139), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_94), .B(n_121), .Y(n_165) );
INVxp67_ASAP7_75t_L g230 ( .A(n_95), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_96), .B(n_139), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_97), .A2(n_130), .B(n_135), .Y(n_129) );
BUFx2_ASAP7_75t_L g512 ( .A(n_98), .Y(n_512) );
BUFx2_ASAP7_75t_L g733 ( .A(n_99), .Y(n_733) );
BUFx2_ASAP7_75t_SL g754 ( .A(n_99), .Y(n_754) );
OAI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_715), .B(n_718), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_113), .B1(n_427), .B2(n_711), .Y(n_103) );
INVx4_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx3_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_SL g720 ( .A1(n_107), .A2(n_113), .B1(n_427), .B2(n_712), .Y(n_720) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_SL g713 ( .A(n_108), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g724 ( .A(n_108), .B(n_109), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_108), .B(n_714), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_109), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
XNOR2xp5_ASAP7_75t_L g740 ( .A(n_113), .B(n_741), .Y(n_740) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_319), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_247), .C(n_297), .Y(n_114) );
OAI211xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_167), .B(n_215), .C(n_236), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_147), .Y(n_116) );
AND2x2_ASAP7_75t_L g246 ( .A(n_117), .B(n_148), .Y(n_246) );
INVx1_ASAP7_75t_L g377 ( .A(n_117), .Y(n_377) );
NOR2x1p5_ASAP7_75t_L g409 ( .A(n_117), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g220 ( .A(n_118), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g268 ( .A(n_118), .Y(n_268) );
OR2x2_ASAP7_75t_L g272 ( .A(n_118), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_118), .B(n_150), .Y(n_284) );
OR2x2_ASAP7_75t_L g306 ( .A(n_118), .B(n_150), .Y(n_306) );
AND2x4_ASAP7_75t_L g312 ( .A(n_118), .B(n_276), .Y(n_312) );
OR2x2_ASAP7_75t_L g329 ( .A(n_118), .B(n_222), .Y(n_329) );
INVx1_ASAP7_75t_L g364 ( .A(n_118), .Y(n_364) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_118), .Y(n_386) );
OR2x2_ASAP7_75t_L g400 ( .A(n_118), .B(n_333), .Y(n_400) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_118), .B(n_222), .Y(n_404) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_144), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_129), .B(n_141), .Y(n_119) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g234 ( .A(n_122), .Y(n_234) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
AND2x6_ASAP7_75t_L g137 ( .A(n_123), .B(n_132), .Y(n_137) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g139 ( .A(n_125), .B(n_134), .Y(n_139) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
AND2x2_ASAP7_75t_L g133 ( .A(n_128), .B(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx3_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
AND2x4_ASAP7_75t_L g180 ( .A(n_133), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g176 ( .A(n_134), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_140), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_137), .B(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_140), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_140), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_140), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_140), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_140), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_140), .A2(n_441), .B(n_442), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_140), .A2(n_449), .B(n_450), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_140), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_140), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_140), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_140), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_140), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_SL g171 ( .A(n_141), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_141), .A2(n_507), .B(n_508), .Y(n_506) );
BUFx4f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_143), .B(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g195 ( .A(n_143), .B(n_146), .Y(n_195) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g356 ( .A(n_148), .B(n_312), .Y(n_356) );
AND2x2_ASAP7_75t_L g403 ( .A(n_148), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_157), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
AND2x2_ASAP7_75t_L g266 ( .A(n_150), .B(n_157), .Y(n_266) );
INVx2_ASAP7_75t_L g273 ( .A(n_150), .Y(n_273) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_150), .Y(n_394) );
BUFx3_ASAP7_75t_L g410 ( .A(n_150), .Y(n_410) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_151), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_151), .A2(n_438), .B(n_439), .Y(n_437) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_151), .A2(n_466), .B(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_157), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g333 ( .A(n_157), .B(n_273), .Y(n_333) );
INVx1_ASAP7_75t_L g351 ( .A(n_157), .Y(n_351) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_157), .Y(n_367) );
INVx1_ASAP7_75t_L g389 ( .A(n_157), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_157), .B(n_268), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_157), .B(n_222), .Y(n_426) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_166), .Y(n_158) );
INVx4_ASAP7_75t_L g231 ( .A(n_159), .Y(n_231) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_159), .A2(n_456), .B(n_462), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_165), .Y(n_160) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_186), .Y(n_168) );
AND2x4_ASAP7_75t_L g240 ( .A(n_169), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g251 ( .A(n_169), .Y(n_251) );
AND2x2_ASAP7_75t_L g256 ( .A(n_169), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g291 ( .A(n_169), .B(n_196), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_169), .B(n_197), .Y(n_301) );
OR2x2_ASAP7_75t_L g381 ( .A(n_169), .B(n_296), .Y(n_381) );
OAI322xp33_ASAP7_75t_L g411 ( .A1(n_169), .A2(n_324), .A3(n_363), .B1(n_396), .B2(n_412), .C1(n_413), .C2(n_414), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_169), .B(n_394), .Y(n_412) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
AOI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_185), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_179), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_174), .A2(n_180), .B1(n_224), .B2(n_226), .Y(n_223) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_178), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_186), .A2(n_358), .B1(n_362), .B2(n_365), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_186), .A2(n_418), .B(n_419), .C(n_422), .Y(n_417) );
AND2x4_ASAP7_75t_SL g186 ( .A(n_187), .B(n_196), .Y(n_186) );
AND2x4_ASAP7_75t_L g239 ( .A(n_187), .B(n_207), .Y(n_239) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
INVx5_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
INVx2_ASAP7_75t_L g264 ( .A(n_187), .Y(n_264) );
AND2x2_ASAP7_75t_L g287 ( .A(n_187), .B(n_197), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_187), .B(n_206), .Y(n_316) );
OR2x2_ASAP7_75t_L g325 ( .A(n_187), .B(n_245), .Y(n_325) );
OR2x2_ASAP7_75t_L g340 ( .A(n_187), .B(n_254), .Y(n_340) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_195), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_195), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_195), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_195), .B(n_230), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g232 ( .A(n_195), .B(n_233), .C(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_195), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_195), .A2(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_196), .B(n_216), .Y(n_215) );
INVx3_ASAP7_75t_SL g324 ( .A(n_196), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_196), .B(n_255), .Y(n_347) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
AND2x2_ASAP7_75t_L g244 ( .A(n_197), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g258 ( .A(n_197), .B(n_207), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_197), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_197), .B(n_207), .Y(n_296) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_197), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_197), .B(n_255), .Y(n_371) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_203), .Y(n_198) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_204), .A2(n_208), .B(n_214), .Y(n_207) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_204), .A2(n_208), .B(n_214), .Y(n_254) );
AOI21x1_ASAP7_75t_L g445 ( .A1(n_204), .A2(n_446), .B(n_452), .Y(n_445) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_207), .Y(n_277) );
AND2x2_ASAP7_75t_L g361 ( .A(n_207), .B(n_245), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_213), .Y(n_208) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_220), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_217), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x6_ASAP7_75t_SL g425 ( .A(n_218), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_219), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_219), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g373 ( .A(n_219), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_220), .A2(n_282), .B1(n_285), .B2(n_292), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_221), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g317 ( .A(n_221), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_221), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_221), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
AND2x2_ASAP7_75t_L g267 ( .A(n_222), .B(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g276 ( .A(n_222), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_222), .A2(n_283), .B1(n_335), .B2(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g342 ( .A(n_222), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_222), .B(n_336), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_222), .B(n_266), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_222), .B(n_273), .Y(n_415) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_228), .Y(n_222) );
INVx3_ASAP7_75t_L g517 ( .A(n_231), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_242), .B(n_246), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
NAND4xp25_ASAP7_75t_SL g285 ( .A(n_238), .B(n_286), .C(n_288), .D(n_290), .Y(n_285) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_239), .B(n_346), .Y(n_375) );
AND2x2_ASAP7_75t_L g402 ( .A(n_239), .B(n_240), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_239), .B(n_262), .Y(n_413) );
INVx1_ASAP7_75t_L g278 ( .A(n_240), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_240), .A2(n_303), .B1(n_314), .B2(n_317), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_240), .B(n_253), .C(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_240), .B(n_255), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_240), .B(n_263), .Y(n_406) );
AND2x2_ASAP7_75t_L g338 ( .A(n_241), .B(n_245), .Y(n_338) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_241), .Y(n_399) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
INVx1_ASAP7_75t_L g384 ( .A(n_244), .Y(n_384) );
AND2x2_ASAP7_75t_L g391 ( .A(n_244), .B(n_255), .Y(n_391) );
BUFx2_ASAP7_75t_L g346 ( .A(n_245), .Y(n_346) );
NAND3xp33_ASAP7_75t_SL g247 ( .A(n_248), .B(n_269), .C(n_281), .Y(n_247) );
OAI31xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_256), .A3(n_259), .B(n_265), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_249), .A2(n_303), .B1(n_307), .B2(n_308), .Y(n_302) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
OR2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_289), .Y(n_288) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_251), .B(n_315), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_252), .A2(n_354), .B(n_384), .C(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_253), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_254), .B(n_262), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_254), .B(n_287), .Y(n_307) );
AND2x2_ASAP7_75t_L g424 ( .A(n_257), .B(n_346), .Y(n_424) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g280 ( .A(n_258), .B(n_264), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_263), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g355 ( .A(n_263), .B(n_338), .Y(n_355) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_264), .B(n_338), .Y(n_344) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g336 ( .A(n_266), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_267), .B(n_367), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_277), .A3(n_278), .B1(n_279), .B2(n_758), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_270), .A2(n_355), .B1(n_391), .B2(n_392), .C(n_395), .Y(n_390) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g283 ( .A(n_275), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g388 ( .A(n_276), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_277), .B(n_299), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_279), .A2(n_322), .B1(n_326), .B2(n_330), .C(n_334), .Y(n_321) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_284), .A2(n_298), .B(n_302), .C(n_313), .Y(n_297) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_290), .A2(n_300), .A3(n_349), .B1(n_396), .B2(n_397), .C1(n_398), .C2(n_400), .Y(n_395) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_293), .A2(n_423), .B(n_425), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g379 ( .A1(n_299), .A2(n_380), .B(n_382), .C(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g421 ( .A(n_306), .B(n_387), .Y(n_421) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_312), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g396 ( .A(n_312), .Y(n_396) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g352 ( .A1(n_316), .A2(n_353), .A3(n_355), .B(n_356), .Y(n_352) );
NOR2x1_ASAP7_75t_L g319 ( .A(n_320), .B(n_378), .Y(n_319) );
NAND5xp2_ASAP7_75t_L g320 ( .A(n_321), .B(n_341), .C(n_352), .D(n_357), .E(n_368), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_324), .A2(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g392 ( .A(n_328), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_345), .C(n_348), .Y(n_341) );
INVxp33_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OR2x2_ASAP7_75t_L g370 ( .A(n_346), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_349), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_SL g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g420 ( .A(n_361), .Y(n_420) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_370), .A2(n_375), .B(n_376), .Y(n_374) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_390), .C(n_401), .D(n_417), .Y(n_378) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_388), .B(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_624), .Y(n_427) );
NOR4xp75_ASAP7_75t_L g428 ( .A(n_429), .B(n_547), .C(n_572), .D(n_599), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_484), .B(n_525), .Y(n_429) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_431), .B(n_468), .C(n_475), .D(n_479), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_453), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_435), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_435), .B(n_472), .Y(n_618) );
AND2x2_ASAP7_75t_L g643 ( .A(n_435), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g668 ( .A(n_435), .B(n_463), .Y(n_668) );
AND2x2_ASAP7_75t_L g709 ( .A(n_435), .B(n_477), .Y(n_709) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_436), .B(n_474), .Y(n_481) );
AND2x2_ASAP7_75t_L g483 ( .A(n_436), .B(n_455), .Y(n_483) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_436), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g544 ( .A(n_436), .Y(n_544) );
AND2x2_ASAP7_75t_L g550 ( .A(n_436), .B(n_477), .Y(n_550) );
BUFx2_ASAP7_75t_L g563 ( .A(n_436), .Y(n_563) );
AND2x4_ASAP7_75t_L g594 ( .A(n_436), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g641 ( .A(n_436), .B(n_642), .Y(n_641) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .Y(n_436) );
INVx1_ASAP7_75t_L g635 ( .A(n_444), .Y(n_635) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
AND2x2_ASAP7_75t_L g477 ( .A(n_445), .B(n_455), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_453), .B(n_653), .Y(n_706) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g543 ( .A(n_454), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_463), .Y(n_454) );
INVx2_ASAP7_75t_L g473 ( .A(n_455), .Y(n_473) );
INVx2_ASAP7_75t_L g534 ( .A(n_455), .Y(n_534) );
AND2x2_ASAP7_75t_L g644 ( .A(n_455), .B(n_474), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
INVx2_ASAP7_75t_L g532 ( .A(n_463), .Y(n_532) );
BUFx3_ASAP7_75t_L g549 ( .A(n_463), .Y(n_549) );
AND2x2_ASAP7_75t_L g576 ( .A(n_463), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AND2x4_ASAP7_75t_L g470 ( .A(n_464), .B(n_465), .Y(n_470) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx2_ASAP7_75t_L g478 ( .A(n_469), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_469), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g647 ( .A(n_469), .B(n_587), .Y(n_647) );
AND2x2_ASAP7_75t_L g671 ( .A(n_469), .B(n_481), .Y(n_671) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g567 ( .A(n_470), .B(n_473), .Y(n_567) );
AND2x2_ASAP7_75t_L g649 ( .A(n_470), .B(n_642), .Y(n_649) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g692 ( .A(n_472), .Y(n_692) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g577 ( .A(n_473), .Y(n_577) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_474), .Y(n_581) );
INVx2_ASAP7_75t_L g589 ( .A(n_474), .Y(n_589) );
INVx1_ASAP7_75t_L g595 ( .A(n_474), .Y(n_595) );
AOI222xp33_ASAP7_75t_SL g525 ( .A1(n_475), .A2(n_526), .B1(n_530), .B2(n_535), .C1(n_542), .C2(n_545), .Y(n_525) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g602 ( .A(n_477), .Y(n_602) );
BUFx2_ASAP7_75t_L g631 ( .A(n_477), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_478), .A2(n_626), .B(n_630), .C(n_638), .Y(n_625) );
OR2x2_ASAP7_75t_L g696 ( .A(n_478), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g704 ( .A(n_478), .B(n_609), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_SL g661 ( .A(n_481), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g679 ( .A(n_481), .B(n_567), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_481), .B(n_659), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_482), .B(n_549), .Y(n_687) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g609 ( .A(n_483), .B(n_581), .Y(n_609) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_504), .Y(n_485) );
INVx1_ASAP7_75t_L g703 ( .A(n_486), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
AND2x2_ASAP7_75t_L g546 ( .A(n_487), .B(n_505), .Y(n_546) );
INVx1_ASAP7_75t_L g623 ( .A(n_487), .Y(n_623) );
OR2x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_505), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_487), .B(n_554), .Y(n_688) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g529 ( .A(n_488), .Y(n_529) );
OR2x2_ASAP7_75t_L g561 ( .A(n_488), .B(n_515), .Y(n_561) );
AND2x2_ASAP7_75t_L g570 ( .A(n_488), .B(n_497), .Y(n_570) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_488), .B(n_505), .Y(n_598) );
AND2x2_ASAP7_75t_L g645 ( .A(n_488), .B(n_540), .Y(n_645) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g528 ( .A(n_497), .Y(n_528) );
INVx1_ASAP7_75t_L g538 ( .A(n_497), .Y(n_538) );
AND2x2_ASAP7_75t_L g554 ( .A(n_497), .B(n_541), .Y(n_554) );
INVx2_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
OR2x2_ASAP7_75t_L g655 ( .A(n_497), .B(n_505), .Y(n_655) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
NOR2x1_ASAP7_75t_SL g540 ( .A(n_505), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_515), .Y(n_571) );
BUFx2_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
INVx2_ASAP7_75t_SL g617 ( .A(n_505), .Y(n_617) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_513), .Y(n_505) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g527 ( .A(n_515), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g673 ( .A(n_515), .B(n_615), .Y(n_673) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_516) );
AO21x1_ASAP7_75t_SL g541 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_526), .A2(n_550), .B(n_690), .C(n_694), .Y(n_689) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_527), .B(n_605), .Y(n_640) );
BUFx2_ASAP7_75t_L g604 ( .A(n_528), .Y(n_604) );
OR2x2_ASAP7_75t_L g552 ( .A(n_529), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g637 ( .A(n_529), .B(n_571), .Y(n_637) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_614), .Y(n_658) );
INVx2_ASAP7_75t_L g665 ( .A(n_529), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_530), .A2(n_671), .B(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g612 ( .A(n_531), .B(n_594), .Y(n_612) );
OR2x2_ASAP7_75t_L g691 ( .A(n_531), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_532), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
AND2x2_ASAP7_75t_L g642 ( .A(n_534), .B(n_589), .Y(n_642) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g627 ( .A(n_537), .B(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_SL g636 ( .A(n_537), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_537), .B(n_546), .Y(n_669) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g545 ( .A(n_538), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g664 ( .A(n_539), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g614 ( .A(n_540), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g584 ( .A(n_541), .B(n_559), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g591 ( .A1(n_542), .A2(n_592), .A3(n_594), .B(n_596), .Y(n_591) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_544), .B(n_567), .Y(n_593) );
AO21x1_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
OR2x2_ASAP7_75t_L g603 ( .A(n_549), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g708 ( .A(n_549), .Y(n_708) );
INVx2_ASAP7_75t_SL g693 ( .A(n_550), .Y(n_693) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g597 ( .A(n_553), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g681 ( .A(n_553), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_554), .B(n_617), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_562), .B1(n_566), .B2(n_568), .Y(n_555) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_556), .A2(n_675), .B(n_676), .Y(n_674) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g629 ( .A(n_561), .B(n_590), .Y(n_629) );
OR2x2_ASAP7_75t_L g654 ( .A(n_561), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_563), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_563), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g653 ( .A(n_563), .Y(n_653) );
INVx2_ASAP7_75t_L g582 ( .A(n_564), .Y(n_582) );
INVx1_ASAP7_75t_L g662 ( .A(n_565), .Y(n_662) );
AND2x2_ASAP7_75t_L g585 ( .A(n_567), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g659 ( .A(n_567), .Y(n_659) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_573), .B(n_591), .Y(n_572) );
OAI321xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .A3(n_583), .B1(n_584), .B2(n_585), .C(n_590), .Y(n_573) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_574), .A2(n_605), .A3(n_700), .B1(n_702), .B2(n_704), .C1(n_705), .C2(n_710), .Y(n_699) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_579), .B(n_659), .Y(n_676) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g684 ( .A(n_582), .Y(n_684) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g616 ( .A(n_584), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI21xp33_ASAP7_75t_SL g683 ( .A1(n_587), .A2(n_593), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx3_ASAP7_75t_L g605 ( .A(n_598), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_619), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B1(n_606), .B2(n_607), .C(n_610), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_602), .Y(n_621) );
AND2x2_ASAP7_75t_L g606 ( .A(n_604), .B(n_605), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_613), .B1(n_616), .B2(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g622 ( .A(n_614), .B(n_623), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_617), .A2(n_706), .B(n_707), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_656), .C(n_677), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_629), .A2(n_664), .B1(n_691), .B2(n_693), .Y(n_690) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B(n_636), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_631), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_637), .A2(n_679), .B1(n_680), .B2(n_683), .C(n_685), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_643), .B2(n_645), .C(n_646), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g675 ( .A(n_641), .Y(n_675) );
INVx1_ASAP7_75t_L g697 ( .A(n_642), .Y(n_697) );
INVx1_ASAP7_75t_SL g695 ( .A(n_643), .Y(n_695) );
AOI31xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .A3(n_650), .B(n_654), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_647), .A2(n_657), .B1(n_659), .B2(n_660), .C(n_759), .Y(n_656) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B(n_666), .C(n_674), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g672 ( .A(n_665), .B(n_673), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_669), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g701 ( .A(n_673), .Y(n_701) );
BUFx2_ASAP7_75t_SL g710 ( .A(n_673), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_689), .C(n_699), .Y(n_677) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B(n_688), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .Y(n_694) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
CKINVDCx11_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_734), .Y(n_727) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_730), .B(n_733), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_SL g749 ( .A(n_731), .B(n_733), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_731), .A2(n_752), .B(n_755), .Y(n_751) );
INVx1_ASAP7_75t_SL g745 ( .A(n_734), .Y(n_745) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_R g738 ( .A(n_735), .Y(n_738) );
BUFx2_ASAP7_75t_L g756 ( .A(n_735), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B(n_744), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx9p33_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx11_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx8_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
endmodule