module real_aes_7850_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_0), .A2(n_205), .B(n_208), .C(n_303), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_1), .A2(n_240), .B(n_330), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_2), .A2(n_171), .B1(n_177), .B2(n_178), .Y(n_170) );
INVx1_ASAP7_75t_L g177 ( .A(n_2), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_3), .B(n_280), .Y(n_337) );
INVx1_ASAP7_75t_L g191 ( .A(n_4), .Y(n_191) );
AND2x6_ASAP7_75t_L g205 ( .A(n_4), .B(n_189), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_4), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g263 ( .A(n_5), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_6), .A2(n_80), .B1(n_81), .B2(n_169), .Y(n_79) );
INVx1_ASAP7_75t_L g169 ( .A(n_6), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_6), .B(n_216), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_7), .A2(n_33), .B1(n_129), .B2(n_134), .Y(n_128) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_29), .B1(n_90), .B2(n_91), .Y(n_89) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_9), .A2(n_69), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_9), .Y(n_174) );
INVx1_ASAP7_75t_L g224 ( .A(n_10), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_11), .A2(n_214), .B(n_288), .C(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_12), .B(n_280), .Y(n_291) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_13), .A2(n_31), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_14), .B(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_15), .A2(n_274), .B(n_275), .C(n_277), .Y(n_273) );
AOI22xp33_ASAP7_75t_SL g157 ( .A1(n_16), .A2(n_19), .B1(n_158), .B2(n_160), .Y(n_157) );
AOI22xp33_ASAP7_75t_SL g139 ( .A1(n_17), .A2(n_38), .B1(n_140), .B2(n_143), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_18), .B(n_216), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_20), .A2(n_73), .B1(n_102), .B2(n_109), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_21), .B(n_216), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_22), .Y(n_320) );
INVx1_ASAP7_75t_L g212 ( .A(n_23), .Y(n_212) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_24), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_25), .Y(n_301) );
AOI22xp33_ASAP7_75t_SL g146 ( .A1(n_26), .A2(n_53), .B1(n_147), .B2(n_152), .Y(n_146) );
INVx1_ASAP7_75t_L g246 ( .A(n_27), .Y(n_246) );
INVx2_ASAP7_75t_L g203 ( .A(n_28), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_30), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g182 ( .A1(n_31), .A2(n_43), .B1(n_51), .B2(n_183), .C(n_184), .Y(n_182) );
INVxp67_ASAP7_75t_L g185 ( .A(n_31), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_32), .A2(n_274), .B(n_333), .C(n_335), .Y(n_332) );
INVxp67_ASAP7_75t_L g247 ( .A(n_34), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_35), .A2(n_208), .B(n_211), .C(n_219), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g331 ( .A(n_36), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_37), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_39), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_40), .Y(n_242) );
INVx1_ASAP7_75t_L g272 ( .A(n_41), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_42), .A2(n_172), .B1(n_173), .B2(n_176), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_42), .Y(n_172) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_43), .A2(n_64), .B1(n_90), .B2(n_94), .Y(n_97) );
INVxp67_ASAP7_75t_L g186 ( .A(n_43), .Y(n_186) );
CKINVDCx14_ASAP7_75t_R g259 ( .A(n_44), .Y(n_259) );
INVx1_ASAP7_75t_L g189 ( .A(n_45), .Y(n_189) );
INVx1_ASAP7_75t_L g223 ( .A(n_46), .Y(n_223) );
INVx1_ASAP7_75t_SL g334 ( .A(n_47), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_48), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_49), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g323 ( .A(n_50), .Y(n_323) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_68), .B1(n_90), .B2(n_91), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_52), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_54), .A2(n_240), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g526 ( .A(n_54), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_55), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_56), .A2(n_240), .B(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g163 ( .A1(n_57), .A2(n_75), .B1(n_164), .B2(n_167), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_58), .A2(n_239), .B(n_241), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_59), .Y(n_206) );
INVx1_ASAP7_75t_L g286 ( .A(n_60), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_61), .A2(n_80), .B1(n_81), .B2(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_61), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_62), .A2(n_240), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g289 ( .A(n_63), .Y(n_289) );
INVx2_ASAP7_75t_L g221 ( .A(n_65), .Y(n_221) );
INVx1_ASAP7_75t_L g304 ( .A(n_66), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_67), .A2(n_208), .B(n_322), .C(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g175 ( .A(n_69), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_70), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_71), .B(n_228), .Y(n_266) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
INVx2_ASAP7_75t_L g276 ( .A(n_74), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_76), .B(n_123), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_179), .B1(n_192), .B2(n_510), .C(n_513), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_170), .Y(n_78) );
AOI22xp5_ASAP7_75t_SL g514 ( .A1(n_80), .A2(n_81), .B1(n_263), .B2(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_138), .C(n_156), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_114), .Y(n_83) );
OAI21xp5_ASAP7_75t_SL g84 ( .A1(n_85), .A2(n_100), .B(n_101), .Y(n_84) );
INVx2_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x6_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x4_ASAP7_75t_L g135 ( .A(n_88), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_93), .Y(n_88) );
AND2x2_ASAP7_75t_L g108 ( .A(n_89), .B(n_97), .Y(n_108) );
INVx2_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx2_ASAP7_75t_L g107 ( .A(n_93), .Y(n_107) );
AND2x2_ASAP7_75t_L g119 ( .A(n_93), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g127 ( .A(n_93), .B(n_120), .Y(n_127) );
INVx1_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
AND2x2_ASAP7_75t_L g141 ( .A(n_95), .B(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g166 ( .A(n_95), .B(n_126), .Y(n_166) );
AND2x4_ASAP7_75t_L g168 ( .A(n_95), .B(n_119), .Y(n_168) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g121 ( .A(n_96), .B(n_99), .Y(n_121) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g151 ( .A(n_97), .B(n_137), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_97), .B(n_99), .Y(n_155) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g106 ( .A(n_99), .Y(n_106) );
INVx1_ASAP7_75t_L g137 ( .A(n_99), .Y(n_137) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g113 ( .A(n_106), .Y(n_113) );
AND2x2_ASAP7_75t_L g142 ( .A(n_107), .B(n_120), .Y(n_142) );
AND2x4_ASAP7_75t_L g112 ( .A(n_108), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g131 ( .A(n_108), .B(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx12f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_122), .C(n_128), .Y(n_114) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
AND2x2_ASAP7_75t_L g150 ( .A(n_119), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g125 ( .A(n_121), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g145 ( .A(n_121), .B(n_142), .Y(n_145) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x6_ASAP7_75t_L g154 ( .A(n_133), .B(n_155), .Y(n_154) );
BUFx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_146), .Y(n_138) );
BUFx2_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g159 ( .A(n_142), .B(n_151), .Y(n_159) );
AND2x4_ASAP7_75t_L g161 ( .A(n_142), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx6_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_163), .Y(n_156) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx11_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_171), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_173), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
AND3x1_ASAP7_75t_SL g181 ( .A(n_182), .B(n_187), .C(n_190), .Y(n_181) );
INVxp67_ASAP7_75t_L g519 ( .A(n_182), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx1_ASAP7_75t_SL g521 ( .A(n_187), .Y(n_521) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_187), .A2(n_201), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g532 ( .A(n_187), .Y(n_532) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_188), .B(n_191), .Y(n_525) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_SL g531 ( .A(n_190), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR5x1_ASAP7_75t_L g193 ( .A(n_194), .B(n_404), .C(n_468), .D(n_484), .E(n_499), .Y(n_193) );
NAND4xp25_ASAP7_75t_L g194 ( .A(n_195), .B(n_338), .C(n_365), .D(n_388), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_281), .B(n_292), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_230), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_SL g315 ( .A(n_198), .Y(n_315) );
AND2x4_ASAP7_75t_L g351 ( .A(n_198), .B(n_340), .Y(n_351) );
OR2x2_ASAP7_75t_L g361 ( .A(n_198), .B(n_317), .Y(n_361) );
OR2x2_ASAP7_75t_L g407 ( .A(n_198), .B(n_233), .Y(n_407) );
AND2x2_ASAP7_75t_L g421 ( .A(n_198), .B(n_316), .Y(n_421) );
AND2x2_ASAP7_75t_L g464 ( .A(n_198), .B(n_354), .Y(n_464) );
AND2x2_ASAP7_75t_L g471 ( .A(n_198), .B(n_328), .Y(n_471) );
AND2x2_ASAP7_75t_L g490 ( .A(n_198), .B(n_380), .Y(n_490) );
AND2x2_ASAP7_75t_L g508 ( .A(n_198), .B(n_350), .Y(n_508) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_225), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_206), .B(n_207), .C(n_220), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_200), .A2(n_301), .B(n_302), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_200), .A2(n_320), .B(n_321), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_201), .B(n_205), .Y(n_200) );
AND2x4_ASAP7_75t_L g240 ( .A(n_201), .B(n_205), .Y(n_240) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx1_ASAP7_75t_L g218 ( .A(n_202), .Y(n_218) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g209 ( .A(n_203), .Y(n_209) );
INVx1_ASAP7_75t_L g278 ( .A(n_203), .Y(n_278) );
INVx1_ASAP7_75t_L g210 ( .A(n_204), .Y(n_210) );
INVx3_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_204), .Y(n_216) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
BUFx3_ASAP7_75t_L g219 ( .A(n_205), .Y(n_219) );
INVx4_ASAP7_75t_SL g250 ( .A(n_205), .Y(n_250) );
INVx5_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
AND2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
BUFx3_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_209), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_215), .C(n_217), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g245 ( .A1(n_213), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_245) );
INVx5_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_214), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g261 ( .A(n_216), .Y(n_261) );
INVx4_ASAP7_75t_L g274 ( .A(n_216), .Y(n_274) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_218), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g254 ( .A(n_220), .Y(n_254) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_220), .A2(n_257), .B(n_266), .Y(n_256) );
INVx1_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g229 ( .A(n_221), .B(n_222), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx3_ASAP7_75t_L g280 ( .A(n_227), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_227), .B(n_310), .Y(n_309) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_227), .A2(n_319), .B(n_326), .Y(n_318) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g236 ( .A(n_229), .Y(n_236) );
INVx1_ASAP7_75t_L g473 ( .A(n_230), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_255), .Y(n_230) );
AND2x2_ASAP7_75t_L g383 ( .A(n_231), .B(n_316), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_231), .B(n_403), .Y(n_402) );
AOI32xp33_ASAP7_75t_L g416 ( .A1(n_231), .A2(n_417), .A3(n_420), .B1(n_422), .B2(n_426), .Y(n_416) );
AND2x2_ASAP7_75t_L g486 ( .A(n_231), .B(n_380), .Y(n_486) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g350 ( .A(n_233), .B(n_317), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_233), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g392 ( .A(n_233), .B(n_339), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_233), .B(n_471), .Y(n_470) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_237), .B(n_251), .Y(n_233) );
INVx1_ASAP7_75t_L g355 ( .A(n_234), .Y(n_355) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_238), .A2(n_252), .B(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_239), .Y(n_512) );
BUFx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_243), .B(n_244), .C(n_250), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_243), .A2(n_250), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_243), .A2(n_250), .B(n_272), .C(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_243), .A2(n_250), .B(n_286), .C(n_287), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_243), .A2(n_250), .B(n_331), .C(n_332), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_248), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_248), .B(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g306 ( .A(n_249), .Y(n_306) );
INVx1_ASAP7_75t_L g325 ( .A(n_250), .Y(n_325) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_254), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g357 ( .A(n_255), .B(n_296), .Y(n_357) );
AND2x2_ASAP7_75t_L g433 ( .A(n_255), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g505 ( .A(n_255), .Y(n_505) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_267), .Y(n_255) );
OR2x2_ASAP7_75t_L g295 ( .A(n_256), .B(n_268), .Y(n_295) );
AND2x2_ASAP7_75t_L g312 ( .A(n_256), .B(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_256), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g364 ( .A(n_256), .Y(n_364) );
AND2x2_ASAP7_75t_L g391 ( .A(n_256), .B(n_268), .Y(n_391) );
BUFx3_ASAP7_75t_L g394 ( .A(n_256), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_256), .B(n_369), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_256), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g515 ( .A(n_263), .Y(n_515) );
INVx2_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
INVx2_ASAP7_75t_L g345 ( .A(n_267), .Y(n_345) );
AND2x2_ASAP7_75t_L g363 ( .A(n_267), .B(n_343), .Y(n_363) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g374 ( .A(n_268), .B(n_283), .Y(n_374) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_268), .Y(n_387) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_279), .Y(n_268) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_269), .A2(n_284), .B(n_291), .Y(n_283) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_269), .A2(n_329), .B(n_337), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_274), .B(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_282), .B(n_394), .Y(n_444) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g313 ( .A(n_283), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_283), .B(n_363), .C(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g370 ( .A(n_283), .B(n_343), .Y(n_370) );
AND2x2_ASAP7_75t_L g390 ( .A(n_283), .B(n_343), .Y(n_390) );
AND2x2_ASAP7_75t_L g434 ( .A(n_283), .B(n_298), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_311), .B(n_314), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x2_ASAP7_75t_L g509 ( .A(n_294), .B(n_434), .Y(n_509) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_295), .A2(n_407), .B1(n_449), .B2(n_451), .Y(n_448) );
OR2x2_ASAP7_75t_L g455 ( .A(n_295), .B(n_370), .Y(n_455) );
OR2x2_ASAP7_75t_L g479 ( .A(n_295), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_295), .B(n_399), .Y(n_492) );
AND2x2_ASAP7_75t_L g385 ( .A(n_296), .B(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_296), .A2(n_458), .B(n_473), .Y(n_472) );
AOI32xp33_ASAP7_75t_L g493 ( .A1(n_296), .A2(n_383), .A3(n_494), .B1(n_496), .B2(n_497), .Y(n_493) );
OR2x2_ASAP7_75t_L g504 ( .A(n_296), .B(n_505), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g372 ( .A(n_297), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_297), .B(n_386), .Y(n_451) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
AND2x2_ASAP7_75t_L g409 ( .A(n_298), .B(n_374), .Y(n_409) );
AND3x2_ASAP7_75t_L g418 ( .A(n_298), .B(n_312), .C(n_419), .Y(n_418) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_309), .Y(n_298) );
O2A1O1Ixp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_307), .C(n_308), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_305), .A2(n_308), .B(n_323), .C(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_313), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_313), .B(n_343), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g339 ( .A(n_315), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g379 ( .A(n_315), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g397 ( .A(n_315), .B(n_328), .Y(n_397) );
AND2x2_ASAP7_75t_L g415 ( .A(n_315), .B(n_317), .Y(n_415) );
OR2x2_ASAP7_75t_L g429 ( .A(n_315), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g475 ( .A(n_315), .B(n_403), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_316), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_328), .Y(n_316) );
AND2x2_ASAP7_75t_L g376 ( .A(n_317), .B(n_354), .Y(n_376) );
OR2x2_ASAP7_75t_L g430 ( .A(n_317), .B(n_354), .Y(n_430) );
AND2x2_ASAP7_75t_L g483 ( .A(n_317), .B(n_340), .Y(n_483) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g381 ( .A(n_318), .Y(n_381) );
AND2x2_ASAP7_75t_L g403 ( .A(n_318), .B(n_328), .Y(n_403) );
INVx2_ASAP7_75t_L g340 ( .A(n_328), .Y(n_340) );
INVx1_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_346), .C(n_358), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_339), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g502 ( .A(n_339), .Y(n_502) );
AND2x2_ASAP7_75t_L g380 ( .A(n_340), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_343), .B(n_344), .Y(n_352) );
INVx1_ASAP7_75t_L g437 ( .A(n_343), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_343), .B(n_364), .Y(n_461) );
AND2x2_ASAP7_75t_L g477 ( .A(n_343), .B(n_391), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_344), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_352), .B1(n_353), .B2(n_356), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_349), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_350), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g375 ( .A(n_351), .B(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_SL g440 ( .A1(n_351), .A2(n_393), .B1(n_441), .B2(n_446), .C(n_448), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_351), .B(n_414), .Y(n_447) );
INVx1_ASAP7_75t_L g507 ( .A(n_353), .Y(n_507) );
BUFx3_ASAP7_75t_L g414 ( .A(n_354), .Y(n_414) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI21xp33_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g423 ( .A(n_360), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_360), .B(n_414), .Y(n_467) );
INVx1_ASAP7_75t_L g424 ( .A(n_361), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_361), .B(n_414), .Y(n_425) );
INVxp67_ASAP7_75t_L g445 ( .A(n_363), .Y(n_445) );
AND2x2_ASAP7_75t_L g386 ( .A(n_364), .B(n_387), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .B(n_375), .C(n_377), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g400 ( .A(n_368), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_369), .B(n_400), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_369), .B(n_391), .Y(n_442) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_372), .A2(n_378), .B1(n_382), .B2(n_384), .Y(n_377) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g393 ( .A(n_374), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_439), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_376), .A2(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_380), .A2(n_389), .B1(n_392), .B2(n_393), .C(n_395), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_380), .B(n_414), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_380), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g496 ( .A(n_386), .Y(n_496) );
INVxp67_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_389), .Y(n_426) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g465 ( .A(n_390), .B(n_394), .Y(n_465) );
INVx1_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_394), .B(n_409), .Y(n_469) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .A3(n_400), .B1(n_401), .B2(n_402), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g408 ( .A(n_403), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_403), .B(n_435), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_403), .B(n_464), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_403), .B(n_414), .Y(n_503) );
NAND5xp2_ASAP7_75t_L g404 ( .A(n_405), .B(n_427), .C(n_440), .D(n_452), .E(n_453), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_410), .B2(n_412), .C(n_416), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_411), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_414), .B(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_415), .A2(n_428), .B1(n_431), .B2(n_435), .Y(n_427) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
OAI211xp5_ASAP7_75t_SL g422 ( .A1(n_418), .A2(n_423), .B(n_424), .C(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g450 ( .A(n_430), .Y(n_450) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_439), .B(n_488), .Y(n_498) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B1(n_458), .B2(n_462), .C1(n_465), .C2(n_466), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_472), .B2(n_474), .C(n_476), .Y(n_468) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g488 ( .A(n_480), .Y(n_488) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_487), .B1(n_489), .B2(n_491), .C(n_493), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B(n_504), .C(n_506), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
OAI322xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_516), .A3(n_520), .B1(n_522), .B2(n_526), .C1(n_527), .C2(n_529), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
endmodule