module fake_netlist_5_2219_n_1846 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1846);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1846;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1668;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_124),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_56),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_50),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_116),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_103),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_19),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_21),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_101),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_33),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_11),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_36),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_127),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_102),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_20),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_55),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_78),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_69),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_13),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_34),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_54),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_168),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_37),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_167),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_88),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_27),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_8),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_64),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_38),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_44),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_67),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_115),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_68),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_24),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_35),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_37),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_157),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_77),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_54),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_94),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_20),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_171),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_33),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_105),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_178),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_164),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_119),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_153),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_147),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_143),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_90),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_64),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_70),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_177),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_170),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_149),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_123),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_60),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_162),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_28),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_63),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_155),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_49),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_152),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_99),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_158),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_53),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_18),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_23),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_29),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_75),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_42),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_145),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_32),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_132),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_2),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_30),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_79),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_130),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_11),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_109),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_135),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_85),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_71),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_154),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_95),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_12),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_82),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_48),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_41),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_96),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_159),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_15),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_179),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_60),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_83),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_24),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_111),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_30),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_110),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_41),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_22),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_97),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_175),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_9),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_50),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_9),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_129),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_131),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_59),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_52),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_144),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_106),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_17),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_48),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_26),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_8),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_197),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_331),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_198),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_214),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_189),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_233),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_228),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_303),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_234),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_223),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_271),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_234),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_280),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_234),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_234),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_348),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_235),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_236),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_196),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_226),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_243),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_261),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_246),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_250),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_227),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_260),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_188),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_229),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_231),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_232),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_267),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_268),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_195),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_237),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_238),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_193),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_200),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_273),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_242),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_189),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_190),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_241),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_277),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_296),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_296),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_282),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_286),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_247),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_248),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_205),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_217),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_230),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_196),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_255),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_254),
.B(n_245),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_288),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_294),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_254),
.B(n_0),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_196),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_297),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_251),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_259),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_300),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_253),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_263),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_265),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_208),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_264),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_345),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_269),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_305),
.B(n_3),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_354),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_377),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_399),
.B(n_245),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_388),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_362),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_393),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_362),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_184),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_249),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_400),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_401),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_402),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_408),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_369),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_411),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_420),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_427),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_428),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_364),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_433),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_419),
.B(n_363),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_386),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_366),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_365),
.B(n_354),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_441),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_371),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_374),
.B(n_184),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_367),
.B(n_266),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_447),
.B(n_206),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_444),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_407),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_448),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_394),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_R g500 ( 
.A(n_450),
.B(n_270),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_384),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_367),
.B(n_292),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_249),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_384),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_385),
.B(n_272),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_418),
.B(n_186),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_410),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_412),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_385),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_389),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_389),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_370),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_391),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_434),
.B(n_252),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_368),
.B(n_252),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_372),
.B(n_274),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_481),
.A2(n_392),
.B1(n_403),
.B2(n_397),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_456),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_375),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_512),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_466),
.B(n_437),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_461),
.Y(n_538)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_459),
.A2(n_451),
.B(n_283),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_466),
.B(n_392),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_512),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_483),
.B(n_502),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_456),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_501),
.Y(n_547)
);

INVx4_ASAP7_75t_SL g548 ( 
.A(n_456),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_466),
.B(n_503),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_483),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_466),
.B(n_397),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_513),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_524),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_403),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_405),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_500),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_513),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_505),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_471),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_505),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_499),
.B(n_405),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_506),
.B(n_376),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_274),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_465),
.B(n_387),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_465),
.B(n_323),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_509),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_517),
.A2(n_390),
.B1(n_279),
.B2(n_317),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_488),
.B(n_323),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_488),
.B(n_416),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_510),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_514),
.B(n_416),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_460),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_413),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_504),
.B(n_195),
.Y(n_587)
);

CKINVDCx14_ASAP7_75t_R g588 ( 
.A(n_461),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_499),
.B(n_421),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_499),
.B(n_425),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_471),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_454),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_525),
.B(n_195),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_464),
.B(n_438),
.C(n_432),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

INVxp33_ASAP7_75t_SL g598 ( 
.A(n_515),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_471),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_471),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_464),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_519),
.B(n_425),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_485),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_485),
.B(n_195),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_516),
.B(n_378),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

INVx6_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_491),
.B(n_195),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_527),
.B(n_426),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_479),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_455),
.B(n_215),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_528),
.A2(n_360),
.B1(n_298),
.B2(n_326),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_455),
.B(n_426),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_494),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_520),
.B(n_435),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_528),
.A2(n_307),
.B1(n_355),
.B2(n_321),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_457),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_495),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_457),
.B(n_435),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_528),
.A2(n_313),
.B1(n_443),
.B2(n_446),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_458),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_495),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_495),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_458),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_463),
.B(n_244),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_462),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_472),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_463),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_520),
.B(n_436),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_496),
.B(n_436),
.Y(n_635)
);

BUFx4f_ASAP7_75t_L g636 ( 
.A(n_522),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_484),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_522),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_496),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_496),
.B(n_439),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_523),
.B(n_430),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_508),
.B(n_439),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_508),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_476),
.B(n_442),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_373),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_528),
.B(n_442),
.Y(n_646)
);

INVx4_ASAP7_75t_SL g647 ( 
.A(n_476),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_489),
.B(n_275),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_526),
.A2(n_191),
.B1(n_211),
.B2(n_311),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_531),
.B(n_431),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_526),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_492),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_529),
.B(n_440),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_492),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

INVxp33_ASAP7_75t_L g657 ( 
.A(n_530),
.Y(n_657)
);

INVx8_ASAP7_75t_L g658 ( 
.A(n_467),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_531),
.B(n_445),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_473),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_531),
.B(n_256),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_473),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_531),
.B(n_186),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_482),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_482),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_482),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_468),
.B(n_379),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_521),
.B(n_276),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_521),
.B(n_257),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_469),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_470),
.B(n_187),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_497),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_474),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_475),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_477),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_487),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_478),
.A2(n_320),
.B1(n_316),
.B2(n_221),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_480),
.A2(n_332),
.B1(n_222),
.B2(n_221),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_486),
.B(n_258),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_493),
.B(n_281),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_597),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_597),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_643),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_549),
.B(n_278),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_553),
.B(n_291),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_554),
.A2(n_383),
.B1(n_325),
.B2(n_318),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_578),
.A2(n_310),
.B1(n_285),
.B2(n_287),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_553),
.B(n_293),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_646),
.B(n_312),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_607),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_534),
.B(n_187),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_578),
.B(n_334),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_603),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_537),
.B(n_335),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_663),
.B(n_338),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_603),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_557),
.B(n_208),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_572),
.A2(n_352),
.B1(n_208),
.B2(n_212),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_663),
.B(n_289),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_619),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_634),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_631),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_424),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_589),
.B(n_290),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_586),
.B(n_449),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_532),
.B(n_295),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_589),
.B(n_299),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_301),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_583),
.B(n_192),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_555),
.A2(n_551),
.B1(n_541),
.B2(n_566),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_592),
.B(n_621),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_583),
.B(n_571),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_SL g716 ( 
.A(n_638),
.B(n_185),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_631),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_654),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_654),
.Y(n_719)
);

NOR3xp33_ASAP7_75t_L g720 ( 
.A(n_677),
.B(n_190),
.C(n_361),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_590),
.B(n_192),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_592),
.B(n_302),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_616),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_621),
.B(n_315),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_557),
.A2(n_324),
.B1(n_328),
.B2(n_322),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_660),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_656),
.B(n_319),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_612),
.A2(n_327),
.B1(n_194),
.B2(n_203),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_641),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_584),
.B(n_194),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_586),
.B(n_449),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_671),
.B(n_329),
.C(n_361),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_671),
.B(n_612),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_660),
.Y(n_734)
);

OAI221xp5_ASAP7_75t_L g735 ( 
.A1(n_620),
.A2(n_336),
.B1(n_359),
.B2(n_358),
.C(n_222),
.Y(n_735)
);

CKINVDCx11_ASAP7_75t_R g736 ( 
.A(n_672),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_SL g737 ( 
.A1(n_598),
.A2(n_306),
.B1(n_339),
.B2(n_240),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_636),
.B(n_208),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_641),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_585),
.B(n_203),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_593),
.B(n_204),
.Y(n_741)
);

AND2x6_ASAP7_75t_SL g742 ( 
.A(n_670),
.B(n_452),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_204),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_625),
.B(n_207),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_636),
.B(n_208),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_642),
.A2(n_344),
.B1(n_207),
.B2(n_340),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_628),
.B(n_632),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_651),
.B(n_208),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_572),
.A2(n_208),
.B1(n_189),
.B2(n_212),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_616),
.B(n_213),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_651),
.B(n_208),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_623),
.B(n_213),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_586),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_662),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_657),
.B(n_216),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_657),
.B(n_535),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_641),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_543),
.B(n_216),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_218),
.B1(n_219),
.B2(n_357),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_545),
.B(n_218),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_SL g762 ( 
.A(n_562),
.B(n_219),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_547),
.B(n_220),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_658),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_563),
.B(n_220),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_565),
.B(n_224),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_680),
.B(n_224),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_567),
.B(n_573),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_640),
.B(n_340),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_574),
.B(n_344),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_643),
.B(n_347),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_601),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_SL g773 ( 
.A(n_556),
.B(n_239),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_579),
.B(n_347),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_622),
.A2(n_353),
.B(n_356),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_668),
.B(n_353),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_556),
.B(n_356),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_648),
.A2(n_357),
.B(n_358),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_617),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_633),
.B(n_284),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_652),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_662),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_650),
.B(n_284),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_602),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_576),
.A2(n_359),
.B(n_351),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_679),
.B(n_199),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_655),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_536),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_536),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_538),
.B(n_333),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_679),
.B(n_575),
.C(n_596),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_588),
.B(n_333),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_540),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_540),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_658),
.B(n_314),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_542),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_570),
.B(n_199),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_613),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_644),
.B(n_201),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_645),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_542),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_594),
.B(n_72),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_650),
.B(n_314),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_552),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_552),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_570),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_658),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_659),
.B(n_314),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_570),
.B(n_201),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_617),
.B(n_626),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_570),
.B(n_342),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_608),
.B(n_81),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_539),
.A2(n_342),
.B(n_350),
.C(n_346),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_570),
.B(n_342),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_558),
.B(n_561),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_598),
.B(n_202),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_645),
.B(n_647),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_560),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_560),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_614),
.B(n_202),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_580),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_617),
.B(n_209),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_614),
.A2(n_336),
.B1(n_350),
.B2(n_346),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_645),
.A2(n_351),
.B1(n_343),
.B2(n_341),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_550),
.B(n_343),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_580),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_558),
.B(n_337),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_594),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_558),
.B(n_210),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_664),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_561),
.B(n_329),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_645),
.A2(n_581),
.B1(n_629),
.B2(n_614),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_626),
.B(n_330),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_626),
.B(n_333),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_626),
.B(n_181),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_678),
.B(n_3),
.C(n_4),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_639),
.B(n_174),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_588),
.B(n_172),
.Y(n_839)
);

BUFx6f_ASAP7_75t_SL g840 ( 
.A(n_672),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_564),
.B(n_161),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_564),
.B(n_156),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_674),
.B(n_5),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_564),
.B(n_142),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_764),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_698),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_715),
.B(n_577),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_806),
.A2(n_587),
.B(n_661),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_733),
.A2(n_606),
.B1(n_568),
.B2(n_673),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_708),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_714),
.A2(n_661),
.B(n_669),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_SL g853 ( 
.A(n_840),
.B(n_582),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_702),
.B(n_544),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_577),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_699),
.A2(n_669),
.B(n_600),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_577),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_691),
.A2(n_666),
.B(n_599),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_699),
.A2(n_600),
.B(n_610),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_810),
.A2(n_815),
.B(n_696),
.Y(n_860)
);

AOI22x1_ASAP7_75t_L g861 ( 
.A1(n_683),
.A2(n_618),
.B1(n_627),
.B2(n_605),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_788),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_702),
.B(n_673),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_694),
.A2(n_649),
.B(n_610),
.C(n_615),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_817),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_723),
.B(n_637),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_786),
.A2(n_675),
.B(n_624),
.C(n_627),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_708),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_810),
.A2(n_533),
.B(n_546),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_697),
.A2(n_828),
.B(n_686),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_711),
.A2(n_533),
.B(n_546),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_723),
.B(n_676),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_767),
.B(n_599),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_703),
.B(n_582),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_757),
.A2(n_690),
.B(n_687),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_768),
.A2(n_599),
.B(n_627),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_790),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_708),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_771),
.A2(n_618),
.B(n_605),
.C(n_613),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_683),
.A2(n_614),
.B(n_629),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_695),
.B(n_639),
.Y(n_882)
);

AO21x1_ASAP7_75t_L g883 ( 
.A1(n_701),
.A2(n_629),
.B(n_604),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_753),
.A2(n_609),
.B1(n_630),
.B2(n_639),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_721),
.B(n_639),
.Y(n_885)
);

BUFx8_ASAP7_75t_SL g886 ( 
.A(n_840),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_693),
.B(n_629),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_784),
.B(n_630),
.Y(n_888)
);

CKINVDCx11_ASAP7_75t_R g889 ( 
.A(n_736),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_752),
.B(n_665),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_716),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_705),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_683),
.A2(n_604),
.B(n_611),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_747),
.A2(n_533),
.B(n_546),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_791),
.B(n_672),
.C(n_658),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_736),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_738),
.A2(n_533),
.B(n_546),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_685),
.Y(n_898)
);

BUFx12f_ASAP7_75t_L g899 ( 
.A(n_742),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_769),
.B(n_665),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_705),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_816),
.B(n_609),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_777),
.B(n_750),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_772),
.B(n_569),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_789),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_722),
.A2(n_569),
.B(n_559),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_731),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_R g908 ( 
.A(n_716),
.B(n_112),
.Y(n_908)
);

OAI321xp33_ASAP7_75t_L g909 ( 
.A1(n_688),
.A2(n_5),
.A3(n_6),
.B1(n_10),
.B2(n_12),
.C(n_14),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_731),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_685),
.A2(n_548),
.B(n_569),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_822),
.A2(n_604),
.B(n_14),
.C(n_15),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_738),
.A2(n_665),
.B(n_591),
.Y(n_913)
);

AND2x2_ASAP7_75t_SL g914 ( 
.A(n_773),
.B(n_665),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_754),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_781),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_798),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_745),
.A2(n_591),
.B(n_559),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_844),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_793),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_745),
.A2(n_591),
.B(n_559),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_840),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_799),
.B(n_611),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_707),
.B(n_10),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_836),
.B(n_16),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_748),
.A2(n_139),
.B(n_136),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_732),
.B(n_16),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_710),
.B(n_17),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_SL g929 ( 
.A(n_764),
.B(n_125),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_787),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_794),
.A2(n_118),
.B(n_117),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_751),
.A2(n_108),
.B(n_107),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_706),
.B(n_18),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_783),
.B(n_19),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_751),
.A2(n_831),
.B(n_829),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_807),
.B(n_23),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_803),
.B(n_25),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_825),
.B(n_29),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_827),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_792),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_756),
.B(n_32),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_804),
.A2(n_104),
.B(n_98),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_729),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_804),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_739),
.A2(n_93),
.B1(n_86),
.B2(n_44),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_808),
.B(n_43),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_724),
.A2(n_43),
.B(n_45),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_776),
.A2(n_45),
.B(n_46),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_818),
.A2(n_46),
.B(n_47),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_812),
.B(n_51),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_819),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_821),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_821),
.A2(n_53),
.B(n_58),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_796),
.A2(n_58),
.B(n_59),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_801),
.A2(n_61),
.B(n_62),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_807),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_817),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_754),
.A2(n_62),
.B(n_63),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_681),
.A2(n_65),
.B(n_66),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_758),
.B(n_66),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_682),
.A2(n_684),
.B(n_734),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_832),
.A2(n_797),
.B1(n_809),
.B2(n_800),
.Y(n_962)
);

AOI21xp33_ASAP7_75t_L g963 ( 
.A1(n_759),
.A2(n_774),
.B(n_761),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_779),
.A2(n_727),
.B(n_811),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_728),
.B(n_746),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_800),
.A2(n_814),
.B1(n_689),
.B2(n_802),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_805),
.A2(n_826),
.B(n_843),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_684),
.B(n_692),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_834),
.B(n_770),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_692),
.B(n_755),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_704),
.A2(n_782),
.B(n_755),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_704),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_834),
.B(n_765),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_717),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_779),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_SL g976 ( 
.A1(n_737),
.A2(n_839),
.B1(n_785),
.B2(n_735),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_837),
.B(n_709),
.C(n_780),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_718),
.A2(n_726),
.B(n_719),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_839),
.B(n_743),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_830),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_779),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_813),
.A2(n_822),
.B(n_833),
.C(n_778),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_730),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_740),
.B(n_744),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_795),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_741),
.B(n_766),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_841),
.A2(n_845),
.B(n_842),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_835),
.A2(n_838),
.B(n_763),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_835),
.A2(n_838),
.B(n_797),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_802),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_809),
.A2(n_820),
.B1(n_833),
.B2(n_725),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_795),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_760),
.B(n_780),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_824),
.B(n_823),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_720),
.B(n_749),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_775),
.B(n_700),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_795),
.B(n_762),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_817),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_817),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_772),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_777),
.B(n_675),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_694),
.A2(n_715),
.B(n_733),
.C(n_691),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_810),
.A2(n_699),
.B(n_714),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_733),
.B(n_702),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_715),
.B(n_723),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_694),
.A2(n_715),
.B(n_733),
.C(n_691),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_806),
.A2(n_557),
.B(n_714),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_699),
.A2(n_806),
.B(n_697),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_817),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_698),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_698),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_715),
.B(n_713),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_840),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_865),
.B(n_870),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_903),
.A2(n_965),
.B(n_1006),
.C(n_1002),
.Y(n_1015)
);

AO31x2_ASAP7_75t_L g1016 ( 
.A1(n_883),
.A2(n_982),
.A3(n_1007),
.B(n_989),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_1001),
.B(n_895),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_1012),
.A2(n_962),
.B1(n_991),
.B2(n_1005),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_865),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_1007),
.A2(n_900),
.B(n_890),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_865),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_914),
.B(n_927),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_1000),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_983),
.B(n_892),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_870),
.B(n_957),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_901),
.B(n_984),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_870),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_885),
.A2(n_964),
.B(n_876),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_981),
.B(n_898),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_878),
.B(n_866),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_967),
.A2(n_978),
.B(n_971),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_986),
.B(n_876),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_873),
.B(n_888),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_940),
.B(n_919),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_916),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_849),
.A2(n_935),
.B(n_871),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_891),
.B(n_850),
.Y(n_1037)
);

AOI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_994),
.A2(n_993),
.B(n_973),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_969),
.B(n_848),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_846),
.B(n_956),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_936),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_963),
.B(n_939),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_849),
.A2(n_852),
.B(n_881),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_852),
.A2(n_987),
.B(n_887),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_941),
.A2(n_864),
.B(n_924),
.C(n_928),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_977),
.A2(n_902),
.B1(n_976),
.B2(n_979),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_857),
.A2(n_874),
.B(n_859),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1004),
.B(n_898),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_875),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_934),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_935),
.A2(n_855),
.B(n_996),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_937),
.B(n_946),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_961),
.B(n_860),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_880),
.A2(n_995),
.B(n_867),
.C(n_938),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_925),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_957),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_854),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_851),
.B(n_868),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_905),
.B(n_920),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_877),
.B(n_869),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_877),
.A2(n_894),
.B(n_906),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_957),
.Y(n_1062)
);

BUFx4f_ASAP7_75t_L g1063 ( 
.A(n_998),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_960),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_913),
.A2(n_859),
.B(n_856),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_951),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_960),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_990),
.A2(n_966),
.B1(n_907),
.B2(n_879),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_910),
.B(n_933),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_950),
.A2(n_923),
.B(n_988),
.C(n_893),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_L g1071 ( 
.A(n_846),
.B(n_956),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_998),
.B(n_999),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_863),
.B(n_847),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_999),
.B(n_1009),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_968),
.A2(n_970),
.B(n_972),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_949),
.A2(n_953),
.A3(n_943),
.B(n_954),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_952),
.B(n_974),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1009),
.B(n_853),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1011),
.A2(n_884),
.B(n_904),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_882),
.A2(n_918),
.B(n_921),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1008),
.B(n_980),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_936),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1008),
.B(n_975),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_992),
.B(n_908),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_L g1086 ( 
.A(n_992),
.B(n_922),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_975),
.B(n_915),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_981),
.B(n_948),
.Y(n_1088)
);

NOR2x1_ASAP7_75t_L g1089 ( 
.A(n_997),
.B(n_936),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_926),
.A2(n_932),
.B(n_929),
.Y(n_1090)
);

AO21x1_ASAP7_75t_L g1091 ( 
.A1(n_912),
.A2(n_947),
.B(n_948),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_949),
.A2(n_953),
.B(n_954),
.Y(n_1092)
);

AND3x4_ASAP7_75t_L g1093 ( 
.A(n_899),
.B(n_889),
.C(n_886),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_947),
.B(n_955),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_958),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_992),
.B(n_1013),
.Y(n_1096)
);

AO21x1_ASAP7_75t_L g1097 ( 
.A1(n_945),
.A2(n_909),
.B(n_985),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1013),
.A2(n_911),
.B(n_872),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_896),
.A2(n_883),
.A3(n_982),
.B(n_1007),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_865),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_849),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_865),
.B(n_870),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1000),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1012),
.B(n_903),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_L g1108 ( 
.A(n_1012),
.B(n_865),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_883),
.A2(n_982),
.A3(n_1007),
.B(n_989),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1000),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1012),
.A2(n_715),
.B1(n_903),
.B2(n_965),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_1012),
.B(n_865),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1005),
.B(n_723),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_L g1115 ( 
.A(n_1001),
.B(n_764),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_886),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1012),
.B(n_903),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1012),
.B(n_903),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_849),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_911),
.A2(n_872),
.B(n_861),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_917),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1007),
.A2(n_557),
.B(n_989),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_917),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_849),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1012),
.B(n_903),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1007),
.A2(n_557),
.B(n_989),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_849),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_862),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1012),
.B(n_903),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1012),
.B(n_903),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_914),
.B(n_850),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_895),
.B(n_675),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_895),
.B(n_675),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_858),
.A2(n_1007),
.B(n_989),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_903),
.Y(n_1136)
);

AOI21xp33_ASAP7_75t_L g1137 ( 
.A1(n_903),
.A2(n_715),
.B(n_712),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_865),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1007),
.A2(n_557),
.B(n_885),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1007),
.A2(n_557),
.B(n_989),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1005),
.B(n_637),
.Y(n_1143)
);

AND2x2_ASAP7_75t_SL g1144 ( 
.A(n_914),
.B(n_927),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1012),
.B(n_903),
.Y(n_1145)
);

INVx11_ASAP7_75t_L g1146 ( 
.A(n_1013),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_911),
.A2(n_872),
.B(n_861),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_959),
.A2(n_942),
.B(n_931),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_L g1149 ( 
.A(n_1001),
.B(n_764),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1012),
.B(n_903),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_903),
.A2(n_694),
.B(n_712),
.C(n_733),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1000),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1012),
.B(n_903),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1012),
.B(n_903),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1137),
.A2(n_1151),
.B(n_1112),
.C(n_1015),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1035),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1096),
.B(n_1121),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1116),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1034),
.B(n_1022),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1056),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1101),
.A2(n_1124),
.B(n_1127),
.C(n_1119),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1032),
.A2(n_1028),
.B(n_1044),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1023),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1118),
.B(n_1125),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1144),
.B(n_1143),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1014),
.B(n_1072),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_L g1172 ( 
.A(n_1118),
.B(n_1125),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1123),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1110),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1032),
.A2(n_1043),
.B(n_1051),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1131),
.B(n_1136),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1104),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1122),
.A2(n_1142),
.B(n_1126),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1063),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_SL g1182 ( 
.A1(n_1038),
.A2(n_1094),
.B(n_1132),
.C(n_1036),
.Y(n_1182)
);

NOR2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1136),
.B(n_1145),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1145),
.B(n_1150),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1056),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1150),
.B(n_1153),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1027),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1018),
.A2(n_1097),
.B1(n_1046),
.B2(n_1154),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1063),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1128),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1153),
.B(n_1154),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1041),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1039),
.B(n_1052),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1045),
.A2(n_1091),
.B(n_1090),
.C(n_1054),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1026),
.B(n_1069),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1146),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_1047),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1026),
.B(n_1057),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1042),
.B(n_1152),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1039),
.B(n_1052),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1083),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1027),
.Y(n_1202)
);

AO21x1_ASAP7_75t_L g1203 ( 
.A1(n_1090),
.A2(n_1068),
.B(n_1094),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1024),
.B(n_1049),
.Y(n_1204)
);

CKINVDCx6p67_ASAP7_75t_R g1205 ( 
.A(n_1027),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1089),
.A2(n_1042),
.B1(n_1058),
.B2(n_1073),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1014),
.B(n_1072),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1024),
.B(n_1050),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1209)
);

CKINVDCx6p67_ASAP7_75t_R g1210 ( 
.A(n_1062),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1048),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1108),
.A2(n_1113),
.B1(n_1079),
.B2(n_1085),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1050),
.B(n_1078),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1103),
.A2(n_1111),
.B(n_1106),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1062),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_1025),
.B(n_1074),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1102),
.B(n_1078),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1102),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1062),
.B(n_1140),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1133),
.A2(n_1134),
.B1(n_1017),
.B2(n_1086),
.Y(n_1220)
);

OR2x2_ASAP7_75t_SL g1221 ( 
.A(n_1140),
.B(n_1048),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1100),
.B(n_1019),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1053),
.A2(n_1020),
.B(n_1092),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1080),
.B(n_1021),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1105),
.A2(n_1139),
.B(n_1138),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1077),
.B(n_1066),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1129),
.A2(n_1141),
.B(n_1020),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1082),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1115),
.B(n_1149),
.Y(n_1230)
);

INVx3_ASAP7_75t_R g1231 ( 
.A(n_1093),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1025),
.B(n_1099),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1099),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1040),
.B(n_1071),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1099),
.B(n_1076),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1098),
.Y(n_1236)
);

NAND2x1_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_1066),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1095),
.A2(n_1088),
.B1(n_1029),
.B2(n_1082),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1087),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1060),
.A2(n_1065),
.B(n_1031),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1076),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1084),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1070),
.B(n_1075),
.C(n_1059),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1076),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_1084),
.Y(n_1245)
);

NOR2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1081),
.B(n_1016),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1016),
.B(n_1109),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1135),
.A2(n_1109),
.B(n_1061),
.C(n_1120),
.Y(n_1248)
);

OAI21xp33_ASAP7_75t_L g1249 ( 
.A1(n_1147),
.A2(n_715),
.B(n_1137),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1143),
.B(n_637),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1143),
.B(n_637),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1035),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1121),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1143),
.B(n_637),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1137),
.A2(n_903),
.B(n_733),
.C(n_1151),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1056),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1121),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1104),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1112),
.A2(n_1107),
.B1(n_1118),
.B2(n_1117),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1137),
.A2(n_903),
.B(n_733),
.C(n_1151),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1104),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1056),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1116),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1112),
.B(n_929),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1137),
.A2(n_715),
.B(n_534),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1056),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1093),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1282)
);

INVx3_ASAP7_75t_SL g1283 ( 
.A(n_1116),
.Y(n_1283)
);

BUFx4_ASAP7_75t_SL g1284 ( 
.A(n_1116),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1023),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1137),
.A2(n_903),
.B(n_733),
.C(n_1151),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1032),
.A2(n_1044),
.B(n_1028),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1096),
.B(n_658),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1096),
.B(n_658),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1027),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1056),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1023),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1178),
.B(n_1193),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1171),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1261),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1292),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1193),
.B(n_1200),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1261),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1253),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1156),
.B(n_1266),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1188),
.A2(n_1276),
.B1(n_1258),
.B2(n_1191),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1265),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1242),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1200),
.B(n_1166),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1265),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1176),
.B(n_1236),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1221),
.Y(n_1309)
);

BUFx8_ASAP7_75t_SL g1310 ( 
.A(n_1281),
.Y(n_1310)
);

BUFx4f_ASAP7_75t_SL g1311 ( 
.A(n_1215),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1166),
.B(n_1168),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1170),
.A2(n_1161),
.B1(n_1263),
.B2(n_1158),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1241),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1174),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1237),
.B(n_1212),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1245),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1263),
.A2(n_1278),
.B1(n_1267),
.B2(n_1269),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1160),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1163),
.B(n_1211),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1169),
.A2(n_1267),
.B1(n_1258),
.B2(n_1262),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1235),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1247),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1183),
.A2(n_1244),
.B1(n_1172),
.B2(n_1271),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1169),
.B(n_1173),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1171),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1233),
.A2(n_1225),
.B1(n_1199),
.B2(n_1257),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1173),
.A2(n_1278),
.B1(n_1257),
.B2(n_1262),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1238),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1232),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1184),
.A2(n_1252),
.B1(n_1269),
.B2(n_1191),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1239),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1184),
.B(n_1186),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1186),
.B(n_1252),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1254),
.Y(n_1336)
);

INVx5_ASAP7_75t_L g1337 ( 
.A(n_1187),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1270),
.B(n_1276),
.Y(n_1338)
);

BUFx2_ASAP7_75t_R g1339 ( 
.A(n_1196),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1284),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1202),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1282),
.A2(n_1206),
.B1(n_1177),
.B2(n_1213),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1207),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1282),
.A2(n_1209),
.B1(n_1195),
.B2(n_1204),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1250),
.A2(n_1255),
.B1(n_1251),
.B2(n_1201),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1208),
.A2(n_1264),
.B1(n_1256),
.B2(n_1287),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1227),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1203),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1211),
.B(n_1155),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1220),
.A2(n_1198),
.B1(n_1217),
.B2(n_1159),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1190),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1217),
.B(n_1207),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1283),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1223),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1249),
.A2(n_1260),
.B1(n_1275),
.B2(n_1192),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1214),
.A2(n_1226),
.B(n_1228),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1246),
.Y(n_1357)
);

CKINVDCx6p67_ASAP7_75t_R g1358 ( 
.A(n_1273),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1216),
.B(n_1182),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1194),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1167),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1288),
.B(n_1164),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1292),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1175),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1219),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_SL g1366 ( 
.A(n_1210),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1243),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1248),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1224),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1224),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1289),
.A2(n_1290),
.B1(n_1230),
.B2(n_1272),
.Y(n_1371)
);

AOI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1240),
.A2(n_1216),
.B(n_1222),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1240),
.Y(n_1373)
);

NOR2x1_ASAP7_75t_R g1374 ( 
.A(n_1181),
.B(n_1189),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1202),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1216),
.B(n_1222),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1162),
.B(n_1185),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1285),
.A2(n_1294),
.B1(n_1290),
.B2(n_1205),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1185),
.A2(n_1234),
.B(n_1209),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1259),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1234),
.Y(n_1381)
);

BUFx2_ASAP7_75t_R g1382 ( 
.A(n_1231),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1218),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1259),
.B(n_1280),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_SL g1385 ( 
.A(n_1268),
.B(n_1280),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1234),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1268),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1165),
.A2(n_1272),
.B1(n_1274),
.B2(n_1291),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1165),
.A2(n_1274),
.B1(n_1286),
.B2(n_1291),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1281),
.A2(n_1137),
.B1(n_965),
.B2(n_1112),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1293),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1292),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1277),
.A2(n_1137),
.B1(n_773),
.B2(n_1112),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1180),
.A2(n_1197),
.B(n_1148),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1277),
.A2(n_1144),
.B1(n_1022),
.B2(n_773),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1229),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1277),
.A2(n_1137),
.B1(n_773),
.B2(n_1112),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1229),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1157),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1279),
.B(n_1112),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1178),
.B(n_1193),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1157),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1157),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1261),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1277),
.A2(n_1137),
.B1(n_965),
.B2(n_1112),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1273),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_R g1408 ( 
.A(n_1196),
.B(n_736),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1277),
.A2(n_1137),
.B1(n_965),
.B2(n_1112),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1215),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1284),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_SL g1414 ( 
.A(n_1353),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1367),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1362),
.A2(n_1356),
.B(n_1368),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1373),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1367),
.Y(n_1418)
);

AO21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1330),
.A2(n_1348),
.B(n_1368),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1369),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1305),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1308),
.Y(n_1423)
);

CKINVDCx10_ASAP7_75t_R g1424 ( 
.A(n_1382),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1370),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1427)
);

AO21x1_ASAP7_75t_L g1428 ( 
.A1(n_1401),
.A2(n_1398),
.B(n_1394),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1349),
.B(n_1314),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1357),
.B(n_1308),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1349),
.B(n_1314),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1333),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1372),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1295),
.B(n_1402),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1346),
.A2(n_1395),
.B(n_1359),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1308),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1360),
.A2(n_1359),
.B(n_1330),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1302),
.B(n_1311),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1303),
.A2(n_1316),
.B(n_1322),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1295),
.B(n_1402),
.Y(n_1441)
);

BUFx4f_ASAP7_75t_L g1442 ( 
.A(n_1316),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1333),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1406),
.A2(n_1409),
.B(n_1391),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1312),
.B(n_1334),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1308),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1447)
);

INVx8_ASAP7_75t_L g1448 ( 
.A(n_1352),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1357),
.B(n_1381),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1399),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1381),
.B(n_1386),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1379),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1301),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1317),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1335),
.B(n_1338),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1335),
.B(n_1338),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1347),
.B(n_1354),
.Y(n_1457)
);

AOI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1378),
.A2(n_1385),
.B(n_1326),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1347),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1319),
.B(n_1404),
.Y(n_1460)
);

BUFx4f_ASAP7_75t_SL g1461 ( 
.A(n_1353),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1300),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1304),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1400),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1329),
.B(n_1332),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1403),
.Y(n_1466)
);

OR2x2_ASAP7_75t_SL g1467 ( 
.A(n_1307),
.B(n_1405),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1309),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1351),
.A2(n_1350),
.B(n_1371),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1336),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1328),
.A2(n_1325),
.B(n_1342),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1315),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1341),
.A2(n_1355),
.B(n_1380),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1380),
.A2(n_1389),
.B(n_1388),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1313),
.B(n_1297),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1315),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1344),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1376),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1376),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1435),
.B(n_1384),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1444),
.A2(n_1396),
.B1(n_1345),
.B2(n_1410),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1435),
.B(n_1412),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1444),
.A2(n_1475),
.B1(n_1465),
.B2(n_1477),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1435),
.B(n_1376),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1435),
.B(n_1412),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1412),
.B(n_1377),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1416),
.B(n_1390),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1478),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1415),
.B(n_1318),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1413),
.B(n_1417),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1413),
.B(n_1377),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1416),
.B(n_1410),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1416),
.B(n_1383),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1467),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1415),
.B(n_1361),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1413),
.B(n_1420),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1420),
.B(n_1296),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1428),
.A2(n_1296),
.B1(n_1343),
.B2(n_1327),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1436),
.B(n_1296),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1425),
.B(n_1296),
.Y(n_1501)
);

BUFx4f_ASAP7_75t_SL g1502 ( 
.A(n_1472),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1465),
.A2(n_1358),
.B1(n_1383),
.B2(n_1327),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1418),
.B(n_1365),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1418),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1467),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1421),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1430),
.Y(n_1508)
);

NAND2x1_ASAP7_75t_L g1509 ( 
.A(n_1440),
.B(n_1375),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1440),
.A2(n_1352),
.B(n_1393),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1459),
.B(n_1445),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1436),
.B(n_1327),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1453),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1438),
.B(n_1343),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1438),
.B(n_1343),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1438),
.B(n_1343),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1475),
.A2(n_1358),
.B1(n_1393),
.B2(n_1366),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1416),
.B(n_1392),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1436),
.B(n_1375),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1428),
.A2(n_1364),
.B1(n_1310),
.B2(n_1320),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1438),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1416),
.B(n_1392),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1433),
.B(n_1392),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_1496),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1490),
.B(n_1462),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1482),
.A2(n_1477),
.B1(n_1442),
.B2(n_1471),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1496),
.B(n_1462),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1484),
.A2(n_1521),
.B(n_1482),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1433),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1471),
.C(n_1454),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1487),
.B(n_1443),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1517),
.A2(n_1432),
.B1(n_1443),
.B2(n_1470),
.C(n_1460),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1503),
.A2(n_1471),
.B1(n_1469),
.B2(n_1430),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1510),
.A2(n_1439),
.B1(n_1471),
.B2(n_1432),
.C(n_1468),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1460),
.C(n_1468),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1454),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1503),
.B(n_1426),
.C(n_1427),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1414),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1510),
.A2(n_1430),
.B(n_1458),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1502),
.A2(n_1442),
.B1(n_1471),
.B2(n_1476),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1493),
.B(n_1427),
.C(n_1426),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1445),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_R g1548 ( 
.A(n_1502),
.B(n_1340),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1495),
.B(n_1442),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1495),
.A2(n_1430),
.B(n_1458),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1506),
.A2(n_1485),
.B(n_1493),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1552)
);

OAI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1493),
.A2(n_1422),
.B(n_1437),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1492),
.B(n_1456),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1483),
.B(n_1456),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1506),
.B(n_1442),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1486),
.B(n_1434),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1494),
.B(n_1474),
.C(n_1450),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1513),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1494),
.B(n_1474),
.C(n_1450),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1494),
.B(n_1488),
.C(n_1504),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1488),
.B(n_1474),
.C(n_1480),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1509),
.A2(n_1476),
.B1(n_1472),
.B2(n_1480),
.C(n_1479),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1485),
.A2(n_1434),
.B1(n_1437),
.B2(n_1422),
.C(n_1455),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1486),
.B(n_1436),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1486),
.B(n_1446),
.Y(n_1566)
);

NAND4xp25_ASAP7_75t_L g1567 ( 
.A(n_1488),
.B(n_1447),
.C(n_1457),
.D(n_1464),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1485),
.B(n_1446),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1509),
.A2(n_1461),
.B1(n_1479),
.B2(n_1455),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1491),
.B(n_1429),
.Y(n_1571)
);

NOR3xp33_ASAP7_75t_L g1572 ( 
.A(n_1489),
.B(n_1473),
.C(n_1452),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1491),
.B(n_1429),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1524),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1491),
.B(n_1431),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_L g1576 ( 
.A(n_1489),
.B(n_1473),
.C(n_1452),
.Y(n_1576)
);

NOR3xp33_ASAP7_75t_L g1577 ( 
.A(n_1489),
.B(n_1473),
.C(n_1452),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1522),
.B(n_1474),
.C(n_1466),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1561),
.B(n_1497),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1407),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1525),
.B(n_1498),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1559),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1532),
.B(n_1501),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1559),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1574),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1508),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1534),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1530),
.B(n_1519),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1535),
.A2(n_1469),
.B1(n_1423),
.B2(n_1446),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1508),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1568),
.B(n_1520),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1534),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1555),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1564),
.B(n_1501),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1565),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1541),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1555),
.B(n_1497),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1529),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1548),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1536),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1531),
.B(n_1514),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1547),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1533),
.B(n_1557),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1533),
.B(n_1497),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1557),
.Y(n_1609)
);

AND2x4_ASAP7_75t_SL g1610 ( 
.A(n_1572),
.B(n_1519),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1554),
.B(n_1514),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1571),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1575),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1546),
.B(n_1518),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1590),
.B(n_1535),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1576),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1618),
.B(n_1558),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1584),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1594),
.B(n_1556),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1614),
.A2(n_1527),
.B1(n_1539),
.B2(n_1538),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1594),
.B(n_1577),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1553),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1586),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1553),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1607),
.B(n_1556),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1601),
.B(n_1580),
.Y(n_1632)
);

AOI322xp5_ASAP7_75t_L g1633 ( 
.A1(n_1591),
.A2(n_1537),
.A3(n_1522),
.B1(n_1514),
.B2(n_1516),
.C1(n_1515),
.C2(n_1507),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1607),
.B(n_1515),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1618),
.B(n_1560),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1596),
.A2(n_1540),
.B1(n_1542),
.B2(n_1545),
.Y(n_1636)
);

AND2x2_ASAP7_75t_SL g1637 ( 
.A(n_1610),
.B(n_1423),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1550),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1595),
.A2(n_1544),
.B(n_1578),
.C(n_1562),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1612),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1515),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1595),
.B(n_1516),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1579),
.B(n_1578),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1579),
.B(n_1524),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1604),
.B(n_1516),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1586),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1589),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1589),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1609),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1524),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1593),
.B(n_1523),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1602),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1609),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1593),
.B(n_1523),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1518),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1505),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1617),
.B(n_1505),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1599),
.Y(n_1659)
);

XNOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1340),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1628),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1620),
.B(n_1603),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1633),
.A2(n_1563),
.B(n_1569),
.C(n_1612),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1593),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1646),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1646),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1657),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1657),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1658),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1650),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1587),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1638),
.B(n_1613),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1639),
.B(n_1613),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1658),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1639),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1613),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1650),
.Y(n_1682)
);

NOR2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1411),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1630),
.B(n_1605),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1619),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1637),
.B(n_1592),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1631),
.B(n_1602),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1640),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1622),
.B(n_1606),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1654),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1635),
.B(n_1600),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1592),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1647),
.Y(n_1698)
);

O2A1O1Ixp5_ASAP7_75t_L g1699 ( 
.A1(n_1635),
.A2(n_1583),
.B(n_1582),
.C(n_1585),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1649),
.B(n_1588),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1633),
.B(n_1643),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1647),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1692),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1689),
.B(n_1621),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1689),
.B(n_1621),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1666),
.B(n_1621),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1680),
.B(n_1659),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1701),
.A2(n_1625),
.B1(n_1624),
.B2(n_1659),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1666),
.B(n_1626),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1674),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1678),
.A2(n_1625),
.B1(n_1665),
.B2(n_1660),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1664),
.B(n_1642),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1686),
.B(n_1644),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1664),
.B(n_1624),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1660),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1678),
.Y(n_1717)
);

AOI21xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1671),
.A2(n_1411),
.B(n_1632),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1674),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1673),
.B(n_1408),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1692),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1675),
.A2(n_1469),
.B1(n_1626),
.B2(n_1449),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1662),
.B(n_1700),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1662),
.B(n_1626),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1700),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1661),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1684),
.B(n_1320),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1685),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1676),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1683),
.B(n_1619),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1677),
.A2(n_1423),
.B1(n_1642),
.B2(n_1446),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1681),
.B(n_1634),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1663),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1667),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1696),
.B(n_1644),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1668),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1685),
.A2(n_1697),
.B1(n_1672),
.B2(n_1679),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1711),
.Y(n_1739)
);

OAI322xp33_ASAP7_75t_L g1740 ( 
.A1(n_1712),
.A2(n_1696),
.A3(n_1694),
.B1(n_1670),
.B2(n_1669),
.C1(n_1698),
.C2(n_1695),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1685),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1711),
.Y(n_1743)
);

OAI21xp33_ASAP7_75t_SL g1744 ( 
.A1(n_1717),
.A2(n_1687),
.B(n_1682),
.Y(n_1744)
);

AOI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1709),
.A2(n_1716),
.B(n_1731),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1716),
.A2(n_1665),
.B(n_1699),
.C(n_1688),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1730),
.B(n_1690),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1720),
.Y(n_1748)
);

AOI222xp33_ASAP7_75t_L g1749 ( 
.A1(n_1715),
.A2(n_1708),
.B1(n_1731),
.B2(n_1726),
.C1(n_1713),
.C2(n_1721),
.Y(n_1749)
);

CKINVDCx14_ASAP7_75t_R g1750 ( 
.A(n_1728),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1718),
.A2(n_1697),
.B(n_1693),
.C(n_1691),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1724),
.B(n_1697),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1704),
.A2(n_1423),
.B1(n_1448),
.B2(n_1702),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1720),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1729),
.A2(n_1469),
.B1(n_1449),
.B2(n_1451),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1704),
.A2(n_1423),
.B1(n_1500),
.B2(n_1512),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1729),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1707),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1703),
.B(n_1688),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1703),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1718),
.B(n_1651),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1719),
.Y(n_1762)
);

OAI33xp33_ASAP7_75t_L g1763 ( 
.A1(n_1727),
.A2(n_1648),
.A3(n_1623),
.B1(n_1653),
.B2(n_1619),
.B3(n_1656),
.Y(n_1763)
);

CKINVDCx6p67_ASAP7_75t_R g1764 ( 
.A(n_1705),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1707),
.B(n_1652),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1757),
.B(n_1706),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1764),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1764),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1758),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1739),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1738),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1739),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1742),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1749),
.B(n_1710),
.Y(n_1774)
);

XOR2x2_ASAP7_75t_L g1775 ( 
.A(n_1761),
.B(n_1424),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1745),
.B(n_1710),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1742),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_SL g1780 ( 
.A(n_1751),
.B(n_1339),
.Y(n_1780)
);

AND2x4_ASAP7_75t_SL g1781 ( 
.A(n_1741),
.B(n_1320),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1765),
.B(n_1706),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1743),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1765),
.B(n_1727),
.Y(n_1785)
);

NAND2xp33_ASAP7_75t_L g1786 ( 
.A(n_1747),
.B(n_1719),
.Y(n_1786)
);

NOR2x1_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1722),
.Y(n_1787)
);

NOR3xp33_ASAP7_75t_L g1788 ( 
.A(n_1768),
.B(n_1750),
.C(n_1740),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1783),
.A2(n_1744),
.B(n_1754),
.C(n_1743),
.Y(n_1789)
);

NOR2xp67_ASAP7_75t_L g1790 ( 
.A(n_1766),
.B(n_1744),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1783),
.A2(n_1763),
.B1(n_1748),
.B2(n_1754),
.C(n_1723),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1780),
.A2(n_1753),
.B1(n_1723),
.B2(n_1755),
.C(n_1756),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1773),
.B(n_1748),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1774),
.A2(n_1755),
.B1(n_1732),
.B2(n_1734),
.C(n_1737),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1776),
.A2(n_1733),
.B1(n_1714),
.B2(n_1736),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1785),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1786),
.A2(n_1762),
.B1(n_1760),
.B2(n_1722),
.C(n_1737),
.Y(n_1797)
);

AOI31xp33_ASAP7_75t_L g1798 ( 
.A1(n_1767),
.A2(n_1424),
.A3(n_1760),
.B(n_1762),
.Y(n_1798)
);

NAND3x1_ASAP7_75t_L g1799 ( 
.A(n_1787),
.B(n_1735),
.C(n_1734),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1767),
.B(n_1714),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1799),
.A2(n_1790),
.B(n_1788),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1800),
.A2(n_1769),
.B1(n_1777),
.B2(n_1771),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1793),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_1789),
.B(n_1786),
.C(n_1777),
.Y(n_1804)
);

NOR3x1_ASAP7_75t_L g1805 ( 
.A(n_1794),
.B(n_1779),
.C(n_1782),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1796),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1795),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_SL g1808 ( 
.A(n_1798),
.B(n_1778),
.Y(n_1808)
);

NOR3x1_ASAP7_75t_L g1809 ( 
.A(n_1792),
.B(n_1784),
.C(n_1772),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_L g1810 ( 
.A(n_1791),
.B(n_1778),
.C(n_1770),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1797),
.B(n_1775),
.Y(n_1811)
);

AO22x2_ASAP7_75t_L g1812 ( 
.A1(n_1804),
.A2(n_1722),
.B1(n_1759),
.B2(n_1735),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_SL g1813 ( 
.A(n_1801),
.B(n_1775),
.C(n_1736),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1759),
.C(n_1781),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1811),
.A2(n_1781),
.B1(n_1759),
.B2(n_1423),
.Y(n_1815)
);

AND4x1_ASAP7_75t_L g1816 ( 
.A(n_1809),
.B(n_1805),
.C(n_1810),
.D(n_1803),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_L g1817 ( 
.A(n_1802),
.B(n_1374),
.C(n_1310),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1807),
.A2(n_1653),
.B(n_1648),
.C(n_1656),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1812),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1813),
.A2(n_1806),
.B1(n_1808),
.B2(n_1364),
.Y(n_1820)
);

AO22x1_ASAP7_75t_L g1821 ( 
.A1(n_1817),
.A2(n_1298),
.B1(n_1363),
.B2(n_1653),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1814),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1818),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1816),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1815),
.Y(n_1825)
);

AOI322xp5_ASAP7_75t_L g1826 ( 
.A1(n_1824),
.A2(n_1641),
.A3(n_1645),
.B1(n_1634),
.B2(n_1655),
.C1(n_1652),
.C2(n_1597),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1820),
.B(n_1655),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1820),
.B(n_1641),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1822),
.B(n_1623),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1823),
.B(n_1363),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_L g1831 ( 
.A(n_1819),
.B(n_1298),
.Y(n_1831)
);

XNOR2xp5_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1825),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1828),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1831),
.B(n_1821),
.Y(n_1834)
);

XNOR2xp5_ASAP7_75t_L g1835 ( 
.A(n_1832),
.B(n_1833),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1835),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1836),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1836),
.Y(n_1838)
);

OAI21xp33_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1832),
.B(n_1829),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1834),
.B(n_1827),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1840),
.B(n_1826),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1839),
.B(n_1651),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1841),
.A2(n_1298),
.B(n_1363),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1843),
.B(n_1842),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_R g1845 ( 
.A1(n_1844),
.A2(n_1448),
.B1(n_1363),
.B2(n_1387),
.C(n_1419),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1363),
.B(n_1375),
.C(n_1387),
.Y(n_1846)
);


endmodule