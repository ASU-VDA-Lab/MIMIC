module real_aes_4301_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_L g98 ( .A1(n_0), .A2(n_37), .B1(n_99), .B2(n_122), .Y(n_98) );
INVx1_ASAP7_75t_L g392 ( .A(n_1), .Y(n_392) );
INVx2_ASAP7_75t_SL g86 ( .A(n_2), .Y(n_86) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_3), .B(n_249), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_4), .A2(n_5), .B1(n_189), .B2(n_191), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_6), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_7), .A2(n_31), .B1(n_291), .B2(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_8), .A2(n_33), .B1(n_309), .B2(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_9), .A2(n_53), .B1(n_354), .B2(n_369), .Y(n_376) );
INVx1_ASAP7_75t_L g387 ( .A(n_10), .Y(n_387) );
INVx1_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_11), .B(n_60), .Y(n_172) );
INVxp67_ASAP7_75t_L g187 ( .A(n_11), .Y(n_187) );
INVx1_ASAP7_75t_L g390 ( .A(n_12), .Y(n_390) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_13), .A2(n_57), .B(n_242), .Y(n_241) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_13), .A2(n_57), .B(n_242), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_14), .B(n_104), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_15), .A2(n_55), .B1(n_354), .B2(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_16), .Y(n_81) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_17), .A2(n_44), .B1(n_143), .B2(n_146), .Y(n_142) );
INVx1_ASAP7_75t_L g384 ( .A(n_18), .Y(n_384) );
INVx1_ASAP7_75t_L g165 ( .A(n_19), .Y(n_165) );
BUFx3_ASAP7_75t_L g201 ( .A(n_20), .Y(n_201) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
AO22x1_ASAP7_75t_L g270 ( .A1(n_22), .A2(n_65), .B1(n_271), .B2(n_275), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_23), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_24), .B(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_24), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_25), .B(n_275), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g160 ( .A1(n_26), .A2(n_43), .B1(n_161), .B2(n_163), .C(n_164), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_27), .A2(n_75), .B1(n_177), .B2(n_179), .Y(n_176) );
AOI22x1_ASAP7_75t_L g353 ( .A1(n_28), .A2(n_74), .B1(n_333), .B2(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g105 ( .A(n_29), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_29), .B(n_59), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_30), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_32), .B(n_246), .Y(n_318) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_34), .A2(n_46), .B1(n_150), .B2(n_155), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_35), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_36), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g242 ( .A(n_38), .Y(n_242) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_39), .Y(n_212) );
AND2x4_ASAP7_75t_L g226 ( .A(n_39), .B(n_210), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_40), .A2(n_64), .B1(n_133), .B2(n_138), .Y(n_132) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_41), .Y(n_224) );
INVx2_ASAP7_75t_L g371 ( .A(n_42), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_45), .A2(n_61), .B1(n_291), .B2(n_333), .Y(n_332) );
CKINVDCx14_ASAP7_75t_R g282 ( .A(n_47), .Y(n_282) );
AND2x2_ASAP7_75t_L g316 ( .A(n_48), .B(n_275), .Y(n_316) );
OA22x2_ASAP7_75t_L g109 ( .A1(n_49), .A2(n_60), .B1(n_104), .B2(n_108), .Y(n_109) );
INVx1_ASAP7_75t_L g129 ( .A(n_49), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_50), .B(n_256), .Y(n_255) );
XOR2xp5_ASAP7_75t_L g635 ( .A(n_51), .B(n_95), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_52), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_54), .B(n_239), .Y(n_238) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_56), .B(n_266), .Y(n_319) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_58), .Y(n_358) );
INVx1_ASAP7_75t_L g121 ( .A(n_59), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_59), .B(n_127), .Y(n_175) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_59), .Y(n_204) );
OAI21xp33_ASAP7_75t_L g130 ( .A1(n_60), .A2(n_66), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_62), .B(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_66), .B(n_73), .Y(n_173) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_67), .Y(n_219) );
BUFx5_ASAP7_75t_L g250 ( .A(n_67), .Y(n_250) );
INVx1_ASAP7_75t_L g274 ( .A(n_67), .Y(n_274) );
INVx2_ASAP7_75t_L g394 ( .A(n_68), .Y(n_394) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_69), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_SL g210 ( .A(n_70), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_71), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_72), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_73), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_76), .B(n_264), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_196), .B1(n_213), .B2(n_227), .C(n_629), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_92), .Y(n_78) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_85), .B1(n_90), .B2(n_91), .Y(n_79) );
INVx1_ASAP7_75t_L g90 ( .A(n_80), .Y(n_90) );
OAI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_80) );
INVx1_ASAP7_75t_L g84 ( .A(n_81), .Y(n_84) );
INVx1_ASAP7_75t_L g83 ( .A(n_82), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_85), .Y(n_91) );
OAI22xp5_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_86), .Y(n_89) );
INVx1_ASAP7_75t_L g88 ( .A(n_87), .Y(n_88) );
AOI22xp5_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_95), .B1(n_194), .B2(n_195), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_93), .Y(n_194) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g195 ( .A(n_95), .Y(n_195) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NOR2x1_ASAP7_75t_L g96 ( .A(n_97), .B(n_159), .Y(n_96) );
NAND4xp25_ASAP7_75t_SL g97 ( .A(n_98), .B(n_132), .C(n_142), .D(n_149), .Y(n_97) );
BUFx4f_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_110), .Y(n_100) );
AND2x4_ASAP7_75t_L g144 ( .A(n_101), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g163 ( .A(n_101), .B(n_157), .Y(n_163) );
AND2x2_ASAP7_75t_L g178 ( .A(n_101), .B(n_153), .Y(n_178) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_109), .Y(n_101) );
INVx1_ASAP7_75t_L g136 ( .A(n_102), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx2_ASAP7_75t_L g108 ( .A(n_104), .Y(n_108) );
INVx3_ASAP7_75t_L g113 ( .A(n_104), .Y(n_113) );
NAND2xp33_ASAP7_75t_L g120 ( .A(n_104), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_104), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_105), .B(n_129), .Y(n_128) );
INVxp67_ASAP7_75t_L g205 ( .A(n_105), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_107), .A2(n_131), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
AND2x2_ASAP7_75t_L g162 ( .A(n_109), .B(n_136), .Y(n_162) );
AND2x2_ASAP7_75t_L g185 ( .A(n_109), .B(n_186), .Y(n_185) );
AND2x4_ASAP7_75t_L g124 ( .A(n_110), .B(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g134 ( .A(n_110), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
OR2x2_ASAP7_75t_L g141 ( .A(n_111), .B(n_116), .Y(n_141) );
AND2x4_ASAP7_75t_L g153 ( .A(n_111), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g158 ( .A(n_111), .Y(n_158) );
AND2x2_ASAP7_75t_L g182 ( .A(n_111), .B(n_183), .Y(n_182) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_113), .B(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g127 ( .A(n_113), .Y(n_127) );
NAND3xp33_ASAP7_75t_L g174 ( .A(n_114), .B(n_126), .C(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx8_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g148 ( .A(n_125), .B(n_140), .Y(n_148) );
AND2x4_ASAP7_75t_L g193 ( .A(n_125), .B(n_157), .Y(n_193) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
BUFx12f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g139 ( .A(n_135), .B(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g152 ( .A(n_135), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g156 ( .A(n_135), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g145 ( .A(n_141), .Y(n_145) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx6_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g161 ( .A(n_153), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g157 ( .A(n_154), .B(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g190 ( .A(n_157), .B(n_162), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .C(n_188), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_174), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_170), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_185), .Y(n_181) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_184), .Y(n_202) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
XOR2xp5_ASAP7_75t_L g630 ( .A(n_195), .B(n_631), .Y(n_630) );
BUFx10_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_207), .Y(n_198) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g634 ( .A(n_200), .B(n_207), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_206), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_211), .Y(n_207) );
OR2x2_ASAP7_75t_L g637 ( .A(n_208), .B(n_212), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_208), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_208), .B(n_211), .Y(n_641) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_215), .B(n_225), .Y(n_214) );
OA21x2_ASAP7_75t_L g639 ( .A1(n_215), .A2(n_640), .B(n_641), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g300 ( .A(n_218), .Y(n_300) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx6_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
INVx3_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
INVx2_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_222), .B(n_293), .Y(n_292) );
OAI22x1_ASAP7_75t_L g347 ( .A1(n_222), .A2(n_348), .B1(n_352), .B2(n_353), .Y(n_347) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_223), .A2(n_245), .B(n_248), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_223), .A2(n_291), .B1(n_292), .B2(n_295), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_223), .B(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_224), .Y(n_258) );
INVxp67_ASAP7_75t_L g314 ( .A(n_224), .Y(n_314) );
INVx1_ASAP7_75t_L g336 ( .A(n_224), .Y(n_336) );
INVx4_ASAP7_75t_L g366 ( .A(n_224), .Y(n_366) );
INVx3_ASAP7_75t_L g375 ( .A(n_224), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_224), .B(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_224), .B(n_387), .Y(n_386) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_225), .A2(n_290), .B(n_298), .Y(n_289) );
AO31x2_ASAP7_75t_L g346 ( .A1(n_225), .A2(n_347), .A3(n_356), .B(n_357), .Y(n_346) );
AO31x2_ASAP7_75t_L g411 ( .A1(n_225), .A2(n_347), .A3(n_356), .B(n_357), .Y(n_411) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
INVx1_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
INVx3_ASAP7_75t_L g331 ( .A(n_226), .Y(n_331) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_531), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_449), .C(n_494), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_425), .Y(n_232) );
AOI211x1_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_361), .B(n_395), .C(n_416), .Y(n_233) );
OAI21xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_285), .B(n_343), .Y(n_234) );
OR2x2_ASAP7_75t_L g440 ( .A(n_235), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g527 ( .A(n_236), .B(n_528), .Y(n_527) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_236), .A2(n_561), .B(n_562), .C(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g572 ( .A(n_236), .B(n_441), .Y(n_572) );
AND2x2_ASAP7_75t_L g575 ( .A(n_236), .B(n_406), .Y(n_575) );
AND2x2_ASAP7_75t_L g605 ( .A(n_236), .B(n_430), .Y(n_605) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_261), .Y(n_236) );
INVx3_ASAP7_75t_L g415 ( .A(n_237), .Y(n_415) );
INVx2_ASAP7_75t_L g445 ( .A(n_237), .Y(n_445) );
AND2x2_ASAP7_75t_L g488 ( .A(n_237), .B(n_404), .Y(n_488) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_239), .B(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_240), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx4_ASAP7_75t_L g267 ( .A(n_241), .Y(n_267) );
BUFx3_ASAP7_75t_L g284 ( .A(n_241), .Y(n_284) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_251), .B(n_259), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g310 ( .A(n_247), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx2_ASAP7_75t_L g291 ( .A(n_249), .Y(n_291) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g256 ( .A(n_250), .Y(n_256) );
INVx2_ASAP7_75t_L g275 ( .A(n_250), .Y(n_275) );
INVx2_ASAP7_75t_L g355 ( .A(n_250), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_255), .B(n_257), .Y(n_251) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
INVx2_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g269 ( .A(n_258), .Y(n_269) );
INVx2_ASAP7_75t_SL g280 ( .A(n_258), .Y(n_280) );
INVxp67_ASAP7_75t_L g302 ( .A(n_258), .Y(n_302) );
INVx2_ASAP7_75t_L g324 ( .A(n_260), .Y(n_324) );
INVx2_ASAP7_75t_SL g404 ( .A(n_261), .Y(n_404) );
AND2x2_ASAP7_75t_L g414 ( .A(n_261), .B(n_415), .Y(n_414) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_268), .B(n_281), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_262), .A2(n_268), .B(n_281), .Y(n_453) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g370 ( .A(n_265), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g323 ( .A(n_267), .Y(n_323) );
AOI21x1_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_276), .Y(n_268) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g351 ( .A(n_274), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_275), .A2(n_300), .B1(n_389), .B2(n_391), .Y(n_388) );
AOI21x1_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_280), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_280), .B(n_319), .Y(n_320) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NOR2xp67_ASAP7_75t_SL g357 ( .A(n_283), .B(n_358), .Y(n_357) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_284), .A2(n_289), .B(n_303), .Y(n_288) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_284), .A2(n_289), .B(n_303), .Y(n_360) );
NOR2x1_ASAP7_75t_SL g489 ( .A(n_285), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_304), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_286), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g566 ( .A(n_286), .B(n_543), .Y(n_566) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g435 ( .A(n_287), .B(n_326), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_287), .B(n_400), .Y(n_467) );
AND2x2_ASAP7_75t_L g608 ( .A(n_287), .B(n_346), .Y(n_608) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g409 ( .A(n_288), .Y(n_409) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_288), .Y(n_511) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_302), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_300), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_326), .Y(n_304) );
INVx1_ASAP7_75t_L g398 ( .A(n_305), .Y(n_398) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g344 ( .A(n_306), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g448 ( .A(n_306), .Y(n_448) );
INVxp67_ASAP7_75t_L g581 ( .A(n_306), .Y(n_581) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_315), .B(n_321), .Y(n_306) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_307), .A2(n_315), .B(n_321), .Y(n_422) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B(n_314), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_309), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
OAI21x1_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B(n_320), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g325 ( .A(n_319), .Y(n_325) );
AOI21xp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B(n_325), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_324), .B(n_366), .C(n_367), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_324), .B(n_367), .C(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g400 ( .A(n_326), .Y(n_400) );
INVx1_ASAP7_75t_L g407 ( .A(n_326), .Y(n_407) );
INVx1_ASAP7_75t_L g625 ( .A(n_326), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_327), .B(n_334), .Y(n_326) );
AND2x2_ASAP7_75t_L g462 ( .A(n_327), .B(n_334), .Y(n_462) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_329), .B(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g342 ( .A(n_330), .Y(n_342) );
INVx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVx1_ASAP7_75t_L g356 ( .A(n_341), .Y(n_356) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_359), .Y(n_343) );
INVx1_ASAP7_75t_L g469 ( .A(n_344), .Y(n_469) );
INVx2_ASAP7_75t_L g424 ( .A(n_345), .Y(n_424) );
INVx1_ASAP7_75t_L g438 ( .A(n_345), .Y(n_438) );
AND2x2_ASAP7_75t_L g471 ( .A(n_345), .B(n_400), .Y(n_471) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_359), .B(n_447), .Y(n_477) );
AND2x2_ASAP7_75t_L g580 ( .A(n_359), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g464 ( .A(n_360), .B(n_422), .Y(n_464) );
AND2x2_ASAP7_75t_L g579 ( .A(n_360), .B(n_462), .Y(n_579) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_362), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g553 ( .A(n_362), .B(n_414), .Y(n_553) );
INVx2_ASAP7_75t_L g562 ( .A(n_362), .Y(n_562) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_377), .Y(n_362) );
INVx1_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_363), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g430 ( .A(n_363), .B(n_378), .Y(n_430) );
INVx1_ASAP7_75t_L g442 ( .A(n_363), .Y(n_442) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_363), .Y(n_456) );
INVx1_ASAP7_75t_L g487 ( .A(n_363), .Y(n_487) );
INVx2_ASAP7_75t_L g493 ( .A(n_363), .Y(n_493) );
AND2x2_ASAP7_75t_L g536 ( .A(n_363), .B(n_415), .Y(n_536) );
OR2x6_ASAP7_75t_L g363 ( .A(n_364), .B(n_372), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B(n_370), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g389 ( .A(n_366), .B(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_366), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g380 ( .A(n_367), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g492 ( .A(n_377), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g403 ( .A(n_378), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
OR2x2_ASAP7_75t_L g452 ( .A(n_378), .B(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g530 ( .A(n_378), .Y(n_530) );
INVx1_ASAP7_75t_L g564 ( .A(n_378), .Y(n_564) );
AO21x2_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_393), .Y(n_378) );
NAND3xp33_ASAP7_75t_SL g381 ( .A(n_382), .B(n_385), .C(n_388), .Y(n_381) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .A3(n_401), .B1(n_405), .B2(n_412), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g595 ( .A(n_398), .B(n_467), .Y(n_595) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g497 ( .A(n_402), .B(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_402), .Y(n_538) );
AND2x4_ASAP7_75t_L g535 ( .A(n_403), .B(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g546 ( .A(n_403), .Y(n_546) );
INVx1_ASAP7_75t_L g507 ( .A(n_404), .Y(n_507) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g501 ( .A(n_407), .Y(n_501) );
INVx1_ASAP7_75t_L g568 ( .A(n_407), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x4_ASAP7_75t_L g421 ( .A(n_409), .B(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_409), .Y(n_591) );
INVx1_ASAP7_75t_L g551 ( .A(n_410), .Y(n_551) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g447 ( .A(n_411), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g526 ( .A(n_411), .B(n_422), .Y(n_526) );
OR2x2_ASAP7_75t_L g543 ( .A(n_411), .B(n_422), .Y(n_543) );
INVx1_ASAP7_75t_L g559 ( .A(n_413), .Y(n_559) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g417 ( .A(n_414), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
AND2x2_ASAP7_75t_L g491 ( .A(n_414), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g506 ( .A(n_415), .Y(n_506) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_417), .A2(n_577), .B1(n_578), .B2(n_580), .Y(n_576) );
INVx2_ASAP7_75t_L g589 ( .A(n_417), .Y(n_589) );
INVx2_ASAP7_75t_L g558 ( .A(n_418), .Y(n_558) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_421), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_421), .B(n_471), .Y(n_485) );
BUFx3_ASAP7_75t_L g519 ( .A(n_421), .Y(n_519) );
INVx1_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
AND2x2_ASAP7_75t_L g552 ( .A(n_423), .B(n_435), .Y(n_552) );
AND2x2_ASAP7_75t_L g573 ( .A(n_423), .B(n_464), .Y(n_573) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g433 ( .A(n_424), .Y(n_433) );
AND2x2_ASAP7_75t_L g516 ( .A(n_424), .B(n_461), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_431), .B(n_439), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g569 ( .A(n_427), .Y(n_569) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_430), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_430), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_432), .B(n_436), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_433), .B(n_575), .Y(n_599) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_436), .A2(n_440), .B1(n_443), .B2(n_446), .Y(n_439) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
NAND2xp67_ASAP7_75t_L g499 ( .A(n_437), .B(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_437), .A2(n_621), .B1(n_627), .B2(n_628), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_438), .B(n_613), .Y(n_619) );
OR2x2_ASAP7_75t_L g504 ( .A(n_441), .B(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_441), .Y(n_601) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g478 ( .A(n_442), .B(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g557 ( .A(n_444), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g561 ( .A(n_444), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_444), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g451 ( .A(n_445), .B(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
AND2x2_ASAP7_75t_L g513 ( .A(n_445), .B(n_487), .Y(n_513) );
AND2x2_ASAP7_75t_L g545 ( .A(n_447), .B(n_525), .Y(n_545) );
AND2x4_ASAP7_75t_L g578 ( .A(n_447), .B(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g596 ( .A(n_447), .Y(n_596) );
BUFx3_ASAP7_75t_L g627 ( .A(n_447), .Y(n_627) );
INVx1_ASAP7_75t_L g512 ( .A(n_448), .Y(n_512) );
OAI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_457), .B(n_472), .C(n_483), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_451), .A2(n_603), .B1(n_604), .B2(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
INVx2_ASAP7_75t_L g479 ( .A(n_452), .Y(n_479) );
BUFx2_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g594 ( .A(n_456), .B(n_479), .Y(n_594) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_465), .C(n_468), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g525 ( .A(n_461), .Y(n_525) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g482 ( .A(n_463), .Y(n_482) );
INVx1_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g550 ( .A(n_467), .Y(n_550) );
NAND2xp33_ASAP7_75t_SL g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_469), .B(n_529), .Y(n_574) );
NOR2x1_ASAP7_75t_R g518 ( .A(n_470), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_471), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_476), .B1(n_478), .B2(n_480), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g628 ( .A(n_478), .B(n_623), .Y(n_628) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_481), .B(n_591), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B(n_489), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g614 ( .A(n_488), .Y(n_614) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_499), .B(n_502), .C(n_517), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g523 ( .A(n_498), .Y(n_523) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g541 ( .A(n_501), .B(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_508), .B1(n_513), .B2(n_514), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2xp67_ASAP7_75t_SL g587 ( .A(n_505), .B(n_564), .Y(n_587) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g540 ( .A(n_506), .Y(n_540) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
NAND2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_546), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g544 ( .A1(n_514), .A2(n_545), .B(n_546), .Y(n_544) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B1(n_524), .B2(n_527), .Y(n_517) );
INVx2_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AND2x2_ASAP7_75t_L g567 ( .A(n_526), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g616 ( .A(n_526), .Y(n_616) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_582), .Y(n_531) );
NOR2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_554), .Y(n_532) );
NAND3xp33_ASAP7_75t_SL g533 ( .A(n_534), .B(n_544), .C(n_547), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_537), .B(n_541), .Y(n_534) );
INVx2_ASAP7_75t_L g618 ( .A(n_535), .Y(n_618) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g623 ( .A(n_540), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_552), .B(n_553), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_552), .B(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_555), .B(n_570), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_565), .B1(n_567), .B2(n_569), .Y(n_555) );
AO21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B(n_560), .Y(n_556) );
OR2x2_ASAP7_75t_L g613 ( .A(n_558), .B(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_563), .Y(n_577) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_571) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_609), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_597), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .C(n_592), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_589), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g603 ( .A(n_591), .Y(n_603) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g626 ( .A(n_594), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_602), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_606), .B(n_618), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_620), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_617), .C(n_619), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_615), .B2(n_616), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI222xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_633), .B2(n_635), .C1(n_636), .C2(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
endmodule