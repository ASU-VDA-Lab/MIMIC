module fake_jpeg_31751_n_42 (n_3, n_2, n_1, n_0, n_4, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_5;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_1),
.Y(n_5)
);

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

A2O1A1Ixp33_ASAP7_75t_L g10 ( 
.A1(n_7),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_6),
.B1(n_9),
.B2(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_10),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.C(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_11),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_22),
.B2(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_6),
.B1(n_14),
.B2(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_23),
.B1(n_6),
.B2(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_2),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_32),
.B(n_27),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_36),
.B(n_4),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_2),
.C(n_3),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_4),
.CI(n_32),
.CON(n_37),
.SN(n_37)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_38),
.B(n_0),
.Y(n_40)
);

OAI311xp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_0),
.A3(n_1),
.B1(n_33),
.C1(n_34),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_40),
.B(n_37),
.C(n_0),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_0),
.Y(n_42)
);


endmodule