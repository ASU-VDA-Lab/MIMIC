module fake_jpeg_14164_n_305 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_305);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_265;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_156;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_70),
.Y(n_98)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_48),
.B1(n_64),
.B2(n_49),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_82),
.B1(n_85),
.B2(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_35),
.B1(n_25),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_92),
.B1(n_104),
.B2(n_66),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_35),
.B1(n_29),
.B2(n_21),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_24),
.C(n_37),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_88),
.C(n_16),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_37),
.C(n_33),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_51),
.B1(n_55),
.B2(n_66),
.Y(n_91)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_65),
.B1(n_54),
.B2(n_53),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_43),
.B1(n_33),
.B2(n_21),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_111),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_96),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_3),
.B(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_42),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_9),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_44),
.A2(n_38),
.B1(n_42),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_38),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_119),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_97),
.B1(n_75),
.B2(n_101),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_118),
.A2(n_122),
.B1(n_105),
.B2(n_76),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_65),
.B1(n_55),
.B2(n_63),
.Y(n_122)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_90),
.B1(n_77),
.B2(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_17),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_9),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_75),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

CKINVDCx12_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_16),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_16),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_108),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_167),
.B1(n_176),
.B2(n_116),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_161),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_80),
.B(n_101),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_180),
.B(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_165),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_75),
.B1(n_91),
.B2(n_79),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_74),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_137),
.B(n_114),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_173),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_91),
.B1(n_110),
.B2(n_109),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_126),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_122),
.A2(n_79),
.B1(n_83),
.B2(n_77),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_179),
.B1(n_146),
.B2(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_83),
.B1(n_77),
.B2(n_110),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_74),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_189),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_123),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_191),
.B(n_196),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_203),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_123),
.B1(n_135),
.B2(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_130),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_140),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_202),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_125),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_199),
.B(n_164),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_141),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_197),
.C(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_204),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_142),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_125),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_125),
.B(n_117),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_113),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_132),
.B1(n_89),
.B2(n_125),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_170),
.B1(n_165),
.B2(n_167),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_150),
.B(n_132),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_90),
.B1(n_116),
.B2(n_127),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_112),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_112),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_223),
.B(n_230),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_170),
.C(n_157),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_169),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_165),
.B1(n_151),
.B2(n_168),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_225),
.B1(n_199),
.B2(n_191),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_159),
.C(n_178),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_186),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_196),
.A2(n_155),
.B(n_172),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_149),
.B1(n_162),
.B2(n_163),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_159),
.C(n_154),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_155),
.C(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_236),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_238),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_203),
.B1(n_198),
.B2(n_207),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_194),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_243),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_204),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_209),
.B(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_205),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_209),
.B1(n_228),
.B2(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_255),
.B(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_220),
.B1(n_214),
.B2(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_253),
.B1(n_187),
.B2(n_184),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_214),
.B1(n_191),
.B2(n_231),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_216),
.B1(n_211),
.B2(n_192),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_211),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_218),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_234),
.B1(n_248),
.B2(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_242),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_237),
.A3(n_238),
.B1(n_244),
.B2(n_184),
.C1(n_242),
.C2(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_181),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_272),
.B(n_273),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_258),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_263),
.B(n_250),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_252),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_195),
.C(n_208),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_261),
.C(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_275),
.C(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_253),
.C(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_149),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_160),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_264),
.B1(n_268),
.B2(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_270),
.B(n_266),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_291),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_269),
.C(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_160),
.C(n_162),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_284),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_283),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_276),
.B1(n_282),
.B2(n_281),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_295),
.B(n_293),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_156),
.C(n_127),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_293),
.B(n_156),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_300),
.C(n_156),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_112),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_112),
.Y(n_305)
);


endmodule