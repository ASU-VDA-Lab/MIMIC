module fake_netlist_5_1299_n_575 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_575);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_575;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_378;
wire n_551;
wire n_382;
wire n_554;
wire n_254;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_559;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_145;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_66),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_51),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_27),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_32),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_43),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_5),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_20),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_77),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_23),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_19),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_49),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

INVx4_ASAP7_75t_R g165 ( 
.A(n_36),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_16),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_37),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_7),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_45),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_28),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_30),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_38),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_39),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_101),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_60),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_26),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_0),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_154),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_136),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_137),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_140),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_156),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_141),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_144),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_157),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_139),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_177),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_143),
.B(n_153),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_172),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_177),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_139),
.Y(n_250)
);

AND2x2_ASAP7_75t_R g251 ( 
.A(n_206),
.B(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_139),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_167),
.B(n_183),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_R g264 ( 
.A(n_203),
.B(n_0),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_216),
.B(n_167),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_185),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_146),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_278),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_149),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_167),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_150),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_167),
.B1(n_181),
.B2(n_176),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_151),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_239),
.B(n_152),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_274),
.B(n_1),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_155),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_160),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_238),
.A2(n_182),
.B1(n_168),
.B2(n_166),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_161),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_1),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_246),
.B(n_262),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_242),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

AO22x2_ASAP7_75t_L g314 ( 
.A1(n_270),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_314)
);

NOR2x1p5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_242),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_4),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_13),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

AND3x1_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_8),
.C(n_9),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_14),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_270),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_243),
.B(n_15),
.Y(n_325)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_267),
.B(n_18),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_234),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_247),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_242),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_231),
.B(n_9),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_231),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_274),
.B(n_10),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

OAI221xp5_ASAP7_75t_L g338 ( 
.A1(n_289),
.A2(n_264),
.B1(n_240),
.B2(n_269),
.C(n_276),
.Y(n_338)
);

AO22x2_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_276),
.B1(n_277),
.B2(n_275),
.Y(n_339)
);

AO22x2_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_251),
.B1(n_273),
.B2(n_12),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_273),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

NAND2x1p5_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_274),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

NAND2x1p5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_274),
.Y(n_349)
);

NAND2x1p5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_254),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_335),
.A2(n_11),
.B1(n_12),
.B2(n_254),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_21),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_250),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_250),
.Y(n_354)
);

NAND2x1p5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_22),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_24),
.Y(n_360)
);

AO22x2_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_303),
.A2(n_250),
.B1(n_253),
.B2(n_235),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_310),
.B(n_253),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_253),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g367 ( 
.A(n_317),
.B(n_41),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_292),
.B(n_250),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g373 ( 
.A(n_280),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_295),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_297),
.B(n_58),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

AO22x2_ASAP7_75t_L g379 ( 
.A1(n_282),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_379)
);

NAND2x1_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_64),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_282),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_287),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_304),
.B(n_75),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_287),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_317),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_387),
.B(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_348),
.B(n_311),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_342),
.B(n_311),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_291),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_366),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_346),
.B(n_311),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_385),
.B(n_352),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_388),
.B(n_302),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_344),
.B(n_299),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_336),
.B(n_302),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_380),
.B(n_325),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_337),
.B(n_309),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_341),
.B(n_284),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_343),
.B(n_284),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_345),
.B(n_284),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_384),
.B(n_333),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_349),
.B(n_286),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_360),
.B(n_370),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_286),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_353),
.B(n_371),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_367),
.B(n_286),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_377),
.B(n_326),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_378),
.B(n_326),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_339),
.B(n_340),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_SL g414 ( 
.A(n_364),
.B(n_321),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_355),
.B(n_321),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_369),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_347),
.B(n_76),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_357),
.B(n_78),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_368),
.B(n_79),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_354),
.B(n_81),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_82),
.Y(n_422)
);

AOI221x1_ASAP7_75t_L g423 ( 
.A1(n_411),
.A2(n_376),
.B1(n_374),
.B2(n_361),
.C(n_362),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_422),
.A2(n_350),
.B(n_365),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_338),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_412),
.A2(n_421),
.B(n_416),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_339),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_351),
.Y(n_429)
);

O2A1O1Ixp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_376),
.B(n_351),
.C(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_362),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

NAND2x1p5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_363),
.Y(n_434)
);

OAI22x1_ASAP7_75t_L g435 ( 
.A1(n_392),
.A2(n_361),
.B1(n_374),
.B2(n_340),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_391),
.A2(n_375),
.B(n_381),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

AO31x2_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_383),
.A3(n_381),
.B(n_379),
.Y(n_438)
);

AOI211x1_ASAP7_75t_L g439 ( 
.A1(n_421),
.A2(n_420),
.B(n_419),
.C(n_417),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_400),
.A2(n_383),
.B(n_375),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_409),
.A2(n_373),
.B(n_85),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_415),
.B(n_84),
.Y(n_442)
);

NOR2x1_ASAP7_75t_R g443 ( 
.A(n_397),
.B(n_86),
.Y(n_443)
);

BUFx12f_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

O2A1O1Ixp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_406),
.B1(n_404),
.B2(n_403),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_402),
.Y(n_449)
);

O2A1O1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_99),
.B(n_100),
.C(n_102),
.Y(n_450)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_431),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_447),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_435),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_124),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_437),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_112),
.B(n_113),
.C(n_117),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

AO21x2_ASAP7_75t_L g461 ( 
.A1(n_427),
.A2(n_118),
.B(n_119),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_436),
.A2(n_123),
.B1(n_441),
.B2(n_434),
.Y(n_462)
);

A2O1A1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_436),
.A2(n_442),
.B(n_445),
.C(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_439),
.Y(n_466)
);

AO21x2_ASAP7_75t_L g467 ( 
.A1(n_438),
.A2(n_424),
.B(n_440),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

AO32x2_ASAP7_75t_L g469 ( 
.A1(n_438),
.A2(n_423),
.A3(n_430),
.B1(n_436),
.B2(n_323),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_453),
.B(n_463),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_467),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_460),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_466),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_458),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

BUFx2_ASAP7_75t_SL g477 ( 
.A(n_457),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

OAI21x1_ASAP7_75t_SL g479 ( 
.A1(n_468),
.A2(n_462),
.B(n_464),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_465),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_461),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_450),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_453),
.A2(n_462),
.B1(n_279),
.B2(n_464),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_451),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_487),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_484),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_475),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_473),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_495),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_R g502 ( 
.A(n_495),
.B(n_488),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_494),
.B(n_470),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_474),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_479),
.B(n_482),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_496),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_R g509 ( 
.A(n_488),
.B(n_480),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_472),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_480),
.B(n_491),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_480),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_R g513 ( 
.A(n_491),
.B(n_482),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_491),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_480),
.B(n_472),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_482),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_496),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_518),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_485),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_508),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_476),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_517),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_515),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_501),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_489),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_519),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_516),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_516),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_516),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_507),
.Y(n_537)
);

AOI211xp5_ASAP7_75t_L g538 ( 
.A1(n_525),
.A2(n_504),
.B(n_493),
.C(n_511),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_524),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_535),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_539),
.B(n_524),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_532),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_530),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_530),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_528),
.Y(n_546)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_531),
.Y(n_547)
);

AO221x2_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_527),
.B1(n_526),
.B2(n_529),
.C(n_522),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_546),
.A2(n_513),
.B1(n_537),
.B2(n_533),
.Y(n_549)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_510),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_546),
.A2(n_513),
.B1(n_537),
.B2(n_533),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_545),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_547),
.B(n_544),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_550),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_549),
.B(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_551),
.Y(n_556)
);

NAND4xp25_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_555),
.C(n_554),
.D(n_538),
.Y(n_557)
);

O2A1O1Ixp5_ASAP7_75t_L g558 ( 
.A1(n_555),
.A2(n_537),
.B(n_511),
.C(n_514),
.Y(n_558)
);

AOI322xp5_ASAP7_75t_L g559 ( 
.A1(n_553),
.A2(n_541),
.A3(n_493),
.B1(n_543),
.B2(n_514),
.C1(n_520),
.C2(n_492),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_552),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_558),
.A2(n_482),
.B(n_507),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_560),
.Y(n_562)
);

NAND4xp25_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_561),
.C(n_559),
.D(n_502),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_563),
.A2(n_529),
.B1(n_503),
.B2(n_506),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_564),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_R g566 ( 
.A(n_565),
.B(n_498),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_482),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_498),
.B1(n_523),
.B2(n_507),
.Y(n_569)
);

AOI31xp33_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_515),
.A3(n_476),
.B(n_492),
.Y(n_570)
);

BUFx2_ASAP7_75t_SL g571 ( 
.A(n_570),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_571),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_572),
.Y(n_573)
);

AOI221xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_523),
.B1(n_472),
.B2(n_481),
.C(n_486),
.Y(n_574)
);

AOI211xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_483),
.B(n_486),
.C(n_471),
.Y(n_575)
);


endmodule