module real_jpeg_1318_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_36),
.B1(n_41),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_3),
.A2(n_36),
.B1(n_41),
.B2(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_31),
.B(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_48),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_24),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_36),
.C(n_84),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_4),
.B(n_38),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_4),
.B(n_89),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_36),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_36),
.B1(n_41),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_67),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_11),
.A2(n_30),
.B1(n_32),
.B2(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_11),
.A2(n_36),
.B1(n_41),
.B2(n_56),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_12),
.A2(n_30),
.B1(n_32),
.B2(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_12),
.A2(n_36),
.B1(n_41),
.B2(n_59),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_81),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_13),
.A2(n_36),
.B1(n_41),
.B2(n_81),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_113),
.B1(n_185),
.B2(n_186),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_19),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_21),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_21),
.B(n_115),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_45),
.CI(n_68),
.CON(n_21),
.SN(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_34),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_24),
.A2(n_25),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_24),
.A2(n_50),
.A3(n_52),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_25),
.B(n_124),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_35),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_35),
.A2(n_38),
.B1(n_128),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_35),
.A2(n_38),
.B1(n_124),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_35),
.A2(n_38),
.B1(n_165),
.B2(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_36),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_36),
.A2(n_41),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_36),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_37),
.A2(n_43),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_37),
.A2(n_105),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_37),
.A2(n_105),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_60),
.C(n_64),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_46),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_57),
.B1(n_77),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_47),
.A2(n_55),
.B1(n_57),
.B2(n_144),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AO22x2_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_50),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_49),
.B(n_53),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_50),
.B(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_70),
.B1(n_74),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_76),
.C(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_90),
.B2(n_91),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_87),
.B2(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_82),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_89),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_82),
.A2(n_89),
.B1(n_135),
.B2(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_88),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_86),
.A2(n_109),
.B1(n_120),
.B2(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_130),
.B(n_184),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_121),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_121),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_179),
.B(n_183),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_148),
.B(n_178),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_138),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_137),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_143),
.C(n_146),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_159),
.B(n_177),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_157),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_171),
.B(n_176),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_170),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_175),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_182),
.Y(n_183)
);


endmodule