module fake_jpeg_28531_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_29),
.B1(n_31),
.B2(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_16),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_47),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_13),
.B1(n_18),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_14),
.B1(n_13),
.B2(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_61),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_26),
.B(n_31),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_56),
.C(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_32),
.B(n_29),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_20),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_18),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_56),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_20),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_16),
.B1(n_18),
.B2(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_12),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

AOI221xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_85),
.B1(n_86),
.B2(n_82),
.C(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_64),
.B1(n_61),
.B2(n_54),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_75),
.B(n_70),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_67),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_70),
.C(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_12),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_68),
.C(n_77),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_85),
.C(n_15),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_97),
.C(n_89),
.Y(n_99)
);

NAND4xp25_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_19),
.C(n_21),
.D(n_9),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_53),
.B1(n_15),
.B2(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_101),
.B1(n_37),
.B2(n_48),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_60),
.B1(n_37),
.B2(n_39),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_105),
.B(n_41),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_95),
.B(n_94),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_99),
.B(n_102),
.C(n_100),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.A3(n_103),
.B1(n_35),
.B2(n_8),
.C1(n_7),
.C2(n_44),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_7),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_8),
.B1(n_41),
.B2(n_44),
.C(n_109),
.Y(n_111)
);


endmodule